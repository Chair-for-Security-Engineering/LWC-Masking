/* modified netlist. Source: module SubCells in file ./test/SubCells.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module SubCells_HPC2_ClockGating_d2 (SubC_in_s0, clk, SubC_in_s1, SubC_in_s2, Fresh, /*rst,*/ SubC_out_s0, SubC_out_s1, SubC_out_s2/*, Synch*/);
    input [127:0] SubC_in_s0 ;
    input clk ;
    input [127:0] SubC_in_s1 ;
    input [127:0] SubC_in_s2 ;
    //input rst ;
    input [575:0] Fresh ;
    output [127:0] SubC_out_s0 ;
    output [127:0] SubC_out_s1 ;
    output [127:0] SubC_out_s2 ;
    //output Synch ;
    wire SB_31_n15 ;
    wire SB_31_n14 ;
    wire SB_31_n13 ;
    wire SB_31_n12 ;
    wire SB_31_n11 ;
    wire SB_31_n10 ;
    wire SB_31_n9 ;
    wire SB_31_T5 ;
    wire SB_31_T4 ;
    wire SB_31_T3 ;
    wire SB_31_T2 ;
    wire SB_31_T1 ;
    wire SB_31_T0 ;
    wire SB_30_n15 ;
    wire SB_30_n14 ;
    wire SB_30_n13 ;
    wire SB_30_n12 ;
    wire SB_30_n11 ;
    wire SB_30_n10 ;
    wire SB_30_n9 ;
    wire SB_30_T5 ;
    wire SB_30_T4 ;
    wire SB_30_T3 ;
    wire SB_30_T2 ;
    wire SB_30_T1 ;
    wire SB_30_T0 ;
    wire SB_29_n15 ;
    wire SB_29_n14 ;
    wire SB_29_n13 ;
    wire SB_29_n12 ;
    wire SB_29_n11 ;
    wire SB_29_n10 ;
    wire SB_29_n9 ;
    wire SB_29_T5 ;
    wire SB_29_T4 ;
    wire SB_29_T3 ;
    wire SB_29_T2 ;
    wire SB_29_T1 ;
    wire SB_29_T0 ;
    wire SB_28_n15 ;
    wire SB_28_n14 ;
    wire SB_28_n13 ;
    wire SB_28_n12 ;
    wire SB_28_n11 ;
    wire SB_28_n10 ;
    wire SB_28_n9 ;
    wire SB_28_T5 ;
    wire SB_28_T4 ;
    wire SB_28_T3 ;
    wire SB_28_T2 ;
    wire SB_28_T1 ;
    wire SB_28_T0 ;
    wire SB_27_n15 ;
    wire SB_27_n14 ;
    wire SB_27_n13 ;
    wire SB_27_n12 ;
    wire SB_27_n11 ;
    wire SB_27_n10 ;
    wire SB_27_n9 ;
    wire SB_27_T5 ;
    wire SB_27_T4 ;
    wire SB_27_T3 ;
    wire SB_27_T2 ;
    wire SB_27_T1 ;
    wire SB_27_T0 ;
    wire SB_26_n15 ;
    wire SB_26_n14 ;
    wire SB_26_n13 ;
    wire SB_26_n12 ;
    wire SB_26_n11 ;
    wire SB_26_n10 ;
    wire SB_26_n9 ;
    wire SB_26_T5 ;
    wire SB_26_T4 ;
    wire SB_26_T3 ;
    wire SB_26_T2 ;
    wire SB_26_T1 ;
    wire SB_26_T0 ;
    wire SB_25_n15 ;
    wire SB_25_n14 ;
    wire SB_25_n13 ;
    wire SB_25_n12 ;
    wire SB_25_n11 ;
    wire SB_25_n10 ;
    wire SB_25_n9 ;
    wire SB_25_T5 ;
    wire SB_25_T4 ;
    wire SB_25_T3 ;
    wire SB_25_T2 ;
    wire SB_25_T1 ;
    wire SB_25_T0 ;
    wire SB_24_n15 ;
    wire SB_24_n14 ;
    wire SB_24_n13 ;
    wire SB_24_n12 ;
    wire SB_24_n11 ;
    wire SB_24_n10 ;
    wire SB_24_n9 ;
    wire SB_24_T5 ;
    wire SB_24_T4 ;
    wire SB_24_T3 ;
    wire SB_24_T2 ;
    wire SB_24_T1 ;
    wire SB_24_T0 ;
    wire SB_23_n15 ;
    wire SB_23_n14 ;
    wire SB_23_n13 ;
    wire SB_23_n12 ;
    wire SB_23_n11 ;
    wire SB_23_n10 ;
    wire SB_23_n9 ;
    wire SB_23_T5 ;
    wire SB_23_T4 ;
    wire SB_23_T3 ;
    wire SB_23_T2 ;
    wire SB_23_T1 ;
    wire SB_23_T0 ;
    wire SB_22_n15 ;
    wire SB_22_n14 ;
    wire SB_22_n13 ;
    wire SB_22_n12 ;
    wire SB_22_n11 ;
    wire SB_22_n10 ;
    wire SB_22_n9 ;
    wire SB_22_T5 ;
    wire SB_22_T4 ;
    wire SB_22_T3 ;
    wire SB_22_T2 ;
    wire SB_22_T1 ;
    wire SB_22_T0 ;
    wire SB_21_n15 ;
    wire SB_21_n14 ;
    wire SB_21_n13 ;
    wire SB_21_n12 ;
    wire SB_21_n11 ;
    wire SB_21_n10 ;
    wire SB_21_n9 ;
    wire SB_21_T5 ;
    wire SB_21_T4 ;
    wire SB_21_T3 ;
    wire SB_21_T2 ;
    wire SB_21_T1 ;
    wire SB_21_T0 ;
    wire SB_20_n15 ;
    wire SB_20_n14 ;
    wire SB_20_n13 ;
    wire SB_20_n12 ;
    wire SB_20_n11 ;
    wire SB_20_n10 ;
    wire SB_20_n9 ;
    wire SB_20_T5 ;
    wire SB_20_T4 ;
    wire SB_20_T3 ;
    wire SB_20_T2 ;
    wire SB_20_T1 ;
    wire SB_20_T0 ;
    wire SB_19_n15 ;
    wire SB_19_n14 ;
    wire SB_19_n13 ;
    wire SB_19_n12 ;
    wire SB_19_n11 ;
    wire SB_19_n10 ;
    wire SB_19_n9 ;
    wire SB_19_T5 ;
    wire SB_19_T4 ;
    wire SB_19_T3 ;
    wire SB_19_T2 ;
    wire SB_19_T1 ;
    wire SB_19_T0 ;
    wire SB_18_n15 ;
    wire SB_18_n14 ;
    wire SB_18_n13 ;
    wire SB_18_n12 ;
    wire SB_18_n11 ;
    wire SB_18_n10 ;
    wire SB_18_n9 ;
    wire SB_18_T5 ;
    wire SB_18_T4 ;
    wire SB_18_T3 ;
    wire SB_18_T2 ;
    wire SB_18_T1 ;
    wire SB_18_T0 ;
    wire SB_17_n15 ;
    wire SB_17_n14 ;
    wire SB_17_n13 ;
    wire SB_17_n12 ;
    wire SB_17_n11 ;
    wire SB_17_n10 ;
    wire SB_17_n9 ;
    wire SB_17_T5 ;
    wire SB_17_T4 ;
    wire SB_17_T3 ;
    wire SB_17_T2 ;
    wire SB_17_T1 ;
    wire SB_17_T0 ;
    wire SB_16_n15 ;
    wire SB_16_n14 ;
    wire SB_16_n13 ;
    wire SB_16_n12 ;
    wire SB_16_n11 ;
    wire SB_16_n10 ;
    wire SB_16_n9 ;
    wire SB_16_T5 ;
    wire SB_16_T4 ;
    wire SB_16_T3 ;
    wire SB_16_T2 ;
    wire SB_16_T1 ;
    wire SB_16_T0 ;
    wire SB_15_n15 ;
    wire SB_15_n14 ;
    wire SB_15_n13 ;
    wire SB_15_n12 ;
    wire SB_15_n11 ;
    wire SB_15_n10 ;
    wire SB_15_n9 ;
    wire SB_15_T5 ;
    wire SB_15_T4 ;
    wire SB_15_T3 ;
    wire SB_15_T2 ;
    wire SB_15_T1 ;
    wire SB_15_T0 ;
    wire SB_14_n15 ;
    wire SB_14_n14 ;
    wire SB_14_n13 ;
    wire SB_14_n12 ;
    wire SB_14_n11 ;
    wire SB_14_n10 ;
    wire SB_14_n9 ;
    wire SB_14_T5 ;
    wire SB_14_T4 ;
    wire SB_14_T3 ;
    wire SB_14_T2 ;
    wire SB_14_T1 ;
    wire SB_14_T0 ;
    wire SB_13_n15 ;
    wire SB_13_n14 ;
    wire SB_13_n13 ;
    wire SB_13_n12 ;
    wire SB_13_n11 ;
    wire SB_13_n10 ;
    wire SB_13_n9 ;
    wire SB_13_T5 ;
    wire SB_13_T4 ;
    wire SB_13_T3 ;
    wire SB_13_T2 ;
    wire SB_13_T1 ;
    wire SB_13_T0 ;
    wire SB_12_n15 ;
    wire SB_12_n14 ;
    wire SB_12_n13 ;
    wire SB_12_n12 ;
    wire SB_12_n11 ;
    wire SB_12_n10 ;
    wire SB_12_n9 ;
    wire SB_12_T5 ;
    wire SB_12_T4 ;
    wire SB_12_T3 ;
    wire SB_12_T2 ;
    wire SB_12_T1 ;
    wire SB_12_T0 ;
    wire SB_11_n15 ;
    wire SB_11_n14 ;
    wire SB_11_n13 ;
    wire SB_11_n12 ;
    wire SB_11_n11 ;
    wire SB_11_n10 ;
    wire SB_11_n9 ;
    wire SB_11_T5 ;
    wire SB_11_T4 ;
    wire SB_11_T3 ;
    wire SB_11_T2 ;
    wire SB_11_T1 ;
    wire SB_11_T0 ;
    wire SB_10_n15 ;
    wire SB_10_n14 ;
    wire SB_10_n13 ;
    wire SB_10_n12 ;
    wire SB_10_n11 ;
    wire SB_10_n10 ;
    wire SB_10_n9 ;
    wire SB_10_T5 ;
    wire SB_10_T4 ;
    wire SB_10_T3 ;
    wire SB_10_T2 ;
    wire SB_10_T1 ;
    wire SB_10_T0 ;
    wire SB_9_n15 ;
    wire SB_9_n14 ;
    wire SB_9_n13 ;
    wire SB_9_n12 ;
    wire SB_9_n11 ;
    wire SB_9_n10 ;
    wire SB_9_n9 ;
    wire SB_9_T5 ;
    wire SB_9_T4 ;
    wire SB_9_T3 ;
    wire SB_9_T2 ;
    wire SB_9_T1 ;
    wire SB_9_T0 ;
    wire SB_8_n15 ;
    wire SB_8_n14 ;
    wire SB_8_n13 ;
    wire SB_8_n12 ;
    wire SB_8_n11 ;
    wire SB_8_n10 ;
    wire SB_8_n9 ;
    wire SB_8_T5 ;
    wire SB_8_T4 ;
    wire SB_8_T3 ;
    wire SB_8_T2 ;
    wire SB_8_T1 ;
    wire SB_8_T0 ;
    wire SB_7_n15 ;
    wire SB_7_n14 ;
    wire SB_7_n13 ;
    wire SB_7_n12 ;
    wire SB_7_n11 ;
    wire SB_7_n10 ;
    wire SB_7_n9 ;
    wire SB_7_T5 ;
    wire SB_7_T4 ;
    wire SB_7_T3 ;
    wire SB_7_T2 ;
    wire SB_7_T1 ;
    wire SB_7_T0 ;
    wire SB_6_n15 ;
    wire SB_6_n14 ;
    wire SB_6_n13 ;
    wire SB_6_n12 ;
    wire SB_6_n11 ;
    wire SB_6_n10 ;
    wire SB_6_n9 ;
    wire SB_6_T5 ;
    wire SB_6_T4 ;
    wire SB_6_T3 ;
    wire SB_6_T2 ;
    wire SB_6_T1 ;
    wire SB_6_T0 ;
    wire SB_5_n15 ;
    wire SB_5_n14 ;
    wire SB_5_n13 ;
    wire SB_5_n12 ;
    wire SB_5_n11 ;
    wire SB_5_n10 ;
    wire SB_5_n9 ;
    wire SB_5_T5 ;
    wire SB_5_T4 ;
    wire SB_5_T3 ;
    wire SB_5_T2 ;
    wire SB_5_T1 ;
    wire SB_5_T0 ;
    wire SB_4_n15 ;
    wire SB_4_n14 ;
    wire SB_4_n13 ;
    wire SB_4_n12 ;
    wire SB_4_n11 ;
    wire SB_4_n10 ;
    wire SB_4_n9 ;
    wire SB_4_T5 ;
    wire SB_4_T4 ;
    wire SB_4_T3 ;
    wire SB_4_T2 ;
    wire SB_4_T1 ;
    wire SB_4_T0 ;
    wire SB_3_n15 ;
    wire SB_3_n14 ;
    wire SB_3_n13 ;
    wire SB_3_n12 ;
    wire SB_3_n11 ;
    wire SB_3_n10 ;
    wire SB_3_n9 ;
    wire SB_3_T5 ;
    wire SB_3_T4 ;
    wire SB_3_T3 ;
    wire SB_3_T2 ;
    wire SB_3_T1 ;
    wire SB_3_T0 ;
    wire SB_2_n15 ;
    wire SB_2_n14 ;
    wire SB_2_n13 ;
    wire SB_2_n12 ;
    wire SB_2_n11 ;
    wire SB_2_n10 ;
    wire SB_2_n9 ;
    wire SB_2_T5 ;
    wire SB_2_T4 ;
    wire SB_2_T3 ;
    wire SB_2_T2 ;
    wire SB_2_T1 ;
    wire SB_2_T0 ;
    wire SB_1_n15 ;
    wire SB_1_n14 ;
    wire SB_1_n13 ;
    wire SB_1_n12 ;
    wire SB_1_n11 ;
    wire SB_1_n10 ;
    wire SB_1_n9 ;
    wire SB_1_T5 ;
    wire SB_1_T4 ;
    wire SB_1_T3 ;
    wire SB_1_T2 ;
    wire SB_1_T1 ;
    wire SB_1_T0 ;
    wire SB_0_n15 ;
    wire SB_0_n14 ;
    wire SB_0_n13 ;
    wire SB_0_n12 ;
    wire SB_0_n11 ;
    wire SB_0_n10 ;
    wire SB_0_n9 ;
    wire SB_0_T5 ;
    wire SB_0_T4 ;
    wire SB_0_T3 ;
    wire SB_0_T2 ;
    wire SB_0_T1 ;
    wire SB_0_T0 ;
    wire new_AGEMA_signal_683 ;
    wire new_AGEMA_signal_684 ;
    wire new_AGEMA_signal_689 ;
    wire new_AGEMA_signal_690 ;
    wire new_AGEMA_signal_691 ;
    wire new_AGEMA_signal_692 ;
    wire new_AGEMA_signal_693 ;
    wire new_AGEMA_signal_694 ;
    wire new_AGEMA_signal_695 ;
    wire new_AGEMA_signal_696 ;
    wire new_AGEMA_signal_697 ;
    wire new_AGEMA_signal_698 ;
    wire new_AGEMA_signal_703 ;
    wire new_AGEMA_signal_704 ;
    wire new_AGEMA_signal_709 ;
    wire new_AGEMA_signal_710 ;
    wire new_AGEMA_signal_711 ;
    wire new_AGEMA_signal_712 ;
    wire new_AGEMA_signal_713 ;
    wire new_AGEMA_signal_714 ;
    wire new_AGEMA_signal_715 ;
    wire new_AGEMA_signal_716 ;
    wire new_AGEMA_signal_717 ;
    wire new_AGEMA_signal_718 ;
    wire new_AGEMA_signal_723 ;
    wire new_AGEMA_signal_724 ;
    wire new_AGEMA_signal_729 ;
    wire new_AGEMA_signal_730 ;
    wire new_AGEMA_signal_731 ;
    wire new_AGEMA_signal_732 ;
    wire new_AGEMA_signal_733 ;
    wire new_AGEMA_signal_734 ;
    wire new_AGEMA_signal_735 ;
    wire new_AGEMA_signal_736 ;
    wire new_AGEMA_signal_737 ;
    wire new_AGEMA_signal_738 ;
    wire new_AGEMA_signal_743 ;
    wire new_AGEMA_signal_744 ;
    wire new_AGEMA_signal_749 ;
    wire new_AGEMA_signal_750 ;
    wire new_AGEMA_signal_751 ;
    wire new_AGEMA_signal_752 ;
    wire new_AGEMA_signal_753 ;
    wire new_AGEMA_signal_754 ;
    wire new_AGEMA_signal_755 ;
    wire new_AGEMA_signal_756 ;
    wire new_AGEMA_signal_757 ;
    wire new_AGEMA_signal_758 ;
    wire new_AGEMA_signal_763 ;
    wire new_AGEMA_signal_764 ;
    wire new_AGEMA_signal_769 ;
    wire new_AGEMA_signal_770 ;
    wire new_AGEMA_signal_771 ;
    wire new_AGEMA_signal_772 ;
    wire new_AGEMA_signal_773 ;
    wire new_AGEMA_signal_774 ;
    wire new_AGEMA_signal_775 ;
    wire new_AGEMA_signal_776 ;
    wire new_AGEMA_signal_777 ;
    wire new_AGEMA_signal_778 ;
    wire new_AGEMA_signal_783 ;
    wire new_AGEMA_signal_784 ;
    wire new_AGEMA_signal_789 ;
    wire new_AGEMA_signal_790 ;
    wire new_AGEMA_signal_791 ;
    wire new_AGEMA_signal_792 ;
    wire new_AGEMA_signal_793 ;
    wire new_AGEMA_signal_794 ;
    wire new_AGEMA_signal_795 ;
    wire new_AGEMA_signal_796 ;
    wire new_AGEMA_signal_797 ;
    wire new_AGEMA_signal_798 ;
    wire new_AGEMA_signal_803 ;
    wire new_AGEMA_signal_804 ;
    wire new_AGEMA_signal_809 ;
    wire new_AGEMA_signal_810 ;
    wire new_AGEMA_signal_811 ;
    wire new_AGEMA_signal_812 ;
    wire new_AGEMA_signal_813 ;
    wire new_AGEMA_signal_814 ;
    wire new_AGEMA_signal_815 ;
    wire new_AGEMA_signal_816 ;
    wire new_AGEMA_signal_817 ;
    wire new_AGEMA_signal_818 ;
    wire new_AGEMA_signal_823 ;
    wire new_AGEMA_signal_824 ;
    wire new_AGEMA_signal_829 ;
    wire new_AGEMA_signal_830 ;
    wire new_AGEMA_signal_831 ;
    wire new_AGEMA_signal_832 ;
    wire new_AGEMA_signal_833 ;
    wire new_AGEMA_signal_834 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_836 ;
    wire new_AGEMA_signal_837 ;
    wire new_AGEMA_signal_838 ;
    wire new_AGEMA_signal_843 ;
    wire new_AGEMA_signal_844 ;
    wire new_AGEMA_signal_849 ;
    wire new_AGEMA_signal_850 ;
    wire new_AGEMA_signal_851 ;
    wire new_AGEMA_signal_852 ;
    wire new_AGEMA_signal_853 ;
    wire new_AGEMA_signal_854 ;
    wire new_AGEMA_signal_855 ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_857 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_863 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_869 ;
    wire new_AGEMA_signal_870 ;
    wire new_AGEMA_signal_871 ;
    wire new_AGEMA_signal_872 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_874 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_878 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_890 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_892 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_896 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_898 ;
    wire new_AGEMA_signal_903 ;
    wire new_AGEMA_signal_904 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_910 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_912 ;
    wire new_AGEMA_signal_913 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_915 ;
    wire new_AGEMA_signal_916 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_924 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_930 ;
    wire new_AGEMA_signal_931 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_934 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U8 ( .a ({SubC_in_s2[63], SubC_in_s1[63], SubC_in_s0[63]}), .b ({SubC_in_s2[95], SubC_in_s1[95], SubC_in_s0[95]}), .c ({new_AGEMA_signal_684, new_AGEMA_signal_683, SB_31_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U3 ( .a ({SubC_in_s2[31], SubC_in_s1[31], SubC_in_s0[31]}), .b ({SubC_in_s2[127], SubC_in_s1[127], SubC_in_s0[127]}), .c ({new_AGEMA_signal_690, new_AGEMA_signal_689, SB_31_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U8 ( .a ({SubC_in_s2[62], SubC_in_s1[62], SubC_in_s0[62]}), .b ({SubC_in_s2[94], SubC_in_s1[94], SubC_in_s0[94]}), .c ({new_AGEMA_signal_704, new_AGEMA_signal_703, SB_30_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U3 ( .a ({SubC_in_s2[30], SubC_in_s1[30], SubC_in_s0[30]}), .b ({SubC_in_s2[126], SubC_in_s1[126], SubC_in_s0[126]}), .c ({new_AGEMA_signal_710, new_AGEMA_signal_709, SB_30_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U8 ( .a ({SubC_in_s2[61], SubC_in_s1[61], SubC_in_s0[61]}), .b ({SubC_in_s2[93], SubC_in_s1[93], SubC_in_s0[93]}), .c ({new_AGEMA_signal_724, new_AGEMA_signal_723, SB_29_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U3 ( .a ({SubC_in_s2[29], SubC_in_s1[29], SubC_in_s0[29]}), .b ({SubC_in_s2[125], SubC_in_s1[125], SubC_in_s0[125]}), .c ({new_AGEMA_signal_730, new_AGEMA_signal_729, SB_29_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U8 ( .a ({SubC_in_s2[60], SubC_in_s1[60], SubC_in_s0[60]}), .b ({SubC_in_s2[92], SubC_in_s1[92], SubC_in_s0[92]}), .c ({new_AGEMA_signal_744, new_AGEMA_signal_743, SB_28_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U3 ( .a ({SubC_in_s2[28], SubC_in_s1[28], SubC_in_s0[28]}), .b ({SubC_in_s2[124], SubC_in_s1[124], SubC_in_s0[124]}), .c ({new_AGEMA_signal_750, new_AGEMA_signal_749, SB_28_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U8 ( .a ({SubC_in_s2[59], SubC_in_s1[59], SubC_in_s0[59]}), .b ({SubC_in_s2[91], SubC_in_s1[91], SubC_in_s0[91]}), .c ({new_AGEMA_signal_764, new_AGEMA_signal_763, SB_27_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U3 ( .a ({SubC_in_s2[27], SubC_in_s1[27], SubC_in_s0[27]}), .b ({SubC_in_s2[123], SubC_in_s1[123], SubC_in_s0[123]}), .c ({new_AGEMA_signal_770, new_AGEMA_signal_769, SB_27_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U8 ( .a ({SubC_in_s2[58], SubC_in_s1[58], SubC_in_s0[58]}), .b ({SubC_in_s2[90], SubC_in_s1[90], SubC_in_s0[90]}), .c ({new_AGEMA_signal_784, new_AGEMA_signal_783, SB_26_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U3 ( .a ({SubC_in_s2[26], SubC_in_s1[26], SubC_in_s0[26]}), .b ({SubC_in_s2[122], SubC_in_s1[122], SubC_in_s0[122]}), .c ({new_AGEMA_signal_790, new_AGEMA_signal_789, SB_26_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U8 ( .a ({SubC_in_s2[57], SubC_in_s1[57], SubC_in_s0[57]}), .b ({SubC_in_s2[89], SubC_in_s1[89], SubC_in_s0[89]}), .c ({new_AGEMA_signal_804, new_AGEMA_signal_803, SB_25_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U3 ( .a ({SubC_in_s2[25], SubC_in_s1[25], SubC_in_s0[25]}), .b ({SubC_in_s2[121], SubC_in_s1[121], SubC_in_s0[121]}), .c ({new_AGEMA_signal_810, new_AGEMA_signal_809, SB_25_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U8 ( .a ({SubC_in_s2[56], SubC_in_s1[56], SubC_in_s0[56]}), .b ({SubC_in_s2[88], SubC_in_s1[88], SubC_in_s0[88]}), .c ({new_AGEMA_signal_824, new_AGEMA_signal_823, SB_24_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U3 ( .a ({SubC_in_s2[24], SubC_in_s1[24], SubC_in_s0[24]}), .b ({SubC_in_s2[120], SubC_in_s1[120], SubC_in_s0[120]}), .c ({new_AGEMA_signal_830, new_AGEMA_signal_829, SB_24_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U8 ( .a ({SubC_in_s2[55], SubC_in_s1[55], SubC_in_s0[55]}), .b ({SubC_in_s2[87], SubC_in_s1[87], SubC_in_s0[87]}), .c ({new_AGEMA_signal_844, new_AGEMA_signal_843, SB_23_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U3 ( .a ({SubC_in_s2[23], SubC_in_s1[23], SubC_in_s0[23]}), .b ({SubC_in_s2[119], SubC_in_s1[119], SubC_in_s0[119]}), .c ({new_AGEMA_signal_850, new_AGEMA_signal_849, SB_23_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U8 ( .a ({SubC_in_s2[54], SubC_in_s1[54], SubC_in_s0[54]}), .b ({SubC_in_s2[86], SubC_in_s1[86], SubC_in_s0[86]}), .c ({new_AGEMA_signal_864, new_AGEMA_signal_863, SB_22_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U3 ( .a ({SubC_in_s2[22], SubC_in_s1[22], SubC_in_s0[22]}), .b ({SubC_in_s2[118], SubC_in_s1[118], SubC_in_s0[118]}), .c ({new_AGEMA_signal_870, new_AGEMA_signal_869, SB_22_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U8 ( .a ({SubC_in_s2[53], SubC_in_s1[53], SubC_in_s0[53]}), .b ({SubC_in_s2[85], SubC_in_s1[85], SubC_in_s0[85]}), .c ({new_AGEMA_signal_884, new_AGEMA_signal_883, SB_21_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U3 ( .a ({SubC_in_s2[21], SubC_in_s1[21], SubC_in_s0[21]}), .b ({SubC_in_s2[117], SubC_in_s1[117], SubC_in_s0[117]}), .c ({new_AGEMA_signal_890, new_AGEMA_signal_889, SB_21_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U8 ( .a ({SubC_in_s2[52], SubC_in_s1[52], SubC_in_s0[52]}), .b ({SubC_in_s2[84], SubC_in_s1[84], SubC_in_s0[84]}), .c ({new_AGEMA_signal_904, new_AGEMA_signal_903, SB_20_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U3 ( .a ({SubC_in_s2[20], SubC_in_s1[20], SubC_in_s0[20]}), .b ({SubC_in_s2[116], SubC_in_s1[116], SubC_in_s0[116]}), .c ({new_AGEMA_signal_910, new_AGEMA_signal_909, SB_20_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U8 ( .a ({SubC_in_s2[51], SubC_in_s1[51], SubC_in_s0[51]}), .b ({SubC_in_s2[83], SubC_in_s1[83], SubC_in_s0[83]}), .c ({new_AGEMA_signal_924, new_AGEMA_signal_923, SB_19_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U3 ( .a ({SubC_in_s2[19], SubC_in_s1[19], SubC_in_s0[19]}), .b ({SubC_in_s2[115], SubC_in_s1[115], SubC_in_s0[115]}), .c ({new_AGEMA_signal_930, new_AGEMA_signal_929, SB_19_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U8 ( .a ({SubC_in_s2[50], SubC_in_s1[50], SubC_in_s0[50]}), .b ({SubC_in_s2[82], SubC_in_s1[82], SubC_in_s0[82]}), .c ({new_AGEMA_signal_944, new_AGEMA_signal_943, SB_18_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U3 ( .a ({SubC_in_s2[18], SubC_in_s1[18], SubC_in_s0[18]}), .b ({SubC_in_s2[114], SubC_in_s1[114], SubC_in_s0[114]}), .c ({new_AGEMA_signal_950, new_AGEMA_signal_949, SB_18_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U8 ( .a ({SubC_in_s2[49], SubC_in_s1[49], SubC_in_s0[49]}), .b ({SubC_in_s2[81], SubC_in_s1[81], SubC_in_s0[81]}), .c ({new_AGEMA_signal_964, new_AGEMA_signal_963, SB_17_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U3 ( .a ({SubC_in_s2[17], SubC_in_s1[17], SubC_in_s0[17]}), .b ({SubC_in_s2[113], SubC_in_s1[113], SubC_in_s0[113]}), .c ({new_AGEMA_signal_970, new_AGEMA_signal_969, SB_17_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U8 ( .a ({SubC_in_s2[48], SubC_in_s1[48], SubC_in_s0[48]}), .b ({SubC_in_s2[80], SubC_in_s1[80], SubC_in_s0[80]}), .c ({new_AGEMA_signal_984, new_AGEMA_signal_983, SB_16_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U3 ( .a ({SubC_in_s2[16], SubC_in_s1[16], SubC_in_s0[16]}), .b ({SubC_in_s2[112], SubC_in_s1[112], SubC_in_s0[112]}), .c ({new_AGEMA_signal_990, new_AGEMA_signal_989, SB_16_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U8 ( .a ({SubC_in_s2[47], SubC_in_s1[47], SubC_in_s0[47]}), .b ({SubC_in_s2[79], SubC_in_s1[79], SubC_in_s0[79]}), .c ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, SB_15_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U3 ( .a ({SubC_in_s2[15], SubC_in_s1[15], SubC_in_s0[15]}), .b ({SubC_in_s2[111], SubC_in_s1[111], SubC_in_s0[111]}), .c ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, SB_15_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U8 ( .a ({SubC_in_s2[46], SubC_in_s1[46], SubC_in_s0[46]}), .b ({SubC_in_s2[78], SubC_in_s1[78], SubC_in_s0[78]}), .c ({new_AGEMA_signal_1024, new_AGEMA_signal_1023, SB_14_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U3 ( .a ({SubC_in_s2[14], SubC_in_s1[14], SubC_in_s0[14]}), .b ({SubC_in_s2[110], SubC_in_s1[110], SubC_in_s0[110]}), .c ({new_AGEMA_signal_1030, new_AGEMA_signal_1029, SB_14_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U8 ( .a ({SubC_in_s2[45], SubC_in_s1[45], SubC_in_s0[45]}), .b ({SubC_in_s2[77], SubC_in_s1[77], SubC_in_s0[77]}), .c ({new_AGEMA_signal_1044, new_AGEMA_signal_1043, SB_13_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U3 ( .a ({SubC_in_s2[13], SubC_in_s1[13], SubC_in_s0[13]}), .b ({SubC_in_s2[109], SubC_in_s1[109], SubC_in_s0[109]}), .c ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SB_13_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U8 ( .a ({SubC_in_s2[44], SubC_in_s1[44], SubC_in_s0[44]}), .b ({SubC_in_s2[76], SubC_in_s1[76], SubC_in_s0[76]}), .c ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SB_12_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U3 ( .a ({SubC_in_s2[12], SubC_in_s1[12], SubC_in_s0[12]}), .b ({SubC_in_s2[108], SubC_in_s1[108], SubC_in_s0[108]}), .c ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, SB_12_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U8 ( .a ({SubC_in_s2[43], SubC_in_s1[43], SubC_in_s0[43]}), .b ({SubC_in_s2[75], SubC_in_s1[75], SubC_in_s0[75]}), .c ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, SB_11_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U3 ( .a ({SubC_in_s2[11], SubC_in_s1[11], SubC_in_s0[11]}), .b ({SubC_in_s2[107], SubC_in_s1[107], SubC_in_s0[107]}), .c ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, SB_11_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U8 ( .a ({SubC_in_s2[42], SubC_in_s1[42], SubC_in_s0[42]}), .b ({SubC_in_s2[74], SubC_in_s1[74], SubC_in_s0[74]}), .c ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, SB_10_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U3 ( .a ({SubC_in_s2[10], SubC_in_s1[10], SubC_in_s0[10]}), .b ({SubC_in_s2[106], SubC_in_s1[106], SubC_in_s0[106]}), .c ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, SB_10_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U8 ( .a ({SubC_in_s2[41], SubC_in_s1[41], SubC_in_s0[41]}), .b ({SubC_in_s2[73], SubC_in_s1[73], SubC_in_s0[73]}), .c ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, SB_9_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U3 ( .a ({SubC_in_s2[9], SubC_in_s1[9], SubC_in_s0[9]}), .b ({SubC_in_s2[105], SubC_in_s1[105], SubC_in_s0[105]}), .c ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SB_9_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U8 ( .a ({SubC_in_s2[40], SubC_in_s1[40], SubC_in_s0[40]}), .b ({SubC_in_s2[72], SubC_in_s1[72], SubC_in_s0[72]}), .c ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SB_8_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U3 ( .a ({SubC_in_s2[8], SubC_in_s1[8], SubC_in_s0[8]}), .b ({SubC_in_s2[104], SubC_in_s1[104], SubC_in_s0[104]}), .c ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, SB_8_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U8 ( .a ({SubC_in_s2[39], SubC_in_s1[39], SubC_in_s0[39]}), .b ({SubC_in_s2[71], SubC_in_s1[71], SubC_in_s0[71]}), .c ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, SB_7_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U3 ( .a ({SubC_in_s2[7], SubC_in_s1[7], SubC_in_s0[7]}), .b ({SubC_in_s2[103], SubC_in_s1[103], SubC_in_s0[103]}), .c ({new_AGEMA_signal_1170, new_AGEMA_signal_1169, SB_7_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U8 ( .a ({SubC_in_s2[38], SubC_in_s1[38], SubC_in_s0[38]}), .b ({SubC_in_s2[70], SubC_in_s1[70], SubC_in_s0[70]}), .c ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, SB_6_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U3 ( .a ({SubC_in_s2[6], SubC_in_s1[6], SubC_in_s0[6]}), .b ({SubC_in_s2[102], SubC_in_s1[102], SubC_in_s0[102]}), .c ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, SB_6_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U8 ( .a ({SubC_in_s2[37], SubC_in_s1[37], SubC_in_s0[37]}), .b ({SubC_in_s2[69], SubC_in_s1[69], SubC_in_s0[69]}), .c ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, SB_5_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U3 ( .a ({SubC_in_s2[5], SubC_in_s1[5], SubC_in_s0[5]}), .b ({SubC_in_s2[101], SubC_in_s1[101], SubC_in_s0[101]}), .c ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SB_5_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U8 ( .a ({SubC_in_s2[36], SubC_in_s1[36], SubC_in_s0[36]}), .b ({SubC_in_s2[68], SubC_in_s1[68], SubC_in_s0[68]}), .c ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SB_4_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U3 ( .a ({SubC_in_s2[4], SubC_in_s1[4], SubC_in_s0[4]}), .b ({SubC_in_s2[100], SubC_in_s1[100], SubC_in_s0[100]}), .c ({new_AGEMA_signal_1230, new_AGEMA_signal_1229, SB_4_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U8 ( .a ({SubC_in_s2[35], SubC_in_s1[35], SubC_in_s0[35]}), .b ({SubC_in_s2[67], SubC_in_s1[67], SubC_in_s0[67]}), .c ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, SB_3_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U3 ( .a ({SubC_in_s2[3], SubC_in_s1[3], SubC_in_s0[3]}), .b ({SubC_in_s2[99], SubC_in_s1[99], SubC_in_s0[99]}), .c ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, SB_3_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U8 ( .a ({SubC_in_s2[34], SubC_in_s1[34], SubC_in_s0[34]}), .b ({SubC_in_s2[66], SubC_in_s1[66], SubC_in_s0[66]}), .c ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, SB_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U3 ( .a ({SubC_in_s2[2], SubC_in_s1[2], SubC_in_s0[2]}), .b ({SubC_in_s2[98], SubC_in_s1[98], SubC_in_s0[98]}), .c ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, SB_2_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U8 ( .a ({SubC_in_s2[33], SubC_in_s1[33], SubC_in_s0[33]}), .b ({SubC_in_s2[65], SubC_in_s1[65], SubC_in_s0[65]}), .c ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, SB_1_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U3 ( .a ({SubC_in_s2[1], SubC_in_s1[1], SubC_in_s0[1]}), .b ({SubC_in_s2[97], SubC_in_s1[97], SubC_in_s0[97]}), .c ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, SB_1_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U8 ( .a ({SubC_in_s2[32], SubC_in_s1[32], SubC_in_s0[32]}), .b ({SubC_in_s2[64], SubC_in_s1[64], SubC_in_s0[64]}), .c ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, SB_0_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U3 ( .a ({SubC_in_s2[0], SubC_in_s1[0], SubC_in_s0[0]}), .b ({SubC_in_s2[96], SubC_in_s1[96], SubC_in_s0[96]}), .c ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, SB_0_n10}) ) ;
    //ClockGatingController #(4) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U11 ( .a ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, SB_31_n15}), .b ({new_AGEMA_signal_684, new_AGEMA_signal_683, SB_31_n14}), .c ({SubC_out_s2[127], SubC_out_s1[127], SubC_out_s0[127]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U9 ( .a ({new_AGEMA_signal_684, new_AGEMA_signal_683, SB_31_n14}), .b ({new_AGEMA_signal_696, new_AGEMA_signal_695, SB_31_T2}), .c ({new_AGEMA_signal_1320, new_AGEMA_signal_1319, SB_31_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U6 ( .a ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, SB_31_n11}), .b ({new_AGEMA_signal_694, new_AGEMA_signal_693, SB_31_T1}), .c ({SubC_out_s2[95], SubC_out_s1[95], SubC_out_s0[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U5 ( .a ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, SB_31_n15}), .b ({SubC_in_s2[63], SubC_in_s1[63], SubC_in_s0[63]}), .c ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, SB_31_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U4 ( .a ({new_AGEMA_signal_690, new_AGEMA_signal_689, SB_31_n10}), .b ({new_AGEMA_signal_692, new_AGEMA_signal_691, SB_31_T0}), .c ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, SB_31_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U1 ( .a ({SubC_in_s2[127], SubC_in_s1[127], SubC_in_s0[127]}), .b ({new_AGEMA_signal_698, new_AGEMA_signal_697, SB_31_T3}), .c ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, SB_31_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_31_t0_AND_U1 ( .a ({SubC_in_s2[127], SubC_in_s1[127], SubC_in_s0[127]}), .b ({SubC_in_s2[95], SubC_in_s1[95], SubC_in_s0[95]}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_692, new_AGEMA_signal_691, SB_31_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_31_t1_AND_U1 ( .a ({SubC_in_s2[127], SubC_in_s1[127], SubC_in_s0[127]}), .b ({SubC_in_s2[63], SubC_in_s1[63], SubC_in_s0[63]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_694, new_AGEMA_signal_693, SB_31_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_31_t2_AND_U1 ( .a ({SubC_in_s2[127], SubC_in_s1[127], SubC_in_s0[127]}), .b ({SubC_in_s2[31], SubC_in_s1[31], SubC_in_s0[31]}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_696, new_AGEMA_signal_695, SB_31_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_31_t3_AND_U1 ( .a ({SubC_in_s2[95], SubC_in_s1[95], SubC_in_s0[95]}), .b ({SubC_in_s2[31], SubC_in_s1[31], SubC_in_s0[31]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_698, new_AGEMA_signal_697, SB_31_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U11 ( .a ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, SB_30_n15}), .b ({new_AGEMA_signal_704, new_AGEMA_signal_703, SB_30_n14}), .c ({SubC_out_s2[126], SubC_out_s1[126], SubC_out_s0[126]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U9 ( .a ({new_AGEMA_signal_704, new_AGEMA_signal_703, SB_30_n14}), .b ({new_AGEMA_signal_716, new_AGEMA_signal_715, SB_30_T2}), .c ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, SB_30_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U6 ( .a ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, SB_30_n11}), .b ({new_AGEMA_signal_714, new_AGEMA_signal_713, SB_30_T1}), .c ({SubC_out_s2[94], SubC_out_s1[94], SubC_out_s0[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U5 ( .a ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, SB_30_n15}), .b ({SubC_in_s2[62], SubC_in_s1[62], SubC_in_s0[62]}), .c ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, SB_30_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U4 ( .a ({new_AGEMA_signal_710, new_AGEMA_signal_709, SB_30_n10}), .b ({new_AGEMA_signal_712, new_AGEMA_signal_711, SB_30_T0}), .c ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, SB_30_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U1 ( .a ({SubC_in_s2[126], SubC_in_s1[126], SubC_in_s0[126]}), .b ({new_AGEMA_signal_718, new_AGEMA_signal_717, SB_30_T3}), .c ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, SB_30_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_30_t0_AND_U1 ( .a ({SubC_in_s2[126], SubC_in_s1[126], SubC_in_s0[126]}), .b ({SubC_in_s2[94], SubC_in_s1[94], SubC_in_s0[94]}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_712, new_AGEMA_signal_711, SB_30_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_30_t1_AND_U1 ( .a ({SubC_in_s2[126], SubC_in_s1[126], SubC_in_s0[126]}), .b ({SubC_in_s2[62], SubC_in_s1[62], SubC_in_s0[62]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_714, new_AGEMA_signal_713, SB_30_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_30_t2_AND_U1 ( .a ({SubC_in_s2[126], SubC_in_s1[126], SubC_in_s0[126]}), .b ({SubC_in_s2[30], SubC_in_s1[30], SubC_in_s0[30]}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_716, new_AGEMA_signal_715, SB_30_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_30_t3_AND_U1 ( .a ({SubC_in_s2[94], SubC_in_s1[94], SubC_in_s0[94]}), .b ({SubC_in_s2[30], SubC_in_s1[30], SubC_in_s0[30]}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_718, new_AGEMA_signal_717, SB_30_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U11 ( .a ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, SB_29_n15}), .b ({new_AGEMA_signal_724, new_AGEMA_signal_723, SB_29_n14}), .c ({SubC_out_s2[125], SubC_out_s1[125], SubC_out_s0[125]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U9 ( .a ({new_AGEMA_signal_724, new_AGEMA_signal_723, SB_29_n14}), .b ({new_AGEMA_signal_736, new_AGEMA_signal_735, SB_29_T2}), .c ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, SB_29_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U6 ( .a ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, SB_29_n11}), .b ({new_AGEMA_signal_734, new_AGEMA_signal_733, SB_29_T1}), .c ({SubC_out_s2[93], SubC_out_s1[93], SubC_out_s0[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U5 ( .a ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, SB_29_n15}), .b ({SubC_in_s2[61], SubC_in_s1[61], SubC_in_s0[61]}), .c ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, SB_29_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U4 ( .a ({new_AGEMA_signal_730, new_AGEMA_signal_729, SB_29_n10}), .b ({new_AGEMA_signal_732, new_AGEMA_signal_731, SB_29_T0}), .c ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, SB_29_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U1 ( .a ({SubC_in_s2[125], SubC_in_s1[125], SubC_in_s0[125]}), .b ({new_AGEMA_signal_738, new_AGEMA_signal_737, SB_29_T3}), .c ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, SB_29_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_29_t0_AND_U1 ( .a ({SubC_in_s2[125], SubC_in_s1[125], SubC_in_s0[125]}), .b ({SubC_in_s2[93], SubC_in_s1[93], SubC_in_s0[93]}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_732, new_AGEMA_signal_731, SB_29_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_29_t1_AND_U1 ( .a ({SubC_in_s2[125], SubC_in_s1[125], SubC_in_s0[125]}), .b ({SubC_in_s2[61], SubC_in_s1[61], SubC_in_s0[61]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_734, new_AGEMA_signal_733, SB_29_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_29_t2_AND_U1 ( .a ({SubC_in_s2[125], SubC_in_s1[125], SubC_in_s0[125]}), .b ({SubC_in_s2[29], SubC_in_s1[29], SubC_in_s0[29]}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_736, new_AGEMA_signal_735, SB_29_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_29_t3_AND_U1 ( .a ({SubC_in_s2[93], SubC_in_s1[93], SubC_in_s0[93]}), .b ({SubC_in_s2[29], SubC_in_s1[29], SubC_in_s0[29]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_738, new_AGEMA_signal_737, SB_29_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U11 ( .a ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, SB_28_n15}), .b ({new_AGEMA_signal_744, new_AGEMA_signal_743, SB_28_n14}), .c ({SubC_out_s2[124], SubC_out_s1[124], SubC_out_s0[124]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U9 ( .a ({new_AGEMA_signal_744, new_AGEMA_signal_743, SB_28_n14}), .b ({new_AGEMA_signal_756, new_AGEMA_signal_755, SB_28_T2}), .c ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, SB_28_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U6 ( .a ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, SB_28_n11}), .b ({new_AGEMA_signal_754, new_AGEMA_signal_753, SB_28_T1}), .c ({SubC_out_s2[92], SubC_out_s1[92], SubC_out_s0[92]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U5 ( .a ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, SB_28_n15}), .b ({SubC_in_s2[60], SubC_in_s1[60], SubC_in_s0[60]}), .c ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, SB_28_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U4 ( .a ({new_AGEMA_signal_750, new_AGEMA_signal_749, SB_28_n10}), .b ({new_AGEMA_signal_752, new_AGEMA_signal_751, SB_28_T0}), .c ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, SB_28_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U1 ( .a ({SubC_in_s2[124], SubC_in_s1[124], SubC_in_s0[124]}), .b ({new_AGEMA_signal_758, new_AGEMA_signal_757, SB_28_T3}), .c ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, SB_28_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_28_t0_AND_U1 ( .a ({SubC_in_s2[124], SubC_in_s1[124], SubC_in_s0[124]}), .b ({SubC_in_s2[92], SubC_in_s1[92], SubC_in_s0[92]}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_752, new_AGEMA_signal_751, SB_28_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_28_t1_AND_U1 ( .a ({SubC_in_s2[124], SubC_in_s1[124], SubC_in_s0[124]}), .b ({SubC_in_s2[60], SubC_in_s1[60], SubC_in_s0[60]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_754, new_AGEMA_signal_753, SB_28_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_28_t2_AND_U1 ( .a ({SubC_in_s2[124], SubC_in_s1[124], SubC_in_s0[124]}), .b ({SubC_in_s2[28], SubC_in_s1[28], SubC_in_s0[28]}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_756, new_AGEMA_signal_755, SB_28_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_28_t3_AND_U1 ( .a ({SubC_in_s2[92], SubC_in_s1[92], SubC_in_s0[92]}), .b ({SubC_in_s2[28], SubC_in_s1[28], SubC_in_s0[28]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_758, new_AGEMA_signal_757, SB_28_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U11 ( .a ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, SB_27_n15}), .b ({new_AGEMA_signal_764, new_AGEMA_signal_763, SB_27_n14}), .c ({SubC_out_s2[123], SubC_out_s1[123], SubC_out_s0[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U9 ( .a ({new_AGEMA_signal_764, new_AGEMA_signal_763, SB_27_n14}), .b ({new_AGEMA_signal_776, new_AGEMA_signal_775, SB_27_T2}), .c ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, SB_27_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U6 ( .a ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, SB_27_n11}), .b ({new_AGEMA_signal_774, new_AGEMA_signal_773, SB_27_T1}), .c ({SubC_out_s2[91], SubC_out_s1[91], SubC_out_s0[91]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U5 ( .a ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, SB_27_n15}), .b ({SubC_in_s2[59], SubC_in_s1[59], SubC_in_s0[59]}), .c ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, SB_27_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U4 ( .a ({new_AGEMA_signal_770, new_AGEMA_signal_769, SB_27_n10}), .b ({new_AGEMA_signal_772, new_AGEMA_signal_771, SB_27_T0}), .c ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, SB_27_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U1 ( .a ({SubC_in_s2[123], SubC_in_s1[123], SubC_in_s0[123]}), .b ({new_AGEMA_signal_778, new_AGEMA_signal_777, SB_27_T3}), .c ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, SB_27_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_27_t0_AND_U1 ( .a ({SubC_in_s2[123], SubC_in_s1[123], SubC_in_s0[123]}), .b ({SubC_in_s2[91], SubC_in_s1[91], SubC_in_s0[91]}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_772, new_AGEMA_signal_771, SB_27_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_27_t1_AND_U1 ( .a ({SubC_in_s2[123], SubC_in_s1[123], SubC_in_s0[123]}), .b ({SubC_in_s2[59], SubC_in_s1[59], SubC_in_s0[59]}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_774, new_AGEMA_signal_773, SB_27_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_27_t2_AND_U1 ( .a ({SubC_in_s2[123], SubC_in_s1[123], SubC_in_s0[123]}), .b ({SubC_in_s2[27], SubC_in_s1[27], SubC_in_s0[27]}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_776, new_AGEMA_signal_775, SB_27_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_27_t3_AND_U1 ( .a ({SubC_in_s2[91], SubC_in_s1[91], SubC_in_s0[91]}), .b ({SubC_in_s2[27], SubC_in_s1[27], SubC_in_s0[27]}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_778, new_AGEMA_signal_777, SB_27_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U11 ( .a ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, SB_26_n15}), .b ({new_AGEMA_signal_784, new_AGEMA_signal_783, SB_26_n14}), .c ({SubC_out_s2[122], SubC_out_s1[122], SubC_out_s0[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U9 ( .a ({new_AGEMA_signal_784, new_AGEMA_signal_783, SB_26_n14}), .b ({new_AGEMA_signal_796, new_AGEMA_signal_795, SB_26_T2}), .c ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, SB_26_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U6 ( .a ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, SB_26_n11}), .b ({new_AGEMA_signal_794, new_AGEMA_signal_793, SB_26_T1}), .c ({SubC_out_s2[90], SubC_out_s1[90], SubC_out_s0[90]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U5 ( .a ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, SB_26_n15}), .b ({SubC_in_s2[58], SubC_in_s1[58], SubC_in_s0[58]}), .c ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, SB_26_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U4 ( .a ({new_AGEMA_signal_790, new_AGEMA_signal_789, SB_26_n10}), .b ({new_AGEMA_signal_792, new_AGEMA_signal_791, SB_26_T0}), .c ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, SB_26_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U1 ( .a ({SubC_in_s2[122], SubC_in_s1[122], SubC_in_s0[122]}), .b ({new_AGEMA_signal_798, new_AGEMA_signal_797, SB_26_T3}), .c ({new_AGEMA_signal_1374, new_AGEMA_signal_1373, SB_26_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_26_t0_AND_U1 ( .a ({SubC_in_s2[122], SubC_in_s1[122], SubC_in_s0[122]}), .b ({SubC_in_s2[90], SubC_in_s1[90], SubC_in_s0[90]}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_792, new_AGEMA_signal_791, SB_26_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_26_t1_AND_U1 ( .a ({SubC_in_s2[122], SubC_in_s1[122], SubC_in_s0[122]}), .b ({SubC_in_s2[58], SubC_in_s1[58], SubC_in_s0[58]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_794, new_AGEMA_signal_793, SB_26_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_26_t2_AND_U1 ( .a ({SubC_in_s2[122], SubC_in_s1[122], SubC_in_s0[122]}), .b ({SubC_in_s2[26], SubC_in_s1[26], SubC_in_s0[26]}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_796, new_AGEMA_signal_795, SB_26_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_26_t3_AND_U1 ( .a ({SubC_in_s2[90], SubC_in_s1[90], SubC_in_s0[90]}), .b ({SubC_in_s2[26], SubC_in_s1[26], SubC_in_s0[26]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_798, new_AGEMA_signal_797, SB_26_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U11 ( .a ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, SB_25_n15}), .b ({new_AGEMA_signal_804, new_AGEMA_signal_803, SB_25_n14}), .c ({SubC_out_s2[121], SubC_out_s1[121], SubC_out_s0[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U9 ( .a ({new_AGEMA_signal_804, new_AGEMA_signal_803, SB_25_n14}), .b ({new_AGEMA_signal_816, new_AGEMA_signal_815, SB_25_T2}), .c ({new_AGEMA_signal_1380, new_AGEMA_signal_1379, SB_25_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U6 ( .a ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, SB_25_n11}), .b ({new_AGEMA_signal_814, new_AGEMA_signal_813, SB_25_T1}), .c ({SubC_out_s2[89], SubC_out_s1[89], SubC_out_s0[89]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U5 ( .a ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, SB_25_n15}), .b ({SubC_in_s2[57], SubC_in_s1[57], SubC_in_s0[57]}), .c ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, SB_25_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U4 ( .a ({new_AGEMA_signal_810, new_AGEMA_signal_809, SB_25_n10}), .b ({new_AGEMA_signal_812, new_AGEMA_signal_811, SB_25_T0}), .c ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, SB_25_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U1 ( .a ({SubC_in_s2[121], SubC_in_s1[121], SubC_in_s0[121]}), .b ({new_AGEMA_signal_818, new_AGEMA_signal_817, SB_25_T3}), .c ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, SB_25_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_25_t0_AND_U1 ( .a ({SubC_in_s2[121], SubC_in_s1[121], SubC_in_s0[121]}), .b ({SubC_in_s2[89], SubC_in_s1[89], SubC_in_s0[89]}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_812, new_AGEMA_signal_811, SB_25_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_25_t1_AND_U1 ( .a ({SubC_in_s2[121], SubC_in_s1[121], SubC_in_s0[121]}), .b ({SubC_in_s2[57], SubC_in_s1[57], SubC_in_s0[57]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_814, new_AGEMA_signal_813, SB_25_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_25_t2_AND_U1 ( .a ({SubC_in_s2[121], SubC_in_s1[121], SubC_in_s0[121]}), .b ({SubC_in_s2[25], SubC_in_s1[25], SubC_in_s0[25]}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_816, new_AGEMA_signal_815, SB_25_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_25_t3_AND_U1 ( .a ({SubC_in_s2[89], SubC_in_s1[89], SubC_in_s0[89]}), .b ({SubC_in_s2[25], SubC_in_s1[25], SubC_in_s0[25]}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_818, new_AGEMA_signal_817, SB_25_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U11 ( .a ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, SB_24_n15}), .b ({new_AGEMA_signal_824, new_AGEMA_signal_823, SB_24_n14}), .c ({SubC_out_s2[120], SubC_out_s1[120], SubC_out_s0[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U9 ( .a ({new_AGEMA_signal_824, new_AGEMA_signal_823, SB_24_n14}), .b ({new_AGEMA_signal_836, new_AGEMA_signal_835, SB_24_T2}), .c ({new_AGEMA_signal_1390, new_AGEMA_signal_1389, SB_24_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U6 ( .a ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, SB_24_n11}), .b ({new_AGEMA_signal_834, new_AGEMA_signal_833, SB_24_T1}), .c ({SubC_out_s2[88], SubC_out_s1[88], SubC_out_s0[88]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U5 ( .a ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, SB_24_n15}), .b ({SubC_in_s2[56], SubC_in_s1[56], SubC_in_s0[56]}), .c ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, SB_24_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U4 ( .a ({new_AGEMA_signal_830, new_AGEMA_signal_829, SB_24_n10}), .b ({new_AGEMA_signal_832, new_AGEMA_signal_831, SB_24_T0}), .c ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, SB_24_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U1 ( .a ({SubC_in_s2[120], SubC_in_s1[120], SubC_in_s0[120]}), .b ({new_AGEMA_signal_838, new_AGEMA_signal_837, SB_24_T3}), .c ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, SB_24_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_24_t0_AND_U1 ( .a ({SubC_in_s2[120], SubC_in_s1[120], SubC_in_s0[120]}), .b ({SubC_in_s2[88], SubC_in_s1[88], SubC_in_s0[88]}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_832, new_AGEMA_signal_831, SB_24_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_24_t1_AND_U1 ( .a ({SubC_in_s2[120], SubC_in_s1[120], SubC_in_s0[120]}), .b ({SubC_in_s2[56], SubC_in_s1[56], SubC_in_s0[56]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_834, new_AGEMA_signal_833, SB_24_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_24_t2_AND_U1 ( .a ({SubC_in_s2[120], SubC_in_s1[120], SubC_in_s0[120]}), .b ({SubC_in_s2[24], SubC_in_s1[24], SubC_in_s0[24]}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_836, new_AGEMA_signal_835, SB_24_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_24_t3_AND_U1 ( .a ({SubC_in_s2[88], SubC_in_s1[88], SubC_in_s0[88]}), .b ({SubC_in_s2[24], SubC_in_s1[24], SubC_in_s0[24]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_838, new_AGEMA_signal_837, SB_24_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U11 ( .a ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, SB_23_n15}), .b ({new_AGEMA_signal_844, new_AGEMA_signal_843, SB_23_n14}), .c ({SubC_out_s2[119], SubC_out_s1[119], SubC_out_s0[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U9 ( .a ({new_AGEMA_signal_844, new_AGEMA_signal_843, SB_23_n14}), .b ({new_AGEMA_signal_856, new_AGEMA_signal_855, SB_23_T2}), .c ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, SB_23_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U6 ( .a ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, SB_23_n11}), .b ({new_AGEMA_signal_854, new_AGEMA_signal_853, SB_23_T1}), .c ({SubC_out_s2[87], SubC_out_s1[87], SubC_out_s0[87]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U5 ( .a ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, SB_23_n15}), .b ({SubC_in_s2[55], SubC_in_s1[55], SubC_in_s0[55]}), .c ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, SB_23_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U4 ( .a ({new_AGEMA_signal_850, new_AGEMA_signal_849, SB_23_n10}), .b ({new_AGEMA_signal_852, new_AGEMA_signal_851, SB_23_T0}), .c ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, SB_23_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U1 ( .a ({SubC_in_s2[119], SubC_in_s1[119], SubC_in_s0[119]}), .b ({new_AGEMA_signal_858, new_AGEMA_signal_857, SB_23_T3}), .c ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, SB_23_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_23_t0_AND_U1 ( .a ({SubC_in_s2[119], SubC_in_s1[119], SubC_in_s0[119]}), .b ({SubC_in_s2[87], SubC_in_s1[87], SubC_in_s0[87]}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_852, new_AGEMA_signal_851, SB_23_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_23_t1_AND_U1 ( .a ({SubC_in_s2[119], SubC_in_s1[119], SubC_in_s0[119]}), .b ({SubC_in_s2[55], SubC_in_s1[55], SubC_in_s0[55]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_854, new_AGEMA_signal_853, SB_23_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_23_t2_AND_U1 ( .a ({SubC_in_s2[119], SubC_in_s1[119], SubC_in_s0[119]}), .b ({SubC_in_s2[23], SubC_in_s1[23], SubC_in_s0[23]}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_856, new_AGEMA_signal_855, SB_23_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_23_t3_AND_U1 ( .a ({SubC_in_s2[87], SubC_in_s1[87], SubC_in_s0[87]}), .b ({SubC_in_s2[23], SubC_in_s1[23], SubC_in_s0[23]}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_858, new_AGEMA_signal_857, SB_23_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U11 ( .a ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, SB_22_n15}), .b ({new_AGEMA_signal_864, new_AGEMA_signal_863, SB_22_n14}), .c ({SubC_out_s2[118], SubC_out_s1[118], SubC_out_s0[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U9 ( .a ({new_AGEMA_signal_864, new_AGEMA_signal_863, SB_22_n14}), .b ({new_AGEMA_signal_876, new_AGEMA_signal_875, SB_22_T2}), .c ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, SB_22_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U6 ( .a ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, SB_22_n11}), .b ({new_AGEMA_signal_874, new_AGEMA_signal_873, SB_22_T1}), .c ({SubC_out_s2[86], SubC_out_s1[86], SubC_out_s0[86]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U5 ( .a ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, SB_22_n15}), .b ({SubC_in_s2[54], SubC_in_s1[54], SubC_in_s0[54]}), .c ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, SB_22_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U4 ( .a ({new_AGEMA_signal_870, new_AGEMA_signal_869, SB_22_n10}), .b ({new_AGEMA_signal_872, new_AGEMA_signal_871, SB_22_T0}), .c ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, SB_22_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U1 ( .a ({SubC_in_s2[118], SubC_in_s1[118], SubC_in_s0[118]}), .b ({new_AGEMA_signal_878, new_AGEMA_signal_877, SB_22_T3}), .c ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, SB_22_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_22_t0_AND_U1 ( .a ({SubC_in_s2[118], SubC_in_s1[118], SubC_in_s0[118]}), .b ({SubC_in_s2[86], SubC_in_s1[86], SubC_in_s0[86]}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_872, new_AGEMA_signal_871, SB_22_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_22_t1_AND_U1 ( .a ({SubC_in_s2[118], SubC_in_s1[118], SubC_in_s0[118]}), .b ({SubC_in_s2[54], SubC_in_s1[54], SubC_in_s0[54]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_874, new_AGEMA_signal_873, SB_22_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_22_t2_AND_U1 ( .a ({SubC_in_s2[118], SubC_in_s1[118], SubC_in_s0[118]}), .b ({SubC_in_s2[22], SubC_in_s1[22], SubC_in_s0[22]}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_876, new_AGEMA_signal_875, SB_22_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_22_t3_AND_U1 ( .a ({SubC_in_s2[86], SubC_in_s1[86], SubC_in_s0[86]}), .b ({SubC_in_s2[22], SubC_in_s1[22], SubC_in_s0[22]}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_878, new_AGEMA_signal_877, SB_22_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U11 ( .a ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, SB_21_n15}), .b ({new_AGEMA_signal_884, new_AGEMA_signal_883, SB_21_n14}), .c ({SubC_out_s2[117], SubC_out_s1[117], SubC_out_s0[117]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U9 ( .a ({new_AGEMA_signal_884, new_AGEMA_signal_883, SB_21_n14}), .b ({new_AGEMA_signal_896, new_AGEMA_signal_895, SB_21_T2}), .c ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, SB_21_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U6 ( .a ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, SB_21_n11}), .b ({new_AGEMA_signal_894, new_AGEMA_signal_893, SB_21_T1}), .c ({SubC_out_s2[85], SubC_out_s1[85], SubC_out_s0[85]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U5 ( .a ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, SB_21_n15}), .b ({SubC_in_s2[53], SubC_in_s1[53], SubC_in_s0[53]}), .c ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, SB_21_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U4 ( .a ({new_AGEMA_signal_890, new_AGEMA_signal_889, SB_21_n10}), .b ({new_AGEMA_signal_892, new_AGEMA_signal_891, SB_21_T0}), .c ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, SB_21_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U1 ( .a ({SubC_in_s2[117], SubC_in_s1[117], SubC_in_s0[117]}), .b ({new_AGEMA_signal_898, new_AGEMA_signal_897, SB_21_T3}), .c ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, SB_21_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_21_t0_AND_U1 ( .a ({SubC_in_s2[117], SubC_in_s1[117], SubC_in_s0[117]}), .b ({SubC_in_s2[85], SubC_in_s1[85], SubC_in_s0[85]}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_892, new_AGEMA_signal_891, SB_21_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_21_t1_AND_U1 ( .a ({SubC_in_s2[117], SubC_in_s1[117], SubC_in_s0[117]}), .b ({SubC_in_s2[53], SubC_in_s1[53], SubC_in_s0[53]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_894, new_AGEMA_signal_893, SB_21_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_21_t2_AND_U1 ( .a ({SubC_in_s2[117], SubC_in_s1[117], SubC_in_s0[117]}), .b ({SubC_in_s2[21], SubC_in_s1[21], SubC_in_s0[21]}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_896, new_AGEMA_signal_895, SB_21_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_21_t3_AND_U1 ( .a ({SubC_in_s2[85], SubC_in_s1[85], SubC_in_s0[85]}), .b ({SubC_in_s2[21], SubC_in_s1[21], SubC_in_s0[21]}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_898, new_AGEMA_signal_897, SB_21_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U11 ( .a ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, SB_20_n15}), .b ({new_AGEMA_signal_904, new_AGEMA_signal_903, SB_20_n14}), .c ({SubC_out_s2[116], SubC_out_s1[116], SubC_out_s0[116]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U9 ( .a ({new_AGEMA_signal_904, new_AGEMA_signal_903, SB_20_n14}), .b ({new_AGEMA_signal_916, new_AGEMA_signal_915, SB_20_T2}), .c ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, SB_20_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U6 ( .a ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, SB_20_n11}), .b ({new_AGEMA_signal_914, new_AGEMA_signal_913, SB_20_T1}), .c ({SubC_out_s2[84], SubC_out_s1[84], SubC_out_s0[84]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U5 ( .a ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, SB_20_n15}), .b ({SubC_in_s2[52], SubC_in_s1[52], SubC_in_s0[52]}), .c ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, SB_20_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U4 ( .a ({new_AGEMA_signal_910, new_AGEMA_signal_909, SB_20_n10}), .b ({new_AGEMA_signal_912, new_AGEMA_signal_911, SB_20_T0}), .c ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, SB_20_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U1 ( .a ({SubC_in_s2[116], SubC_in_s1[116], SubC_in_s0[116]}), .b ({new_AGEMA_signal_918, new_AGEMA_signal_917, SB_20_T3}), .c ({new_AGEMA_signal_1434, new_AGEMA_signal_1433, SB_20_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_20_t0_AND_U1 ( .a ({SubC_in_s2[116], SubC_in_s1[116], SubC_in_s0[116]}), .b ({SubC_in_s2[84], SubC_in_s1[84], SubC_in_s0[84]}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_912, new_AGEMA_signal_911, SB_20_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_20_t1_AND_U1 ( .a ({SubC_in_s2[116], SubC_in_s1[116], SubC_in_s0[116]}), .b ({SubC_in_s2[52], SubC_in_s1[52], SubC_in_s0[52]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_914, new_AGEMA_signal_913, SB_20_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_20_t2_AND_U1 ( .a ({SubC_in_s2[116], SubC_in_s1[116], SubC_in_s0[116]}), .b ({SubC_in_s2[20], SubC_in_s1[20], SubC_in_s0[20]}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_916, new_AGEMA_signal_915, SB_20_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_20_t3_AND_U1 ( .a ({SubC_in_s2[84], SubC_in_s1[84], SubC_in_s0[84]}), .b ({SubC_in_s2[20], SubC_in_s1[20], SubC_in_s0[20]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_918, new_AGEMA_signal_917, SB_20_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U11 ( .a ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, SB_19_n15}), .b ({new_AGEMA_signal_924, new_AGEMA_signal_923, SB_19_n14}), .c ({SubC_out_s2[115], SubC_out_s1[115], SubC_out_s0[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U9 ( .a ({new_AGEMA_signal_924, new_AGEMA_signal_923, SB_19_n14}), .b ({new_AGEMA_signal_936, new_AGEMA_signal_935, SB_19_T2}), .c ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, SB_19_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U6 ( .a ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, SB_19_n11}), .b ({new_AGEMA_signal_934, new_AGEMA_signal_933, SB_19_T1}), .c ({SubC_out_s2[83], SubC_out_s1[83], SubC_out_s0[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U5 ( .a ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, SB_19_n15}), .b ({SubC_in_s2[51], SubC_in_s1[51], SubC_in_s0[51]}), .c ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, SB_19_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U4 ( .a ({new_AGEMA_signal_930, new_AGEMA_signal_929, SB_19_n10}), .b ({new_AGEMA_signal_932, new_AGEMA_signal_931, SB_19_T0}), .c ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, SB_19_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U1 ( .a ({SubC_in_s2[115], SubC_in_s1[115], SubC_in_s0[115]}), .b ({new_AGEMA_signal_938, new_AGEMA_signal_937, SB_19_T3}), .c ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, SB_19_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_19_t0_AND_U1 ( .a ({SubC_in_s2[115], SubC_in_s1[115], SubC_in_s0[115]}), .b ({SubC_in_s2[83], SubC_in_s1[83], SubC_in_s0[83]}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_932, new_AGEMA_signal_931, SB_19_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_19_t1_AND_U1 ( .a ({SubC_in_s2[115], SubC_in_s1[115], SubC_in_s0[115]}), .b ({SubC_in_s2[51], SubC_in_s1[51], SubC_in_s0[51]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_934, new_AGEMA_signal_933, SB_19_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_19_t2_AND_U1 ( .a ({SubC_in_s2[115], SubC_in_s1[115], SubC_in_s0[115]}), .b ({SubC_in_s2[19], SubC_in_s1[19], SubC_in_s0[19]}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_936, new_AGEMA_signal_935, SB_19_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_19_t3_AND_U1 ( .a ({SubC_in_s2[83], SubC_in_s1[83], SubC_in_s0[83]}), .b ({SubC_in_s2[19], SubC_in_s1[19], SubC_in_s0[19]}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_938, new_AGEMA_signal_937, SB_19_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U11 ( .a ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, SB_18_n15}), .b ({new_AGEMA_signal_944, new_AGEMA_signal_943, SB_18_n14}), .c ({SubC_out_s2[114], SubC_out_s1[114], SubC_out_s0[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U9 ( .a ({new_AGEMA_signal_944, new_AGEMA_signal_943, SB_18_n14}), .b ({new_AGEMA_signal_956, new_AGEMA_signal_955, SB_18_T2}), .c ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, SB_18_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U6 ( .a ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, SB_18_n11}), .b ({new_AGEMA_signal_954, new_AGEMA_signal_953, SB_18_T1}), .c ({SubC_out_s2[82], SubC_out_s1[82], SubC_out_s0[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U5 ( .a ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, SB_18_n15}), .b ({SubC_in_s2[50], SubC_in_s1[50], SubC_in_s0[50]}), .c ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, SB_18_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U4 ( .a ({new_AGEMA_signal_950, new_AGEMA_signal_949, SB_18_n10}), .b ({new_AGEMA_signal_952, new_AGEMA_signal_951, SB_18_T0}), .c ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, SB_18_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U1 ( .a ({SubC_in_s2[114], SubC_in_s1[114], SubC_in_s0[114]}), .b ({new_AGEMA_signal_958, new_AGEMA_signal_957, SB_18_T3}), .c ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, SB_18_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_18_t0_AND_U1 ( .a ({SubC_in_s2[114], SubC_in_s1[114], SubC_in_s0[114]}), .b ({SubC_in_s2[82], SubC_in_s1[82], SubC_in_s0[82]}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_952, new_AGEMA_signal_951, SB_18_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_18_t1_AND_U1 ( .a ({SubC_in_s2[114], SubC_in_s1[114], SubC_in_s0[114]}), .b ({SubC_in_s2[50], SubC_in_s1[50], SubC_in_s0[50]}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_954, new_AGEMA_signal_953, SB_18_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_18_t2_AND_U1 ( .a ({SubC_in_s2[114], SubC_in_s1[114], SubC_in_s0[114]}), .b ({SubC_in_s2[18], SubC_in_s1[18], SubC_in_s0[18]}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_956, new_AGEMA_signal_955, SB_18_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_18_t3_AND_U1 ( .a ({SubC_in_s2[82], SubC_in_s1[82], SubC_in_s0[82]}), .b ({SubC_in_s2[18], SubC_in_s1[18], SubC_in_s0[18]}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_958, new_AGEMA_signal_957, SB_18_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U11 ( .a ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, SB_17_n15}), .b ({new_AGEMA_signal_964, new_AGEMA_signal_963, SB_17_n14}), .c ({SubC_out_s2[113], SubC_out_s1[113], SubC_out_s0[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U9 ( .a ({new_AGEMA_signal_964, new_AGEMA_signal_963, SB_17_n14}), .b ({new_AGEMA_signal_976, new_AGEMA_signal_975, SB_17_T2}), .c ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, SB_17_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U6 ( .a ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, SB_17_n11}), .b ({new_AGEMA_signal_974, new_AGEMA_signal_973, SB_17_T1}), .c ({SubC_out_s2[81], SubC_out_s1[81], SubC_out_s0[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U5 ( .a ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, SB_17_n15}), .b ({SubC_in_s2[49], SubC_in_s1[49], SubC_in_s0[49]}), .c ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, SB_17_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U4 ( .a ({new_AGEMA_signal_970, new_AGEMA_signal_969, SB_17_n10}), .b ({new_AGEMA_signal_972, new_AGEMA_signal_971, SB_17_T0}), .c ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, SB_17_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U1 ( .a ({SubC_in_s2[113], SubC_in_s1[113], SubC_in_s0[113]}), .b ({new_AGEMA_signal_978, new_AGEMA_signal_977, SB_17_T3}), .c ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, SB_17_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_17_t0_AND_U1 ( .a ({SubC_in_s2[113], SubC_in_s1[113], SubC_in_s0[113]}), .b ({SubC_in_s2[81], SubC_in_s1[81], SubC_in_s0[81]}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_972, new_AGEMA_signal_971, SB_17_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_17_t1_AND_U1 ( .a ({SubC_in_s2[113], SubC_in_s1[113], SubC_in_s0[113]}), .b ({SubC_in_s2[49], SubC_in_s1[49], SubC_in_s0[49]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_974, new_AGEMA_signal_973, SB_17_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_17_t2_AND_U1 ( .a ({SubC_in_s2[113], SubC_in_s1[113], SubC_in_s0[113]}), .b ({SubC_in_s2[17], SubC_in_s1[17], SubC_in_s0[17]}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_976, new_AGEMA_signal_975, SB_17_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_17_t3_AND_U1 ( .a ({SubC_in_s2[81], SubC_in_s1[81], SubC_in_s0[81]}), .b ({SubC_in_s2[17], SubC_in_s1[17], SubC_in_s0[17]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_978, new_AGEMA_signal_977, SB_17_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U11 ( .a ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, SB_16_n15}), .b ({new_AGEMA_signal_984, new_AGEMA_signal_983, SB_16_n14}), .c ({SubC_out_s2[112], SubC_out_s1[112], SubC_out_s0[112]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U9 ( .a ({new_AGEMA_signal_984, new_AGEMA_signal_983, SB_16_n14}), .b ({new_AGEMA_signal_996, new_AGEMA_signal_995, SB_16_T2}), .c ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, SB_16_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U6 ( .a ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, SB_16_n11}), .b ({new_AGEMA_signal_994, new_AGEMA_signal_993, SB_16_T1}), .c ({SubC_out_s2[80], SubC_out_s1[80], SubC_out_s0[80]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U5 ( .a ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, SB_16_n15}), .b ({SubC_in_s2[48], SubC_in_s1[48], SubC_in_s0[48]}), .c ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, SB_16_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U4 ( .a ({new_AGEMA_signal_990, new_AGEMA_signal_989, SB_16_n10}), .b ({new_AGEMA_signal_992, new_AGEMA_signal_991, SB_16_T0}), .c ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, SB_16_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U1 ( .a ({SubC_in_s2[112], SubC_in_s1[112], SubC_in_s0[112]}), .b ({new_AGEMA_signal_998, new_AGEMA_signal_997, SB_16_T3}), .c ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, SB_16_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_16_t0_AND_U1 ( .a ({SubC_in_s2[112], SubC_in_s1[112], SubC_in_s0[112]}), .b ({SubC_in_s2[80], SubC_in_s1[80], SubC_in_s0[80]}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_992, new_AGEMA_signal_991, SB_16_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_16_t1_AND_U1 ( .a ({SubC_in_s2[112], SubC_in_s1[112], SubC_in_s0[112]}), .b ({SubC_in_s2[48], SubC_in_s1[48], SubC_in_s0[48]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_994, new_AGEMA_signal_993, SB_16_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_16_t2_AND_U1 ( .a ({SubC_in_s2[112], SubC_in_s1[112], SubC_in_s0[112]}), .b ({SubC_in_s2[16], SubC_in_s1[16], SubC_in_s0[16]}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_996, new_AGEMA_signal_995, SB_16_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_16_t3_AND_U1 ( .a ({SubC_in_s2[80], SubC_in_s1[80], SubC_in_s0[80]}), .b ({SubC_in_s2[16], SubC_in_s1[16], SubC_in_s0[16]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_998, new_AGEMA_signal_997, SB_16_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U11 ( .a ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, SB_15_n15}), .b ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, SB_15_n14}), .c ({SubC_out_s2[111], SubC_out_s1[111], SubC_out_s0[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U9 ( .a ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, SB_15_n14}), .b ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, SB_15_T2}), .c ({new_AGEMA_signal_1480, new_AGEMA_signal_1479, SB_15_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U6 ( .a ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, SB_15_n11}), .b ({new_AGEMA_signal_1014, new_AGEMA_signal_1013, SB_15_T1}), .c ({SubC_out_s2[79], SubC_out_s1[79], SubC_out_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U5 ( .a ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, SB_15_n15}), .b ({SubC_in_s2[47], SubC_in_s1[47], SubC_in_s0[47]}), .c ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, SB_15_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U4 ( .a ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, SB_15_n10}), .b ({new_AGEMA_signal_1012, new_AGEMA_signal_1011, SB_15_T0}), .c ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, SB_15_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U1 ( .a ({SubC_in_s2[111], SubC_in_s1[111], SubC_in_s0[111]}), .b ({new_AGEMA_signal_1018, new_AGEMA_signal_1017, SB_15_T3}), .c ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, SB_15_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_15_t0_AND_U1 ( .a ({SubC_in_s2[111], SubC_in_s1[111], SubC_in_s0[111]}), .b ({SubC_in_s2[79], SubC_in_s1[79], SubC_in_s0[79]}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1012, new_AGEMA_signal_1011, SB_15_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_15_t1_AND_U1 ( .a ({SubC_in_s2[111], SubC_in_s1[111], SubC_in_s0[111]}), .b ({SubC_in_s2[47], SubC_in_s1[47], SubC_in_s0[47]}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_1014, new_AGEMA_signal_1013, SB_15_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_15_t2_AND_U1 ( .a ({SubC_in_s2[111], SubC_in_s1[111], SubC_in_s0[111]}), .b ({SubC_in_s2[15], SubC_in_s1[15], SubC_in_s0[15]}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, SB_15_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_15_t3_AND_U1 ( .a ({SubC_in_s2[79], SubC_in_s1[79], SubC_in_s0[79]}), .b ({SubC_in_s2[15], SubC_in_s1[15], SubC_in_s0[15]}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_1018, new_AGEMA_signal_1017, SB_15_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U11 ( .a ({new_AGEMA_signal_1492, new_AGEMA_signal_1491, SB_14_n15}), .b ({new_AGEMA_signal_1024, new_AGEMA_signal_1023, SB_14_n14}), .c ({SubC_out_s2[110], SubC_out_s1[110], SubC_out_s0[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U9 ( .a ({new_AGEMA_signal_1024, new_AGEMA_signal_1023, SB_14_n14}), .b ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, SB_14_T2}), .c ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, SB_14_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U6 ( .a ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, SB_14_n11}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SB_14_T1}), .c ({SubC_out_s2[78], SubC_out_s1[78], SubC_out_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U5 ( .a ({new_AGEMA_signal_1492, new_AGEMA_signal_1491, SB_14_n15}), .b ({SubC_in_s2[46], SubC_in_s1[46], SubC_in_s0[46]}), .c ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, SB_14_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U4 ( .a ({new_AGEMA_signal_1030, new_AGEMA_signal_1029, SB_14_n10}), .b ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SB_14_T0}), .c ({new_AGEMA_signal_1492, new_AGEMA_signal_1491, SB_14_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U1 ( .a ({SubC_in_s2[110], SubC_in_s1[110], SubC_in_s0[110]}), .b ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, SB_14_T3}), .c ({new_AGEMA_signal_1494, new_AGEMA_signal_1493, SB_14_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_14_t0_AND_U1 ( .a ({SubC_in_s2[110], SubC_in_s1[110], SubC_in_s0[110]}), .b ({SubC_in_s2[78], SubC_in_s1[78], SubC_in_s0[78]}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, SB_14_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_14_t1_AND_U1 ( .a ({SubC_in_s2[110], SubC_in_s1[110], SubC_in_s0[110]}), .b ({SubC_in_s2[46], SubC_in_s1[46], SubC_in_s0[46]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, SB_14_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_14_t2_AND_U1 ( .a ({SubC_in_s2[110], SubC_in_s1[110], SubC_in_s0[110]}), .b ({SubC_in_s2[14], SubC_in_s1[14], SubC_in_s0[14]}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, SB_14_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_14_t3_AND_U1 ( .a ({SubC_in_s2[78], SubC_in_s1[78], SubC_in_s0[78]}), .b ({SubC_in_s2[14], SubC_in_s1[14], SubC_in_s0[14]}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, SB_14_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U11 ( .a ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, SB_13_n15}), .b ({new_AGEMA_signal_1044, new_AGEMA_signal_1043, SB_13_n14}), .c ({SubC_out_s2[109], SubC_out_s1[109], SubC_out_s0[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U9 ( .a ({new_AGEMA_signal_1044, new_AGEMA_signal_1043, SB_13_n14}), .b ({new_AGEMA_signal_1056, new_AGEMA_signal_1055, SB_13_T2}), .c ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, SB_13_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U6 ( .a ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, SB_13_n11}), .b ({new_AGEMA_signal_1054, new_AGEMA_signal_1053, SB_13_T1}), .c ({SubC_out_s2[77], SubC_out_s1[77], SubC_out_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U5 ( .a ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, SB_13_n15}), .b ({SubC_in_s2[45], SubC_in_s1[45], SubC_in_s0[45]}), .c ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, SB_13_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U4 ( .a ({new_AGEMA_signal_1050, new_AGEMA_signal_1049, SB_13_n10}), .b ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, SB_13_T0}), .c ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, SB_13_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U1 ( .a ({SubC_in_s2[109], SubC_in_s1[109], SubC_in_s0[109]}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, SB_13_T3}), .c ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, SB_13_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_13_t0_AND_U1 ( .a ({SubC_in_s2[109], SubC_in_s1[109], SubC_in_s0[109]}), .b ({SubC_in_s2[77], SubC_in_s1[77], SubC_in_s0[77]}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, SB_13_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_13_t1_AND_U1 ( .a ({SubC_in_s2[109], SubC_in_s1[109], SubC_in_s0[109]}), .b ({SubC_in_s2[45], SubC_in_s1[45], SubC_in_s0[45]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_1054, new_AGEMA_signal_1053, SB_13_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_13_t2_AND_U1 ( .a ({SubC_in_s2[109], SubC_in_s1[109], SubC_in_s0[109]}), .b ({SubC_in_s2[13], SubC_in_s1[13], SubC_in_s0[13]}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1056, new_AGEMA_signal_1055, SB_13_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_13_t3_AND_U1 ( .a ({SubC_in_s2[77], SubC_in_s1[77], SubC_in_s0[77]}), .b ({SubC_in_s2[13], SubC_in_s1[13], SubC_in_s0[13]}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, SB_13_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U11 ( .a ({new_AGEMA_signal_1512, new_AGEMA_signal_1511, SB_12_n15}), .b ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SB_12_n14}), .c ({SubC_out_s2[108], SubC_out_s1[108], SubC_out_s0[108]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U9 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, SB_12_n14}), .b ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, SB_12_T2}), .c ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, SB_12_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U6 ( .a ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, SB_12_n11}), .b ({new_AGEMA_signal_1074, new_AGEMA_signal_1073, SB_12_T1}), .c ({SubC_out_s2[76], SubC_out_s1[76], SubC_out_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U5 ( .a ({new_AGEMA_signal_1512, new_AGEMA_signal_1511, SB_12_n15}), .b ({SubC_in_s2[44], SubC_in_s1[44], SubC_in_s0[44]}), .c ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, SB_12_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U4 ( .a ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, SB_12_n10}), .b ({new_AGEMA_signal_1072, new_AGEMA_signal_1071, SB_12_T0}), .c ({new_AGEMA_signal_1512, new_AGEMA_signal_1511, SB_12_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U1 ( .a ({SubC_in_s2[108], SubC_in_s1[108], SubC_in_s0[108]}), .b ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, SB_12_T3}), .c ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, SB_12_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_12_t0_AND_U1 ( .a ({SubC_in_s2[108], SubC_in_s1[108], SubC_in_s0[108]}), .b ({SubC_in_s2[76], SubC_in_s1[76], SubC_in_s0[76]}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1072, new_AGEMA_signal_1071, SB_12_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_12_t1_AND_U1 ( .a ({SubC_in_s2[108], SubC_in_s1[108], SubC_in_s0[108]}), .b ({SubC_in_s2[44], SubC_in_s1[44], SubC_in_s0[44]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_1074, new_AGEMA_signal_1073, SB_12_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_12_t2_AND_U1 ( .a ({SubC_in_s2[108], SubC_in_s1[108], SubC_in_s0[108]}), .b ({SubC_in_s2[12], SubC_in_s1[12], SubC_in_s0[12]}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, SB_12_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_12_t3_AND_U1 ( .a ({SubC_in_s2[76], SubC_in_s1[76], SubC_in_s0[76]}), .b ({SubC_in_s2[12], SubC_in_s1[12], SubC_in_s0[12]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, SB_12_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U11 ( .a ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, SB_11_n15}), .b ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, SB_11_n14}), .c ({SubC_out_s2[107], SubC_out_s1[107], SubC_out_s0[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U9 ( .a ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, SB_11_n14}), .b ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SB_11_T2}), .c ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, SB_11_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U6 ( .a ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, SB_11_n11}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, SB_11_T1}), .c ({SubC_out_s2[75], SubC_out_s1[75], SubC_out_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U5 ( .a ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, SB_11_n15}), .b ({SubC_in_s2[43], SubC_in_s1[43], SubC_in_s0[43]}), .c ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, SB_11_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U4 ( .a ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, SB_11_n10}), .b ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, SB_11_T0}), .c ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, SB_11_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U1 ( .a ({SubC_in_s2[107], SubC_in_s1[107], SubC_in_s0[107]}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SB_11_T3}), .c ({new_AGEMA_signal_1524, new_AGEMA_signal_1523, SB_11_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_11_t0_AND_U1 ( .a ({SubC_in_s2[107], SubC_in_s1[107], SubC_in_s0[107]}), .b ({SubC_in_s2[75], SubC_in_s1[75], SubC_in_s0[75]}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, SB_11_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_11_t1_AND_U1 ( .a ({SubC_in_s2[107], SubC_in_s1[107], SubC_in_s0[107]}), .b ({SubC_in_s2[43], SubC_in_s1[43], SubC_in_s0[43]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, SB_11_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_11_t2_AND_U1 ( .a ({SubC_in_s2[107], SubC_in_s1[107], SubC_in_s0[107]}), .b ({SubC_in_s2[11], SubC_in_s1[11], SubC_in_s0[11]}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SB_11_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_11_t3_AND_U1 ( .a ({SubC_in_s2[75], SubC_in_s1[75], SubC_in_s0[75]}), .b ({SubC_in_s2[11], SubC_in_s1[11], SubC_in_s0[11]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SB_11_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U11 ( .a ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, SB_10_n15}), .b ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, SB_10_n14}), .c ({SubC_out_s2[106], SubC_out_s1[106], SubC_out_s0[106]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U9 ( .a ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, SB_10_n14}), .b ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, SB_10_T2}), .c ({new_AGEMA_signal_1530, new_AGEMA_signal_1529, SB_10_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U6 ( .a ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, SB_10_n11}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SB_10_T1}), .c ({SubC_out_s2[74], SubC_out_s1[74], SubC_out_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U5 ( .a ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, SB_10_n15}), .b ({SubC_in_s2[42], SubC_in_s1[42], SubC_in_s0[42]}), .c ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, SB_10_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U4 ( .a ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, SB_10_n10}), .b ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SB_10_T0}), .c ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, SB_10_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U1 ( .a ({SubC_in_s2[106], SubC_in_s1[106], SubC_in_s0[106]}), .b ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, SB_10_T3}), .c ({new_AGEMA_signal_1534, new_AGEMA_signal_1533, SB_10_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_10_t0_AND_U1 ( .a ({SubC_in_s2[106], SubC_in_s1[106], SubC_in_s0[106]}), .b ({SubC_in_s2[74], SubC_in_s1[74], SubC_in_s0[74]}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, SB_10_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_10_t1_AND_U1 ( .a ({SubC_in_s2[106], SubC_in_s1[106], SubC_in_s0[106]}), .b ({SubC_in_s2[42], SubC_in_s1[42], SubC_in_s0[42]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, SB_10_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_10_t2_AND_U1 ( .a ({SubC_in_s2[106], SubC_in_s1[106], SubC_in_s0[106]}), .b ({SubC_in_s2[10], SubC_in_s1[10], SubC_in_s0[10]}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, SB_10_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_10_t3_AND_U1 ( .a ({SubC_in_s2[74], SubC_in_s1[74], SubC_in_s0[74]}), .b ({SubC_in_s2[10], SubC_in_s1[10], SubC_in_s0[10]}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, SB_10_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U11 ( .a ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, SB_9_n15}), .b ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, SB_9_n14}), .c ({SubC_out_s2[105], SubC_out_s1[105], SubC_out_s0[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U9 ( .a ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, SB_9_n14}), .b ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, SB_9_T2}), .c ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, SB_9_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U6 ( .a ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, SB_9_n11}), .b ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, SB_9_T1}), .c ({SubC_out_s2[73], SubC_out_s1[73], SubC_out_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U5 ( .a ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, SB_9_n15}), .b ({SubC_in_s2[41], SubC_in_s1[41], SubC_in_s0[41]}), .c ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, SB_9_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U4 ( .a ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, SB_9_n10}), .b ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, SB_9_T0}), .c ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, SB_9_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U1 ( .a ({SubC_in_s2[105], SubC_in_s1[105], SubC_in_s0[105]}), .b ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, SB_9_T3}), .c ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, SB_9_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_9_t0_AND_U1 ( .a ({SubC_in_s2[105], SubC_in_s1[105], SubC_in_s0[105]}), .b ({SubC_in_s2[73], SubC_in_s1[73], SubC_in_s0[73]}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, SB_9_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_9_t1_AND_U1 ( .a ({SubC_in_s2[105], SubC_in_s1[105], SubC_in_s0[105]}), .b ({SubC_in_s2[41], SubC_in_s1[41], SubC_in_s0[41]}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, SB_9_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_9_t2_AND_U1 ( .a ({SubC_in_s2[105], SubC_in_s1[105], SubC_in_s0[105]}), .b ({SubC_in_s2[9], SubC_in_s1[9], SubC_in_s0[9]}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, SB_9_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_9_t3_AND_U1 ( .a ({SubC_in_s2[73], SubC_in_s1[73], SubC_in_s0[73]}), .b ({SubC_in_s2[9], SubC_in_s1[9], SubC_in_s0[9]}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, SB_9_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U11 ( .a ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, SB_8_n15}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SB_8_n14}), .c ({SubC_out_s2[104], SubC_out_s1[104], SubC_out_s0[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U9 ( .a ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, SB_8_n14}), .b ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, SB_8_T2}), .c ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, SB_8_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U6 ( .a ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, SB_8_n11}), .b ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, SB_8_T1}), .c ({SubC_out_s2[72], SubC_out_s1[72], SubC_out_s0[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U5 ( .a ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, SB_8_n15}), .b ({SubC_in_s2[40], SubC_in_s1[40], SubC_in_s0[40]}), .c ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, SB_8_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U4 ( .a ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, SB_8_n10}), .b ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, SB_8_T0}), .c ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, SB_8_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U1 ( .a ({SubC_in_s2[104], SubC_in_s1[104], SubC_in_s0[104]}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, SB_8_T3}), .c ({new_AGEMA_signal_1554, new_AGEMA_signal_1553, SB_8_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_8_t0_AND_U1 ( .a ({SubC_in_s2[104], SubC_in_s1[104], SubC_in_s0[104]}), .b ({SubC_in_s2[72], SubC_in_s1[72], SubC_in_s0[72]}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, SB_8_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_8_t1_AND_U1 ( .a ({SubC_in_s2[104], SubC_in_s1[104], SubC_in_s0[104]}), .b ({SubC_in_s2[40], SubC_in_s1[40], SubC_in_s0[40]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, SB_8_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_8_t2_AND_U1 ( .a ({SubC_in_s2[104], SubC_in_s1[104], SubC_in_s0[104]}), .b ({SubC_in_s2[8], SubC_in_s1[8], SubC_in_s0[8]}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, SB_8_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_8_t3_AND_U1 ( .a ({SubC_in_s2[72], SubC_in_s1[72], SubC_in_s0[72]}), .b ({SubC_in_s2[8], SubC_in_s1[8], SubC_in_s0[8]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, SB_8_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U11 ( .a ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, SB_7_n15}), .b ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, SB_7_n14}), .c ({SubC_out_s2[103], SubC_out_s1[103], SubC_out_s0[103]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U9 ( .a ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, SB_7_n14}), .b ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SB_7_T2}), .c ({new_AGEMA_signal_1560, new_AGEMA_signal_1559, SB_7_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U6 ( .a ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, SB_7_n11}), .b ({new_AGEMA_signal_1174, new_AGEMA_signal_1173, SB_7_T1}), .c ({SubC_out_s2[71], SubC_out_s1[71], SubC_out_s0[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U5 ( .a ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, SB_7_n15}), .b ({SubC_in_s2[39], SubC_in_s1[39], SubC_in_s0[39]}), .c ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, SB_7_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U4 ( .a ({new_AGEMA_signal_1170, new_AGEMA_signal_1169, SB_7_n10}), .b ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, SB_7_T0}), .c ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, SB_7_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U1 ( .a ({SubC_in_s2[103], SubC_in_s1[103], SubC_in_s0[103]}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SB_7_T3}), .c ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, SB_7_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_7_t0_AND_U1 ( .a ({SubC_in_s2[103], SubC_in_s1[103], SubC_in_s0[103]}), .b ({SubC_in_s2[71], SubC_in_s1[71], SubC_in_s0[71]}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, SB_7_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_7_t1_AND_U1 ( .a ({SubC_in_s2[103], SubC_in_s1[103], SubC_in_s0[103]}), .b ({SubC_in_s2[39], SubC_in_s1[39], SubC_in_s0[39]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_1174, new_AGEMA_signal_1173, SB_7_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_7_t2_AND_U1 ( .a ({SubC_in_s2[103], SubC_in_s1[103], SubC_in_s0[103]}), .b ({SubC_in_s2[7], SubC_in_s1[7], SubC_in_s0[7]}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SB_7_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_7_t3_AND_U1 ( .a ({SubC_in_s2[71], SubC_in_s1[71], SubC_in_s0[71]}), .b ({SubC_in_s2[7], SubC_in_s1[7], SubC_in_s0[7]}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SB_7_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U11 ( .a ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, SB_6_n15}), .b ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, SB_6_n14}), .c ({SubC_out_s2[102], SubC_out_s1[102], SubC_out_s0[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U9 ( .a ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, SB_6_n14}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, SB_6_T2}), .c ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, SB_6_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U6 ( .a ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, SB_6_n11}), .b ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SB_6_T1}), .c ({SubC_out_s2[70], SubC_out_s1[70], SubC_out_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U5 ( .a ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, SB_6_n15}), .b ({SubC_in_s2[38], SubC_in_s1[38], SubC_in_s0[38]}), .c ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, SB_6_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U4 ( .a ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, SB_6_n10}), .b ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SB_6_T0}), .c ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, SB_6_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U1 ( .a ({SubC_in_s2[102], SubC_in_s1[102], SubC_in_s0[102]}), .b ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, SB_6_T3}), .c ({new_AGEMA_signal_1574, new_AGEMA_signal_1573, SB_6_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_6_t0_AND_U1 ( .a ({SubC_in_s2[102], SubC_in_s1[102], SubC_in_s0[102]}), .b ({SubC_in_s2[70], SubC_in_s1[70], SubC_in_s0[70]}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, SB_6_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_6_t1_AND_U1 ( .a ({SubC_in_s2[102], SubC_in_s1[102], SubC_in_s0[102]}), .b ({SubC_in_s2[38], SubC_in_s1[38], SubC_in_s0[38]}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_1194, new_AGEMA_signal_1193, SB_6_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_6_t2_AND_U1 ( .a ({SubC_in_s2[102], SubC_in_s1[102], SubC_in_s0[102]}), .b ({SubC_in_s2[6], SubC_in_s1[6], SubC_in_s0[6]}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, SB_6_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_6_t3_AND_U1 ( .a ({SubC_in_s2[70], SubC_in_s1[70], SubC_in_s0[70]}), .b ({SubC_in_s2[6], SubC_in_s1[6], SubC_in_s0[6]}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, SB_6_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U11 ( .a ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, SB_5_n15}), .b ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, SB_5_n14}), .c ({SubC_out_s2[101], SubC_out_s1[101], SubC_out_s0[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U9 ( .a ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, SB_5_n14}), .b ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, SB_5_T2}), .c ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, SB_5_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U6 ( .a ({new_AGEMA_signal_1852, new_AGEMA_signal_1851, SB_5_n11}), .b ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, SB_5_T1}), .c ({SubC_out_s2[69], SubC_out_s1[69], SubC_out_s0[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U5 ( .a ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, SB_5_n15}), .b ({SubC_in_s2[37], SubC_in_s1[37], SubC_in_s0[37]}), .c ({new_AGEMA_signal_1852, new_AGEMA_signal_1851, SB_5_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U4 ( .a ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, SB_5_n10}), .b ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, SB_5_T0}), .c ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, SB_5_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U1 ( .a ({SubC_in_s2[101], SubC_in_s1[101], SubC_in_s0[101]}), .b ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, SB_5_T3}), .c ({new_AGEMA_signal_1584, new_AGEMA_signal_1583, SB_5_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_5_t0_AND_U1 ( .a ({SubC_in_s2[101], SubC_in_s1[101], SubC_in_s0[101]}), .b ({SubC_in_s2[69], SubC_in_s1[69], SubC_in_s0[69]}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, SB_5_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_5_t1_AND_U1 ( .a ({SubC_in_s2[101], SubC_in_s1[101], SubC_in_s0[101]}), .b ({SubC_in_s2[37], SubC_in_s1[37], SubC_in_s0[37]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, SB_5_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_5_t2_AND_U1 ( .a ({SubC_in_s2[101], SubC_in_s1[101], SubC_in_s0[101]}), .b ({SubC_in_s2[5], SubC_in_s1[5], SubC_in_s0[5]}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, SB_5_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_5_t3_AND_U1 ( .a ({SubC_in_s2[69], SubC_in_s1[69], SubC_in_s0[69]}), .b ({SubC_in_s2[5], SubC_in_s1[5], SubC_in_s0[5]}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, SB_5_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U11 ( .a ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, SB_4_n15}), .b ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SB_4_n14}), .c ({SubC_out_s2[100], SubC_out_s1[100], SubC_out_s0[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U9 ( .a ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, SB_4_n14}), .b ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, SB_4_T2}), .c ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, SB_4_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U6 ( .a ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, SB_4_n11}), .b ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, SB_4_T1}), .c ({SubC_out_s2[68], SubC_out_s1[68], SubC_out_s0[68]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U5 ( .a ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, SB_4_n15}), .b ({SubC_in_s2[36], SubC_in_s1[36], SubC_in_s0[36]}), .c ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, SB_4_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U4 ( .a ({new_AGEMA_signal_1230, new_AGEMA_signal_1229, SB_4_n10}), .b ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, SB_4_T0}), .c ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, SB_4_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U1 ( .a ({SubC_in_s2[100], SubC_in_s1[100], SubC_in_s0[100]}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, SB_4_T3}), .c ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, SB_4_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_4_t0_AND_U1 ( .a ({SubC_in_s2[100], SubC_in_s1[100], SubC_in_s0[100]}), .b ({SubC_in_s2[68], SubC_in_s1[68], SubC_in_s0[68]}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, SB_4_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_4_t1_AND_U1 ( .a ({SubC_in_s2[100], SubC_in_s1[100], SubC_in_s0[100]}), .b ({SubC_in_s2[36], SubC_in_s1[36], SubC_in_s0[36]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, SB_4_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_4_t2_AND_U1 ( .a ({SubC_in_s2[100], SubC_in_s1[100], SubC_in_s0[100]}), .b ({SubC_in_s2[4], SubC_in_s1[4], SubC_in_s0[4]}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, SB_4_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_4_t3_AND_U1 ( .a ({SubC_in_s2[68], SubC_in_s1[68], SubC_in_s0[68]}), .b ({SubC_in_s2[4], SubC_in_s1[4], SubC_in_s0[4]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, SB_4_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U11 ( .a ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, SB_3_n15}), .b ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, SB_3_n14}), .c ({SubC_out_s2[99], SubC_out_s1[99], SubC_out_s0[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U9 ( .a ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, SB_3_n14}), .b ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SB_3_T2}), .c ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, SB_3_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U6 ( .a ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, SB_3_n11}), .b ({new_AGEMA_signal_1254, new_AGEMA_signal_1253, SB_3_T1}), .c ({SubC_out_s2[67], SubC_out_s1[67], SubC_out_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U5 ( .a ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, SB_3_n15}), .b ({SubC_in_s2[35], SubC_in_s1[35], SubC_in_s0[35]}), .c ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, SB_3_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U4 ( .a ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, SB_3_n10}), .b ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, SB_3_T0}), .c ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, SB_3_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U1 ( .a ({SubC_in_s2[99], SubC_in_s1[99], SubC_in_s0[99]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SB_3_T3}), .c ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, SB_3_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_3_t0_AND_U1 ( .a ({SubC_in_s2[99], SubC_in_s1[99], SubC_in_s0[99]}), .b ({SubC_in_s2[67], SubC_in_s1[67], SubC_in_s0[67]}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, SB_3_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_3_t1_AND_U1 ( .a ({SubC_in_s2[99], SubC_in_s1[99], SubC_in_s0[99]}), .b ({SubC_in_s2[35], SubC_in_s1[35], SubC_in_s0[35]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_1254, new_AGEMA_signal_1253, SB_3_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_3_t2_AND_U1 ( .a ({SubC_in_s2[99], SubC_in_s1[99], SubC_in_s0[99]}), .b ({SubC_in_s2[3], SubC_in_s1[3], SubC_in_s0[3]}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SB_3_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_3_t3_AND_U1 ( .a ({SubC_in_s2[67], SubC_in_s1[67], SubC_in_s0[67]}), .b ({SubC_in_s2[3], SubC_in_s1[3], SubC_in_s0[3]}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SB_3_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U11 ( .a ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, SB_2_n15}), .b ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, SB_2_n14}), .c ({SubC_out_s2[98], SubC_out_s1[98], SubC_out_s0[98]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U9 ( .a ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, SB_2_n14}), .b ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SB_2_T2}), .c ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, SB_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U6 ( .a ({new_AGEMA_signal_1876, new_AGEMA_signal_1875, SB_2_n11}), .b ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SB_2_T1}), .c ({SubC_out_s2[66], SubC_out_s1[66], SubC_out_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U5 ( .a ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, SB_2_n15}), .b ({SubC_in_s2[34], SubC_in_s1[34], SubC_in_s0[34]}), .c ({new_AGEMA_signal_1876, new_AGEMA_signal_1875, SB_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U4 ( .a ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, SB_2_n10}), .b ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SB_2_T0}), .c ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, SB_2_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U1 ( .a ({SubC_in_s2[98], SubC_in_s1[98], SubC_in_s0[98]}), .b ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SB_2_T3}), .c ({new_AGEMA_signal_1614, new_AGEMA_signal_1613, SB_2_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_2_t0_AND_U1 ( .a ({SubC_in_s2[98], SubC_in_s1[98], SubC_in_s0[98]}), .b ({SubC_in_s2[66], SubC_in_s1[66], SubC_in_s0[66]}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, SB_2_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_2_t1_AND_U1 ( .a ({SubC_in_s2[98], SubC_in_s1[98], SubC_in_s0[98]}), .b ({SubC_in_s2[34], SubC_in_s1[34], SubC_in_s0[34]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, SB_2_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_2_t2_AND_U1 ( .a ({SubC_in_s2[98], SubC_in_s1[98], SubC_in_s0[98]}), .b ({SubC_in_s2[2], SubC_in_s1[2], SubC_in_s0[2]}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SB_2_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_2_t3_AND_U1 ( .a ({SubC_in_s2[66], SubC_in_s1[66], SubC_in_s0[66]}), .b ({SubC_in_s2[2], SubC_in_s1[2], SubC_in_s0[2]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SB_2_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U11 ( .a ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, SB_1_n15}), .b ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, SB_1_n14}), .c ({SubC_out_s2[97], SubC_out_s1[97], SubC_out_s0[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U9 ( .a ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, SB_1_n14}), .b ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, SB_1_T2}), .c ({new_AGEMA_signal_1620, new_AGEMA_signal_1619, SB_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U6 ( .a ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, SB_1_n11}), .b ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, SB_1_T1}), .c ({SubC_out_s2[65], SubC_out_s1[65], SubC_out_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U5 ( .a ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, SB_1_n15}), .b ({SubC_in_s2[33], SubC_in_s1[33], SubC_in_s0[33]}), .c ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, SB_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U4 ( .a ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, SB_1_n10}), .b ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, SB_1_T0}), .c ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, SB_1_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U1 ( .a ({SubC_in_s2[97], SubC_in_s1[97], SubC_in_s0[97]}), .b ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SB_1_T3}), .c ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, SB_1_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_1_t0_AND_U1 ( .a ({SubC_in_s2[97], SubC_in_s1[97], SubC_in_s0[97]}), .b ({SubC_in_s2[65], SubC_in_s1[65], SubC_in_s0[65]}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, SB_1_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_1_t1_AND_U1 ( .a ({SubC_in_s2[97], SubC_in_s1[97], SubC_in_s0[97]}), .b ({SubC_in_s2[33], SubC_in_s1[33], SubC_in_s0[33]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, SB_1_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_1_t2_AND_U1 ( .a ({SubC_in_s2[97], SubC_in_s1[97], SubC_in_s0[97]}), .b ({SubC_in_s2[1], SubC_in_s1[1], SubC_in_s0[1]}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, SB_1_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_1_t3_AND_U1 ( .a ({SubC_in_s2[65], SubC_in_s1[65], SubC_in_s0[65]}), .b ({SubC_in_s2[1], SubC_in_s1[1], SubC_in_s0[1]}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SB_1_T3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U11 ( .a ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, SB_0_n15}), .b ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, SB_0_n14}), .c ({SubC_out_s2[96], SubC_out_s1[96], SubC_out_s0[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U9 ( .a ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, SB_0_n14}), .b ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, SB_0_T2}), .c ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, SB_0_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U6 ( .a ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, SB_0_n11}), .b ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, SB_0_T1}), .c ({SubC_out_s2[64], SubC_out_s1[64], SubC_out_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U5 ( .a ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, SB_0_n15}), .b ({SubC_in_s2[32], SubC_in_s1[32], SubC_in_s0[32]}), .c ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, SB_0_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U4 ( .a ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, SB_0_n10}), .b ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, SB_0_T0}), .c ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, SB_0_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U1 ( .a ({SubC_in_s2[96], SubC_in_s1[96], SubC_in_s0[96]}), .b ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, SB_0_T3}), .c ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, SB_0_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_0_t0_AND_U1 ( .a ({SubC_in_s2[96], SubC_in_s1[96], SubC_in_s0[96]}), .b ({SubC_in_s2[64], SubC_in_s1[64], SubC_in_s0[64]}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, SB_0_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_0_t1_AND_U1 ( .a ({SubC_in_s2[96], SubC_in_s1[96], SubC_in_s0[96]}), .b ({SubC_in_s2[32], SubC_in_s1[32], SubC_in_s0[32]}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_1314, new_AGEMA_signal_1313, SB_0_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_0_t2_AND_U1 ( .a ({SubC_in_s2[96], SubC_in_s1[96], SubC_in_s0[96]}), .b ({SubC_in_s2[0], SubC_in_s1[0], SubC_in_s0[0]}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, SB_0_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_0_t3_AND_U1 ( .a ({SubC_in_s2[64], SubC_in_s1[64], SubC_in_s0[64]}), .b ({SubC_in_s2[0], SubC_in_s1[0], SubC_in_s0[0]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, SB_0_T3}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U10 ( .a ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, SB_31_n13}), .b ({new_AGEMA_signal_1320, new_AGEMA_signal_1319, SB_31_n12}), .c ({SubC_out_s2[63], SubC_out_s1[63], SubC_out_s0[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U7 ( .a ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, SB_31_T4}), .b ({new_AGEMA_signal_698, new_AGEMA_signal_697, SB_31_T3}), .c ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, SB_31_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_31_U2 ( .a ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, SB_31_n9}), .b ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, SB_31_T5}), .c ({SubC_out_s2[31], SubC_out_s1[31], SubC_out_s0[31]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_31_t4_AND_U1 ( .a ({SubC_in_s2[63], SubC_in_s1[63], SubC_in_s0[63]}), .b ({new_AGEMA_signal_698, new_AGEMA_signal_697, SB_31_T3}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, SB_31_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_31_t5_AND_U1 ( .a ({SubC_in_s2[63], SubC_in_s1[63], SubC_in_s0[63]}), .b ({new_AGEMA_signal_696, new_AGEMA_signal_695, SB_31_T2}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, SB_31_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U10 ( .a ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, SB_30_n13}), .b ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, SB_30_n12}), .c ({SubC_out_s2[62], SubC_out_s1[62], SubC_out_s0[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U7 ( .a ({new_AGEMA_signal_1336, new_AGEMA_signal_1335, SB_30_T4}), .b ({new_AGEMA_signal_718, new_AGEMA_signal_717, SB_30_T3}), .c ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, SB_30_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_30_U2 ( .a ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, SB_30_n9}), .b ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, SB_30_T5}), .c ({SubC_out_s2[30], SubC_out_s1[30], SubC_out_s0[30]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_30_t4_AND_U1 ( .a ({SubC_in_s2[62], SubC_in_s1[62], SubC_in_s0[62]}), .b ({new_AGEMA_signal_718, new_AGEMA_signal_717, SB_30_T3}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1336, new_AGEMA_signal_1335, SB_30_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_30_t5_AND_U1 ( .a ({SubC_in_s2[62], SubC_in_s1[62], SubC_in_s0[62]}), .b ({new_AGEMA_signal_716, new_AGEMA_signal_715, SB_30_T2}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, SB_30_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U10 ( .a ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, SB_29_n13}), .b ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, SB_29_n12}), .c ({SubC_out_s2[61], SubC_out_s1[61], SubC_out_s0[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U7 ( .a ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, SB_29_T4}), .b ({new_AGEMA_signal_738, new_AGEMA_signal_737, SB_29_T3}), .c ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, SB_29_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_29_U2 ( .a ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, SB_29_n9}), .b ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, SB_29_T5}), .c ({SubC_out_s2[29], SubC_out_s1[29], SubC_out_s0[29]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_29_t4_AND_U1 ( .a ({SubC_in_s2[61], SubC_in_s1[61], SubC_in_s0[61]}), .b ({new_AGEMA_signal_738, new_AGEMA_signal_737, SB_29_T3}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, SB_29_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_29_t5_AND_U1 ( .a ({SubC_in_s2[61], SubC_in_s1[61], SubC_in_s0[61]}), .b ({new_AGEMA_signal_736, new_AGEMA_signal_735, SB_29_T2}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, SB_29_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U10 ( .a ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, SB_28_n13}), .b ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, SB_28_n12}), .c ({SubC_out_s2[60], SubC_out_s1[60], SubC_out_s0[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U7 ( .a ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, SB_28_T4}), .b ({new_AGEMA_signal_758, new_AGEMA_signal_757, SB_28_T3}), .c ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, SB_28_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_28_U2 ( .a ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, SB_28_n9}), .b ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, SB_28_T5}), .c ({SubC_out_s2[28], SubC_out_s1[28], SubC_out_s0[28]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_28_t4_AND_U1 ( .a ({SubC_in_s2[60], SubC_in_s1[60], SubC_in_s0[60]}), .b ({new_AGEMA_signal_758, new_AGEMA_signal_757, SB_28_T3}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, SB_28_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_28_t5_AND_U1 ( .a ({SubC_in_s2[60], SubC_in_s1[60], SubC_in_s0[60]}), .b ({new_AGEMA_signal_756, new_AGEMA_signal_755, SB_28_T2}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, SB_28_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U10 ( .a ({new_AGEMA_signal_1674, new_AGEMA_signal_1673, SB_27_n13}), .b ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, SB_27_n12}), .c ({SubC_out_s2[59], SubC_out_s1[59], SubC_out_s0[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U7 ( .a ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, SB_27_T4}), .b ({new_AGEMA_signal_778, new_AGEMA_signal_777, SB_27_T3}), .c ({new_AGEMA_signal_1674, new_AGEMA_signal_1673, SB_27_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_27_U2 ( .a ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, SB_27_n9}), .b ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, SB_27_T5}), .c ({SubC_out_s2[27], SubC_out_s1[27], SubC_out_s0[27]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_27_t4_AND_U1 ( .a ({SubC_in_s2[59], SubC_in_s1[59], SubC_in_s0[59]}), .b ({new_AGEMA_signal_778, new_AGEMA_signal_777, SB_27_T3}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, SB_27_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_27_t5_AND_U1 ( .a ({SubC_in_s2[59], SubC_in_s1[59], SubC_in_s0[59]}), .b ({new_AGEMA_signal_776, new_AGEMA_signal_775, SB_27_T2}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, SB_27_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U10 ( .a ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, SB_26_n13}), .b ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, SB_26_n12}), .c ({SubC_out_s2[58], SubC_out_s1[58], SubC_out_s0[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U7 ( .a ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, SB_26_T4}), .b ({new_AGEMA_signal_798, new_AGEMA_signal_797, SB_26_T3}), .c ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, SB_26_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_26_U2 ( .a ({new_AGEMA_signal_1374, new_AGEMA_signal_1373, SB_26_n9}), .b ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, SB_26_T5}), .c ({SubC_out_s2[26], SubC_out_s1[26], SubC_out_s0[26]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_26_t4_AND_U1 ( .a ({SubC_in_s2[58], SubC_in_s1[58], SubC_in_s0[58]}), .b ({new_AGEMA_signal_798, new_AGEMA_signal_797, SB_26_T3}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, SB_26_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_26_t5_AND_U1 ( .a ({SubC_in_s2[58], SubC_in_s1[58], SubC_in_s0[58]}), .b ({new_AGEMA_signal_796, new_AGEMA_signal_795, SB_26_T2}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, SB_26_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U10 ( .a ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, SB_25_n13}), .b ({new_AGEMA_signal_1380, new_AGEMA_signal_1379, SB_25_n12}), .c ({SubC_out_s2[57], SubC_out_s1[57], SubC_out_s0[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U7 ( .a ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, SB_25_T4}), .b ({new_AGEMA_signal_818, new_AGEMA_signal_817, SB_25_T3}), .c ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, SB_25_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_25_U2 ( .a ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, SB_25_n9}), .b ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, SB_25_T5}), .c ({SubC_out_s2[25], SubC_out_s1[25], SubC_out_s0[25]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_25_t4_AND_U1 ( .a ({SubC_in_s2[57], SubC_in_s1[57], SubC_in_s0[57]}), .b ({new_AGEMA_signal_818, new_AGEMA_signal_817, SB_25_T3}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, SB_25_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_25_t5_AND_U1 ( .a ({SubC_in_s2[57], SubC_in_s1[57], SubC_in_s0[57]}), .b ({new_AGEMA_signal_816, new_AGEMA_signal_815, SB_25_T2}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, SB_25_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U10 ( .a ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, SB_24_n13}), .b ({new_AGEMA_signal_1390, new_AGEMA_signal_1389, SB_24_n12}), .c ({SubC_out_s2[56], SubC_out_s1[56], SubC_out_s0[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U7 ( .a ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, SB_24_T4}), .b ({new_AGEMA_signal_838, new_AGEMA_signal_837, SB_24_T3}), .c ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, SB_24_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_24_U2 ( .a ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, SB_24_n9}), .b ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, SB_24_T5}), .c ({SubC_out_s2[24], SubC_out_s1[24], SubC_out_s0[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_24_t4_AND_U1 ( .a ({SubC_in_s2[56], SubC_in_s1[56], SubC_in_s0[56]}), .b ({new_AGEMA_signal_838, new_AGEMA_signal_837, SB_24_T3}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, SB_24_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_24_t5_AND_U1 ( .a ({SubC_in_s2[56], SubC_in_s1[56], SubC_in_s0[56]}), .b ({new_AGEMA_signal_836, new_AGEMA_signal_835, SB_24_T2}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, SB_24_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U10 ( .a ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, SB_23_n13}), .b ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, SB_23_n12}), .c ({SubC_out_s2[55], SubC_out_s1[55], SubC_out_s0[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U7 ( .a ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, SB_23_T4}), .b ({new_AGEMA_signal_858, new_AGEMA_signal_857, SB_23_T3}), .c ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, SB_23_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_23_U2 ( .a ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, SB_23_n9}), .b ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, SB_23_T5}), .c ({SubC_out_s2[23], SubC_out_s1[23], SubC_out_s0[23]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_23_t4_AND_U1 ( .a ({SubC_in_s2[55], SubC_in_s1[55], SubC_in_s0[55]}), .b ({new_AGEMA_signal_858, new_AGEMA_signal_857, SB_23_T3}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, SB_23_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_23_t5_AND_U1 ( .a ({SubC_in_s2[55], SubC_in_s1[55], SubC_in_s0[55]}), .b ({new_AGEMA_signal_856, new_AGEMA_signal_855, SB_23_T2}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, SB_23_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U10 ( .a ({new_AGEMA_signal_1714, new_AGEMA_signal_1713, SB_22_n13}), .b ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, SB_22_n12}), .c ({SubC_out_s2[54], SubC_out_s1[54], SubC_out_s0[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U7 ( .a ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, SB_22_T4}), .b ({new_AGEMA_signal_878, new_AGEMA_signal_877, SB_22_T3}), .c ({new_AGEMA_signal_1714, new_AGEMA_signal_1713, SB_22_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_22_U2 ( .a ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, SB_22_n9}), .b ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, SB_22_T5}), .c ({SubC_out_s2[22], SubC_out_s1[22], SubC_out_s0[22]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_22_t4_AND_U1 ( .a ({SubC_in_s2[54], SubC_in_s1[54], SubC_in_s0[54]}), .b ({new_AGEMA_signal_878, new_AGEMA_signal_877, SB_22_T3}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, SB_22_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_22_t5_AND_U1 ( .a ({SubC_in_s2[54], SubC_in_s1[54], SubC_in_s0[54]}), .b ({new_AGEMA_signal_876, new_AGEMA_signal_875, SB_22_T2}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, SB_22_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U10 ( .a ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, SB_21_n13}), .b ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, SB_21_n12}), .c ({SubC_out_s2[53], SubC_out_s1[53], SubC_out_s0[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U7 ( .a ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, SB_21_T4}), .b ({new_AGEMA_signal_898, new_AGEMA_signal_897, SB_21_T3}), .c ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, SB_21_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_21_U2 ( .a ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, SB_21_n9}), .b ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, SB_21_T5}), .c ({SubC_out_s2[21], SubC_out_s1[21], SubC_out_s0[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_21_t4_AND_U1 ( .a ({SubC_in_s2[53], SubC_in_s1[53], SubC_in_s0[53]}), .b ({new_AGEMA_signal_898, new_AGEMA_signal_897, SB_21_T3}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, SB_21_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_21_t5_AND_U1 ( .a ({SubC_in_s2[53], SubC_in_s1[53], SubC_in_s0[53]}), .b ({new_AGEMA_signal_896, new_AGEMA_signal_895, SB_21_T2}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, SB_21_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U10 ( .a ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, SB_20_n13}), .b ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, SB_20_n12}), .c ({SubC_out_s2[52], SubC_out_s1[52], SubC_out_s0[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U7 ( .a ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, SB_20_T4}), .b ({new_AGEMA_signal_918, new_AGEMA_signal_917, SB_20_T3}), .c ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, SB_20_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_20_U2 ( .a ({new_AGEMA_signal_1434, new_AGEMA_signal_1433, SB_20_n9}), .b ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, SB_20_T5}), .c ({SubC_out_s2[20], SubC_out_s1[20], SubC_out_s0[20]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_20_t4_AND_U1 ( .a ({SubC_in_s2[52], SubC_in_s1[52], SubC_in_s0[52]}), .b ({new_AGEMA_signal_918, new_AGEMA_signal_917, SB_20_T3}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, SB_20_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_20_t5_AND_U1 ( .a ({SubC_in_s2[52], SubC_in_s1[52], SubC_in_s0[52]}), .b ({new_AGEMA_signal_916, new_AGEMA_signal_915, SB_20_T2}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, SB_20_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U10 ( .a ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, SB_19_n13}), .b ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, SB_19_n12}), .c ({SubC_out_s2[51], SubC_out_s1[51], SubC_out_s0[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U7 ( .a ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, SB_19_T4}), .b ({new_AGEMA_signal_938, new_AGEMA_signal_937, SB_19_T3}), .c ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, SB_19_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_19_U2 ( .a ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, SB_19_n9}), .b ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, SB_19_T5}), .c ({SubC_out_s2[19], SubC_out_s1[19], SubC_out_s0[19]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_19_t4_AND_U1 ( .a ({SubC_in_s2[51], SubC_in_s1[51], SubC_in_s0[51]}), .b ({new_AGEMA_signal_938, new_AGEMA_signal_937, SB_19_T3}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, SB_19_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_19_t5_AND_U1 ( .a ({SubC_in_s2[51], SubC_in_s1[51], SubC_in_s0[51]}), .b ({new_AGEMA_signal_936, new_AGEMA_signal_935, SB_19_T2}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, SB_19_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U10 ( .a ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, SB_18_n13}), .b ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, SB_18_n12}), .c ({SubC_out_s2[50], SubC_out_s1[50], SubC_out_s0[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U7 ( .a ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, SB_18_T4}), .b ({new_AGEMA_signal_958, new_AGEMA_signal_957, SB_18_T3}), .c ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, SB_18_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_18_U2 ( .a ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, SB_18_n9}), .b ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, SB_18_T5}), .c ({SubC_out_s2[18], SubC_out_s1[18], SubC_out_s0[18]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_18_t4_AND_U1 ( .a ({SubC_in_s2[50], SubC_in_s1[50], SubC_in_s0[50]}), .b ({new_AGEMA_signal_958, new_AGEMA_signal_957, SB_18_T3}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, SB_18_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_18_t5_AND_U1 ( .a ({SubC_in_s2[50], SubC_in_s1[50], SubC_in_s0[50]}), .b ({new_AGEMA_signal_956, new_AGEMA_signal_955, SB_18_T2}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, SB_18_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U10 ( .a ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, SB_17_n13}), .b ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, SB_17_n12}), .c ({SubC_out_s2[49], SubC_out_s1[49], SubC_out_s0[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U7 ( .a ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, SB_17_T4}), .b ({new_AGEMA_signal_978, new_AGEMA_signal_977, SB_17_T3}), .c ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, SB_17_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_17_U2 ( .a ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, SB_17_n9}), .b ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, SB_17_T5}), .c ({SubC_out_s2[17], SubC_out_s1[17], SubC_out_s0[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_17_t4_AND_U1 ( .a ({SubC_in_s2[49], SubC_in_s1[49], SubC_in_s0[49]}), .b ({new_AGEMA_signal_978, new_AGEMA_signal_977, SB_17_T3}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, SB_17_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_17_t5_AND_U1 ( .a ({SubC_in_s2[49], SubC_in_s1[49], SubC_in_s0[49]}), .b ({new_AGEMA_signal_976, new_AGEMA_signal_975, SB_17_T2}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, SB_17_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U10 ( .a ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, SB_16_n13}), .b ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, SB_16_n12}), .c ({SubC_out_s2[48], SubC_out_s1[48], SubC_out_s0[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U7 ( .a ({new_AGEMA_signal_1476, new_AGEMA_signal_1475, SB_16_T4}), .b ({new_AGEMA_signal_998, new_AGEMA_signal_997, SB_16_T3}), .c ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, SB_16_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_16_U2 ( .a ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, SB_16_n9}), .b ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, SB_16_T5}), .c ({SubC_out_s2[16], SubC_out_s1[16], SubC_out_s0[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_16_t4_AND_U1 ( .a ({SubC_in_s2[48], SubC_in_s1[48], SubC_in_s0[48]}), .b ({new_AGEMA_signal_998, new_AGEMA_signal_997, SB_16_T3}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1476, new_AGEMA_signal_1475, SB_16_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_16_t5_AND_U1 ( .a ({SubC_in_s2[48], SubC_in_s1[48], SubC_in_s0[48]}), .b ({new_AGEMA_signal_996, new_AGEMA_signal_995, SB_16_T2}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, SB_16_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U10 ( .a ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, SB_15_n13}), .b ({new_AGEMA_signal_1480, new_AGEMA_signal_1479, SB_15_n12}), .c ({SubC_out_s2[47], SubC_out_s1[47], SubC_out_s0[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U7 ( .a ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, SB_15_T4}), .b ({new_AGEMA_signal_1018, new_AGEMA_signal_1017, SB_15_T3}), .c ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, SB_15_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_15_U2 ( .a ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, SB_15_n9}), .b ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, SB_15_T5}), .c ({SubC_out_s2[15], SubC_out_s1[15], SubC_out_s0[15]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_15_t4_AND_U1 ( .a ({SubC_in_s2[47], SubC_in_s1[47], SubC_in_s0[47]}), .b ({new_AGEMA_signal_1018, new_AGEMA_signal_1017, SB_15_T3}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, SB_15_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_15_t5_AND_U1 ( .a ({SubC_in_s2[47], SubC_in_s1[47], SubC_in_s0[47]}), .b ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, SB_15_T2}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, SB_15_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U10 ( .a ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, SB_14_n13}), .b ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, SB_14_n12}), .c ({SubC_out_s2[46], SubC_out_s1[46], SubC_out_s0[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U7 ( .a ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, SB_14_T4}), .b ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, SB_14_T3}), .c ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, SB_14_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_14_U2 ( .a ({new_AGEMA_signal_1494, new_AGEMA_signal_1493, SB_14_n9}), .b ({new_AGEMA_signal_1498, new_AGEMA_signal_1497, SB_14_T5}), .c ({SubC_out_s2[14], SubC_out_s1[14], SubC_out_s0[14]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_14_t4_AND_U1 ( .a ({SubC_in_s2[46], SubC_in_s1[46], SubC_in_s0[46]}), .b ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, SB_14_T3}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, SB_14_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_14_t5_AND_U1 ( .a ({SubC_in_s2[46], SubC_in_s1[46], SubC_in_s0[46]}), .b ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, SB_14_T2}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_1498, new_AGEMA_signal_1497, SB_14_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U10 ( .a ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, SB_13_n13}), .b ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, SB_13_n12}), .c ({SubC_out_s2[45], SubC_out_s1[45], SubC_out_s0[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U7 ( .a ({new_AGEMA_signal_1506, new_AGEMA_signal_1505, SB_13_T4}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, SB_13_T3}), .c ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, SB_13_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_13_U2 ( .a ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, SB_13_n9}), .b ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, SB_13_T5}), .c ({SubC_out_s2[13], SubC_out_s1[13], SubC_out_s0[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_13_t4_AND_U1 ( .a ({SubC_in_s2[45], SubC_in_s1[45], SubC_in_s0[45]}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, SB_13_T3}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1506, new_AGEMA_signal_1505, SB_13_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_13_t5_AND_U1 ( .a ({SubC_in_s2[45], SubC_in_s1[45], SubC_in_s0[45]}), .b ({new_AGEMA_signal_1056, new_AGEMA_signal_1055, SB_13_T2}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, SB_13_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U10 ( .a ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, SB_12_n13}), .b ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, SB_12_n12}), .c ({SubC_out_s2[44], SubC_out_s1[44], SubC_out_s0[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U7 ( .a ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, SB_12_T4}), .b ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, SB_12_T3}), .c ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, SB_12_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_12_U2 ( .a ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, SB_12_n9}), .b ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, SB_12_T5}), .c ({SubC_out_s2[12], SubC_out_s1[12], SubC_out_s0[12]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_12_t4_AND_U1 ( .a ({SubC_in_s2[44], SubC_in_s1[44], SubC_in_s0[44]}), .b ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, SB_12_T3}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, SB_12_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_12_t5_AND_U1 ( .a ({SubC_in_s2[44], SubC_in_s1[44], SubC_in_s0[44]}), .b ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, SB_12_T2}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, SB_12_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U10 ( .a ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, SB_11_n13}), .b ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, SB_11_n12}), .c ({SubC_out_s2[43], SubC_out_s1[43], SubC_out_s0[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U7 ( .a ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, SB_11_T4}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SB_11_T3}), .c ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, SB_11_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_11_U2 ( .a ({new_AGEMA_signal_1524, new_AGEMA_signal_1523, SB_11_n9}), .b ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, SB_11_T5}), .c ({SubC_out_s2[11], SubC_out_s1[11], SubC_out_s0[11]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_11_t4_AND_U1 ( .a ({SubC_in_s2[43], SubC_in_s1[43], SubC_in_s0[43]}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, SB_11_T3}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, SB_11_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_11_t5_AND_U1 ( .a ({SubC_in_s2[43], SubC_in_s1[43], SubC_in_s0[43]}), .b ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, SB_11_T2}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, SB_11_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U10 ( .a ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, SB_10_n13}), .b ({new_AGEMA_signal_1530, new_AGEMA_signal_1529, SB_10_n12}), .c ({SubC_out_s2[42], SubC_out_s1[42], SubC_out_s0[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U7 ( .a ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, SB_10_T4}), .b ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, SB_10_T3}), .c ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, SB_10_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_10_U2 ( .a ({new_AGEMA_signal_1534, new_AGEMA_signal_1533, SB_10_n9}), .b ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, SB_10_T5}), .c ({SubC_out_s2[10], SubC_out_s1[10], SubC_out_s0[10]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_10_t4_AND_U1 ( .a ({SubC_in_s2[42], SubC_in_s1[42], SubC_in_s0[42]}), .b ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, SB_10_T3}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, SB_10_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_10_t5_AND_U1 ( .a ({SubC_in_s2[42], SubC_in_s1[42], SubC_in_s0[42]}), .b ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, SB_10_T2}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, SB_10_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U10 ( .a ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, SB_9_n13}), .b ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, SB_9_n12}), .c ({SubC_out_s2[41], SubC_out_s1[41], SubC_out_s0[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U7 ( .a ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, SB_9_T4}), .b ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, SB_9_T3}), .c ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, SB_9_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_9_U2 ( .a ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, SB_9_n9}), .b ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, SB_9_T5}), .c ({SubC_out_s2[9], SubC_out_s1[9], SubC_out_s0[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_9_t4_AND_U1 ( .a ({SubC_in_s2[41], SubC_in_s1[41], SubC_in_s0[41]}), .b ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, SB_9_T3}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, SB_9_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_9_t5_AND_U1 ( .a ({SubC_in_s2[41], SubC_in_s1[41], SubC_in_s0[41]}), .b ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, SB_9_T2}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, SB_9_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U10 ( .a ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, SB_8_n13}), .b ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, SB_8_n12}), .c ({SubC_out_s2[40], SubC_out_s1[40], SubC_out_s0[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U7 ( .a ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, SB_8_T4}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, SB_8_T3}), .c ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, SB_8_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_8_U2 ( .a ({new_AGEMA_signal_1554, new_AGEMA_signal_1553, SB_8_n9}), .b ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, SB_8_T5}), .c ({SubC_out_s2[8], SubC_out_s1[8], SubC_out_s0[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_8_t4_AND_U1 ( .a ({SubC_in_s2[40], SubC_in_s1[40], SubC_in_s0[40]}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, SB_8_T3}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, SB_8_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_8_t5_AND_U1 ( .a ({SubC_in_s2[40], SubC_in_s1[40], SubC_in_s0[40]}), .b ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, SB_8_T2}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, SB_8_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U10 ( .a ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, SB_7_n13}), .b ({new_AGEMA_signal_1560, new_AGEMA_signal_1559, SB_7_n12}), .c ({SubC_out_s2[39], SubC_out_s1[39], SubC_out_s0[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U7 ( .a ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, SB_7_T4}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SB_7_T3}), .c ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, SB_7_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_7_U2 ( .a ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, SB_7_n9}), .b ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, SB_7_T5}), .c ({SubC_out_s2[7], SubC_out_s1[7], SubC_out_s0[7]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_7_t4_AND_U1 ( .a ({SubC_in_s2[39], SubC_in_s1[39], SubC_in_s0[39]}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, SB_7_T3}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, SB_7_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_7_t5_AND_U1 ( .a ({SubC_in_s2[39], SubC_in_s1[39], SubC_in_s0[39]}), .b ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, SB_7_T2}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, SB_7_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U10 ( .a ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, SB_6_n13}), .b ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, SB_6_n12}), .c ({SubC_out_s2[38], SubC_out_s1[38], SubC_out_s0[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U7 ( .a ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, SB_6_T4}), .b ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, SB_6_T3}), .c ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, SB_6_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_6_U2 ( .a ({new_AGEMA_signal_1574, new_AGEMA_signal_1573, SB_6_n9}), .b ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, SB_6_T5}), .c ({SubC_out_s2[6], SubC_out_s1[6], SubC_out_s0[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_6_t4_AND_U1 ( .a ({SubC_in_s2[38], SubC_in_s1[38], SubC_in_s0[38]}), .b ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, SB_6_T3}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, SB_6_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_6_t5_AND_U1 ( .a ({SubC_in_s2[38], SubC_in_s1[38], SubC_in_s0[38]}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, SB_6_T2}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, SB_6_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U10 ( .a ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, SB_5_n13}), .b ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, SB_5_n12}), .c ({SubC_out_s2[37], SubC_out_s1[37], SubC_out_s0[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U7 ( .a ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, SB_5_T4}), .b ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, SB_5_T3}), .c ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, SB_5_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_5_U2 ( .a ({new_AGEMA_signal_1584, new_AGEMA_signal_1583, SB_5_n9}), .b ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, SB_5_T5}), .c ({SubC_out_s2[5], SubC_out_s1[5], SubC_out_s0[5]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_5_t4_AND_U1 ( .a ({SubC_in_s2[37], SubC_in_s1[37], SubC_in_s0[37]}), .b ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, SB_5_T3}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, SB_5_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_5_t5_AND_U1 ( .a ({SubC_in_s2[37], SubC_in_s1[37], SubC_in_s0[37]}), .b ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, SB_5_T2}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, SB_5_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U10 ( .a ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, SB_4_n13}), .b ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, SB_4_n12}), .c ({SubC_out_s2[36], SubC_out_s1[36], SubC_out_s0[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U7 ( .a ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, SB_4_T4}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, SB_4_T3}), .c ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, SB_4_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_4_U2 ( .a ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, SB_4_n9}), .b ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, SB_4_T5}), .c ({SubC_out_s2[4], SubC_out_s1[4], SubC_out_s0[4]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_4_t4_AND_U1 ( .a ({SubC_in_s2[36], SubC_in_s1[36], SubC_in_s0[36]}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, SB_4_T3}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, SB_4_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_4_t5_AND_U1 ( .a ({SubC_in_s2[36], SubC_in_s1[36], SubC_in_s0[36]}), .b ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, SB_4_T2}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, SB_4_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U10 ( .a ({new_AGEMA_signal_1866, new_AGEMA_signal_1865, SB_3_n13}), .b ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, SB_3_n12}), .c ({SubC_out_s2[35], SubC_out_s1[35], SubC_out_s0[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U7 ( .a ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, SB_3_T4}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SB_3_T3}), .c ({new_AGEMA_signal_1866, new_AGEMA_signal_1865, SB_3_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_3_U2 ( .a ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, SB_3_n9}), .b ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, SB_3_T5}), .c ({SubC_out_s2[3], SubC_out_s1[3], SubC_out_s0[3]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_3_t4_AND_U1 ( .a ({SubC_in_s2[35], SubC_in_s1[35], SubC_in_s0[35]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, SB_3_T3}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, SB_3_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_3_t5_AND_U1 ( .a ({SubC_in_s2[35], SubC_in_s1[35], SubC_in_s0[35]}), .b ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, SB_3_T2}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, SB_3_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U10 ( .a ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, SB_2_n13}), .b ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, SB_2_n12}), .c ({SubC_out_s2[34], SubC_out_s1[34], SubC_out_s0[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U7 ( .a ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, SB_2_T4}), .b ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SB_2_T3}), .c ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, SB_2_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_2_U2 ( .a ({new_AGEMA_signal_1614, new_AGEMA_signal_1613, SB_2_n9}), .b ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, SB_2_T5}), .c ({SubC_out_s2[2], SubC_out_s1[2], SubC_out_s0[2]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_2_t4_AND_U1 ( .a ({SubC_in_s2[34], SubC_in_s1[34], SubC_in_s0[34]}), .b ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, SB_2_T3}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, SB_2_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_2_t5_AND_U1 ( .a ({SubC_in_s2[34], SubC_in_s1[34], SubC_in_s0[34]}), .b ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, SB_2_T2}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, SB_2_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U10 ( .a ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, SB_1_n13}), .b ({new_AGEMA_signal_1620, new_AGEMA_signal_1619, SB_1_n12}), .c ({SubC_out_s2[33], SubC_out_s1[33], SubC_out_s0[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U7 ( .a ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, SB_1_T4}), .b ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SB_1_T3}), .c ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, SB_1_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_1_U2 ( .a ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, SB_1_n9}), .b ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, SB_1_T5}), .c ({SubC_out_s2[1], SubC_out_s1[1], SubC_out_s0[1]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_1_t4_AND_U1 ( .a ({SubC_in_s2[33], SubC_in_s1[33], SubC_in_s0[33]}), .b ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, SB_1_T3}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, SB_1_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_1_t5_AND_U1 ( .a ({SubC_in_s2[33], SubC_in_s1[33], SubC_in_s0[33]}), .b ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, SB_1_T2}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, SB_1_T5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U10 ( .a ({new_AGEMA_signal_1890, new_AGEMA_signal_1889, SB_0_n13}), .b ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, SB_0_n12}), .c ({SubC_out_s2[32], SubC_out_s1[32], SubC_out_s0[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U7 ( .a ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, SB_0_T4}), .b ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, SB_0_T3}), .c ({new_AGEMA_signal_1890, new_AGEMA_signal_1889, SB_0_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SB_0_U2 ( .a ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, SB_0_n9}), .b ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, SB_0_T5}), .c ({SubC_out_s2[0], SubC_out_s1[0], SubC_out_s0[0]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_0_t4_AND_U1 ( .a ({SubC_in_s2[32], SubC_in_s1[32], SubC_in_s0[32]}), .b ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, SB_0_T3}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, SB_0_T4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SB_0_t5_AND_U1 ( .a ({SubC_in_s2[32], SubC_in_s1[32], SubC_in_s0[32]}), .b ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, SB_0_T2}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, SB_0_T5}) ) ;

endmodule
