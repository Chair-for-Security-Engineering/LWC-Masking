/* clock gating is added to the circuit, the latency increased 10 time(s)  */

module arx_round_HPC2_ClockGating_d1 (round_constant, round, x_round_in_s0, y_round_in_s0, clk, y_round_in_s1, x_round_in_s1, Fresh, /*rst,*/ x_round_out_s0, y_round_out_s0, x_round_out_s1, y_round_out_s1/*, Synch*/);
    input [31:0] round_constant ;
    input [1:0] round ;
    input [31:0] x_round_in_s0 ;
    input [31:0] y_round_in_s0 ;
    input clk ;
    input [31:0] y_round_in_s1 ;
    input [31:0] x_round_in_s1 ;
    //input rst ;
    input [255:0] Fresh ;
    output [31:0] x_round_out_s0 ;
    output [31:0] y_round_out_s0 ;
    output [31:0] x_round_out_s1 ;
    output [31:0] y_round_out_s1 ;
    //output Synch ;
    wire AdderIns_s2_gc_0_a1_t ;
    wire AdderIns_s2_bc_0_a1_t ;
    wire AdderIns_s2_bc_1_a1_t ;
    wire AdderIns_s2_bc_2_a1_t ;
    wire AdderIns_s2_bc_3_a1_t ;
    wire AdderIns_s2_bc_4_a1_t ;
    wire AdderIns_s2_bc_5_a1_t ;
    wire AdderIns_s2_bc_6_a1_t ;
    wire AdderIns_s2_bc_7_a1_t ;
    wire AdderIns_s2_bc_8_a1_t ;
    wire AdderIns_s2_bc_9_a1_t ;
    wire AdderIns_s2_bc_10_a1_t ;
    wire AdderIns_s2_bc_11_a1_t ;
    wire AdderIns_s2_bc_12_a1_t ;
    wire AdderIns_s2_bc_13_a1_t ;
    wire AdderIns_s2_bc_14_a1_t ;
    wire AdderIns_s2_bc_15_a1_t ;
    wire AdderIns_s2_bc_16_a1_t ;
    wire AdderIns_s2_bc_17_a1_t ;
    wire AdderIns_s2_bc_18_a1_t ;
    wire AdderIns_s2_bc_19_a1_t ;
    wire AdderIns_s2_bc_20_a1_t ;
    wire AdderIns_s2_bc_21_a1_t ;
    wire AdderIns_s2_bc_22_a1_t ;
    wire AdderIns_s2_bc_23_a1_t ;
    wire AdderIns_s2_bc_24_a1_t ;
    wire AdderIns_s2_bc_25_a1_t ;
    wire AdderIns_s2_bc_26_a1_t ;
    wire AdderIns_s2_bc_27_a1_t ;
    wire AdderIns_s2_bc_28_a1_t ;
    wire AdderIns_s2_bc_29_a1_t ;
    wire AdderIns_s3_gc_0_a1_t ;
    wire AdderIns_s3_gc_1_a1_t ;
    wire AdderIns_s3_bc_0_a1_t ;
    wire AdderIns_s3_bc_1_a1_t ;
    wire AdderIns_s3_bc_2_a1_t ;
    wire AdderIns_s3_bc_3_a1_t ;
    wire AdderIns_s3_bc_4_a1_t ;
    wire AdderIns_s3_bc_5_a1_t ;
    wire AdderIns_s3_bc_6_a1_t ;
    wire AdderIns_s3_bc_7_a1_t ;
    wire AdderIns_s3_bc_8_a1_t ;
    wire AdderIns_s3_bc_9_a1_t ;
    wire AdderIns_s3_bc_10_a1_t ;
    wire AdderIns_s3_bc_11_a1_t ;
    wire AdderIns_s3_bc_12_a1_t ;
    wire AdderIns_s3_bc_13_a1_t ;
    wire AdderIns_s3_bc_14_a1_t ;
    wire AdderIns_s3_bc_15_a1_t ;
    wire AdderIns_s3_bc_16_a1_t ;
    wire AdderIns_s3_bc_17_a1_t ;
    wire AdderIns_s3_bc_18_a1_t ;
    wire AdderIns_s3_bc_19_a1_t ;
    wire AdderIns_s3_bc_20_a1_t ;
    wire AdderIns_s3_bc_21_a1_t ;
    wire AdderIns_s3_bc_22_a1_t ;
    wire AdderIns_s3_bc_23_a1_t ;
    wire AdderIns_s3_bc_24_a1_t ;
    wire AdderIns_s3_bc_25_a1_t ;
    wire AdderIns_s3_bc_26_a1_t ;
    wire AdderIns_s3_bc_27_a1_t ;
    wire AdderIns_s4_gc_0_a1_t ;
    wire AdderIns_s4_gc_1_a1_t ;
    wire AdderIns_s4_gc_2_a1_t ;
    wire AdderIns_s4_gc_3_a1_t ;
    wire AdderIns_s4_bc_0_a1_t ;
    wire AdderIns_s4_bc_1_a1_t ;
    wire AdderIns_s4_bc_2_a1_t ;
    wire AdderIns_s4_bc_3_a1_t ;
    wire AdderIns_s4_bc_4_a1_t ;
    wire AdderIns_s4_bc_5_a1_t ;
    wire AdderIns_s4_bc_6_a1_t ;
    wire AdderIns_s4_bc_7_a1_t ;
    wire AdderIns_s4_bc_8_a1_t ;
    wire AdderIns_s4_bc_9_a1_t ;
    wire AdderIns_s4_bc_10_a1_t ;
    wire AdderIns_s4_bc_11_a1_t ;
    wire AdderIns_s4_bc_12_a1_t ;
    wire AdderIns_s4_bc_13_a1_t ;
    wire AdderIns_s4_bc_14_a1_t ;
    wire AdderIns_s4_bc_15_a1_t ;
    wire AdderIns_s4_bc_16_a1_t ;
    wire AdderIns_s4_bc_17_a1_t ;
    wire AdderIns_s4_bc_18_a1_t ;
    wire AdderIns_s4_bc_19_a1_t ;
    wire AdderIns_s4_bc_20_a1_t ;
    wire AdderIns_s4_bc_21_a1_t ;
    wire AdderIns_s4_bc_22_a1_t ;
    wire AdderIns_s4_bc_23_a1_t ;
    wire AdderIns_s5_gc_0_a1_t ;
    wire AdderIns_s5_gc_1_a1_t ;
    wire AdderIns_s5_gc_2_a1_t ;
    wire AdderIns_s5_gc_3_a1_t ;
    wire AdderIns_s5_gc_4_a1_t ;
    wire AdderIns_s5_gc_5_a1_t ;
    wire AdderIns_s5_gc_6_a1_t ;
    wire AdderIns_s5_gc_7_a1_t ;
    wire AdderIns_s5_bc_0_a1_t ;
    wire AdderIns_s5_bc_1_a1_t ;
    wire AdderIns_s5_bc_2_a1_t ;
    wire AdderIns_s5_bc_3_a1_t ;
    wire AdderIns_s5_bc_4_a1_t ;
    wire AdderIns_s5_bc_5_a1_t ;
    wire AdderIns_s5_bc_6_a1_t ;
    wire AdderIns_s5_bc_7_a1_t ;
    wire AdderIns_s5_bc_8_a1_t ;
    wire AdderIns_s5_bc_9_a1_t ;
    wire AdderIns_s5_bc_10_a1_t ;
    wire AdderIns_s5_bc_11_a1_t ;
    wire AdderIns_s5_bc_12_a1_t ;
    wire AdderIns_s5_bc_13_a1_t ;
    wire AdderIns_s5_bc_14_a1_t ;
    wire AdderIns_s5_bc_15_a1_t ;
    wire AdderIns_s6_gc_1_a1_t ;
    wire AdderIns_s6_gc_2_a1_t ;
    wire AdderIns_s6_gc_3_a1_t ;
    wire AdderIns_s6_gc_4_a1_t ;
    wire AdderIns_s6_gc_5_a1_t ;
    wire AdderIns_s6_gc_6_a1_t ;
    wire AdderIns_s6_gc_7_a1_t ;
    wire AdderIns_s6_gc_8_a1_t ;
    wire AdderIns_s6_gc_9_a1_t ;
    wire AdderIns_s6_gc_10_a1_t ;
    wire AdderIns_s6_gc_11_a1_t ;
    wire AdderIns_s6_gc_12_a1_t ;
    wire AdderIns_s6_gc_13_a1_t ;
    wire AdderIns_s6_gc_14_a1_t ;
    wire AdderIns_s6_gc_15_a1_t ;
    wire [31:0] y_rotated01 ;
    wire [31:0] y_rotated23 ;
    wire [31:0] y_rotated ;
    wire [31:0] sum ;
    wire [31:0] sum_rotated01 ;
    wire [31:0] sum_rotated23 ;
    wire [31:0] sum_rotated ;
    wire [30:0] AdderIns_g6 ;
    wire [31:1] AdderIns_p6 ;
    wire [30:16] AdderIns_g5 ;
    wire [15:1] AdderIns_p5 ;
    wire [30:7] AdderIns_g4 ;
    wire [23:0] AdderIns_p4 ;
    wire [30:3] AdderIns_g3 ;
    wire [27:0] AdderIns_p3 ;
    wire [30:1] AdderIns_g2 ;
    wire [29:0] AdderIns_p2 ;
    wire [30:0] AdderIns_g1 ;
    wire new_AGEMA_signal_826 ;
    wire new_AGEMA_signal_829 ;
    wire new_AGEMA_signal_832 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_838 ;
    wire new_AGEMA_signal_841 ;
    wire new_AGEMA_signal_844 ;
    wire new_AGEMA_signal_847 ;
    wire new_AGEMA_signal_850 ;
    wire new_AGEMA_signal_853 ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_859 ;
    wire new_AGEMA_signal_862 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_869 ;
    wire new_AGEMA_signal_871 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_874 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_878 ;
    wire new_AGEMA_signal_879 ;
    wire new_AGEMA_signal_880 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_886 ;
    wire new_AGEMA_signal_887 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_890 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_892 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_896 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_898 ;
    wire new_AGEMA_signal_899 ;
    wire new_AGEMA_signal_900 ;
    wire new_AGEMA_signal_901 ;
    wire new_AGEMA_signal_902 ;
    wire new_AGEMA_signal_903 ;
    wire new_AGEMA_signal_904 ;
    wire new_AGEMA_signal_905 ;
    wire new_AGEMA_signal_906 ;
    wire new_AGEMA_signal_907 ;
    wire new_AGEMA_signal_908 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_910 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_912 ;
    wire new_AGEMA_signal_913 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_915 ;
    wire new_AGEMA_signal_916 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_919 ;
    wire new_AGEMA_signal_920 ;
    wire new_AGEMA_signal_921 ;
    wire new_AGEMA_signal_922 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_924 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_928 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_930 ;
    wire new_AGEMA_signal_931 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_934 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_939 ;
    wire new_AGEMA_signal_940 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_942 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) U129 ( .a ({1'b0, round_constant[0]}), .b ({new_AGEMA_signal_953, sum[0]}), .c ({x_round_out_s1[0], x_round_out_s0[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_0_U1 ( .s (round[0]), .b ({y_round_in_s1[31], y_round_in_s0[31]}), .a ({y_round_in_s1[17], y_round_in_s0[17]}), .c ({new_AGEMA_signal_826, y_rotated01[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_1_U1 ( .s (round[0]), .b ({y_round_in_s1[0], y_round_in_s0[0]}), .a ({y_round_in_s1[18], y_round_in_s0[18]}), .c ({new_AGEMA_signal_829, y_rotated01[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_2_U1 ( .s (round[0]), .b ({y_round_in_s1[1], y_round_in_s0[1]}), .a ({y_round_in_s1[19], y_round_in_s0[19]}), .c ({new_AGEMA_signal_832, y_rotated01[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_3_U1 ( .s (round[0]), .b ({y_round_in_s1[2], y_round_in_s0[2]}), .a ({y_round_in_s1[20], y_round_in_s0[20]}), .c ({new_AGEMA_signal_835, y_rotated01[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_4_U1 ( .s (round[0]), .b ({y_round_in_s1[3], y_round_in_s0[3]}), .a ({y_round_in_s1[21], y_round_in_s0[21]}), .c ({new_AGEMA_signal_838, y_rotated01[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_5_U1 ( .s (round[0]), .b ({y_round_in_s1[4], y_round_in_s0[4]}), .a ({y_round_in_s1[22], y_round_in_s0[22]}), .c ({new_AGEMA_signal_841, y_rotated01[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_6_U1 ( .s (round[0]), .b ({y_round_in_s1[5], y_round_in_s0[5]}), .a ({y_round_in_s1[23], y_round_in_s0[23]}), .c ({new_AGEMA_signal_844, y_rotated01[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_7_U1 ( .s (round[0]), .b ({y_round_in_s1[6], y_round_in_s0[6]}), .a ({y_round_in_s1[24], y_round_in_s0[24]}), .c ({new_AGEMA_signal_847, y_rotated01[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_8_U1 ( .s (round[0]), .b ({y_round_in_s1[7], y_round_in_s0[7]}), .a ({y_round_in_s1[25], y_round_in_s0[25]}), .c ({new_AGEMA_signal_850, y_rotated01[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_9_U1 ( .s (round[0]), .b ({y_round_in_s1[8], y_round_in_s0[8]}), .a ({y_round_in_s1[26], y_round_in_s0[26]}), .c ({new_AGEMA_signal_853, y_rotated01[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_10_U1 ( .s (round[0]), .b ({y_round_in_s1[9], y_round_in_s0[9]}), .a ({y_round_in_s1[27], y_round_in_s0[27]}), .c ({new_AGEMA_signal_856, y_rotated01[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_11_U1 ( .s (round[0]), .b ({y_round_in_s1[10], y_round_in_s0[10]}), .a ({y_round_in_s1[28], y_round_in_s0[28]}), .c ({new_AGEMA_signal_859, y_rotated01[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_12_U1 ( .s (round[0]), .b ({y_round_in_s1[11], y_round_in_s0[11]}), .a ({y_round_in_s1[29], y_round_in_s0[29]}), .c ({new_AGEMA_signal_862, y_rotated01[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_13_U1 ( .s (round[0]), .b ({y_round_in_s1[12], y_round_in_s0[12]}), .a ({y_round_in_s1[30], y_round_in_s0[30]}), .c ({new_AGEMA_signal_865, y_rotated01[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_14_U1 ( .s (round[0]), .b ({y_round_in_s1[13], y_round_in_s0[13]}), .a ({y_round_in_s1[31], y_round_in_s0[31]}), .c ({new_AGEMA_signal_867, y_rotated01[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_15_U1 ( .s (round[0]), .b ({y_round_in_s1[14], y_round_in_s0[14]}), .a ({y_round_in_s1[0], y_round_in_s0[0]}), .c ({new_AGEMA_signal_869, y_rotated01[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_16_U1 ( .s (round[0]), .b ({y_round_in_s1[15], y_round_in_s0[15]}), .a ({y_round_in_s1[1], y_round_in_s0[1]}), .c ({new_AGEMA_signal_871, y_rotated01[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_17_U1 ( .s (round[0]), .b ({y_round_in_s1[16], y_round_in_s0[16]}), .a ({y_round_in_s1[2], y_round_in_s0[2]}), .c ({new_AGEMA_signal_873, y_rotated01[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_18_U1 ( .s (round[0]), .b ({y_round_in_s1[17], y_round_in_s0[17]}), .a ({y_round_in_s1[3], y_round_in_s0[3]}), .c ({new_AGEMA_signal_874, y_rotated01[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_19_U1 ( .s (round[0]), .b ({y_round_in_s1[18], y_round_in_s0[18]}), .a ({y_round_in_s1[4], y_round_in_s0[4]}), .c ({new_AGEMA_signal_875, y_rotated01[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_20_U1 ( .s (round[0]), .b ({y_round_in_s1[19], y_round_in_s0[19]}), .a ({y_round_in_s1[5], y_round_in_s0[5]}), .c ({new_AGEMA_signal_876, y_rotated01[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_21_U1 ( .s (round[0]), .b ({y_round_in_s1[20], y_round_in_s0[20]}), .a ({y_round_in_s1[6], y_round_in_s0[6]}), .c ({new_AGEMA_signal_877, y_rotated01[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_22_U1 ( .s (round[0]), .b ({y_round_in_s1[21], y_round_in_s0[21]}), .a ({y_round_in_s1[7], y_round_in_s0[7]}), .c ({new_AGEMA_signal_878, y_rotated01[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_23_U1 ( .s (round[0]), .b ({y_round_in_s1[22], y_round_in_s0[22]}), .a ({y_round_in_s1[8], y_round_in_s0[8]}), .c ({new_AGEMA_signal_879, y_rotated01[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_24_U1 ( .s (round[0]), .b ({y_round_in_s1[23], y_round_in_s0[23]}), .a ({y_round_in_s1[9], y_round_in_s0[9]}), .c ({new_AGEMA_signal_880, y_rotated01[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_25_U1 ( .s (round[0]), .b ({y_round_in_s1[24], y_round_in_s0[24]}), .a ({y_round_in_s1[10], y_round_in_s0[10]}), .c ({new_AGEMA_signal_881, y_rotated01[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_26_U1 ( .s (round[0]), .b ({y_round_in_s1[25], y_round_in_s0[25]}), .a ({y_round_in_s1[11], y_round_in_s0[11]}), .c ({new_AGEMA_signal_882, y_rotated01[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_27_U1 ( .s (round[0]), .b ({y_round_in_s1[26], y_round_in_s0[26]}), .a ({y_round_in_s1[12], y_round_in_s0[12]}), .c ({new_AGEMA_signal_883, y_rotated01[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_28_U1 ( .s (round[0]), .b ({y_round_in_s1[27], y_round_in_s0[27]}), .a ({y_round_in_s1[13], y_round_in_s0[13]}), .c ({new_AGEMA_signal_884, y_rotated01[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_29_U1 ( .s (round[0]), .b ({y_round_in_s1[28], y_round_in_s0[28]}), .a ({y_round_in_s1[14], y_round_in_s0[14]}), .c ({new_AGEMA_signal_885, y_rotated01[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_30_U1 ( .s (round[0]), .b ({y_round_in_s1[29], y_round_in_s0[29]}), .a ({y_round_in_s1[15], y_round_in_s0[15]}), .c ({new_AGEMA_signal_886, y_rotated01[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M0_mux_inst_31_U1 ( .s (round[0]), .b ({y_round_in_s1[30], y_round_in_s0[30]}), .a ({y_round_in_s1[16], y_round_in_s0[16]}), .c ({new_AGEMA_signal_887, y_rotated01[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_0_U1 ( .s (round[0]), .b ({y_round_in_s1[0], y_round_in_s0[0]}), .a ({y_round_in_s1[24], y_round_in_s0[24]}), .c ({new_AGEMA_signal_888, y_rotated23[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_1_U1 ( .s (round[0]), .b ({y_round_in_s1[1], y_round_in_s0[1]}), .a ({y_round_in_s1[25], y_round_in_s0[25]}), .c ({new_AGEMA_signal_889, y_rotated23[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_2_U1 ( .s (round[0]), .b ({y_round_in_s1[2], y_round_in_s0[2]}), .a ({y_round_in_s1[26], y_round_in_s0[26]}), .c ({new_AGEMA_signal_890, y_rotated23[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_3_U1 ( .s (round[0]), .b ({y_round_in_s1[3], y_round_in_s0[3]}), .a ({y_round_in_s1[27], y_round_in_s0[27]}), .c ({new_AGEMA_signal_891, y_rotated23[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_4_U1 ( .s (round[0]), .b ({y_round_in_s1[4], y_round_in_s0[4]}), .a ({y_round_in_s1[28], y_round_in_s0[28]}), .c ({new_AGEMA_signal_892, y_rotated23[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_5_U1 ( .s (round[0]), .b ({y_round_in_s1[5], y_round_in_s0[5]}), .a ({y_round_in_s1[29], y_round_in_s0[29]}), .c ({new_AGEMA_signal_893, y_rotated23[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_6_U1 ( .s (round[0]), .b ({y_round_in_s1[6], y_round_in_s0[6]}), .a ({y_round_in_s1[30], y_round_in_s0[30]}), .c ({new_AGEMA_signal_894, y_rotated23[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_7_U1 ( .s (round[0]), .b ({y_round_in_s1[7], y_round_in_s0[7]}), .a ({y_round_in_s1[31], y_round_in_s0[31]}), .c ({new_AGEMA_signal_895, y_rotated23[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_8_U1 ( .s (round[0]), .b ({y_round_in_s1[8], y_round_in_s0[8]}), .a ({y_round_in_s1[0], y_round_in_s0[0]}), .c ({new_AGEMA_signal_896, y_rotated23[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_9_U1 ( .s (round[0]), .b ({y_round_in_s1[9], y_round_in_s0[9]}), .a ({y_round_in_s1[1], y_round_in_s0[1]}), .c ({new_AGEMA_signal_897, y_rotated23[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_10_U1 ( .s (round[0]), .b ({y_round_in_s1[10], y_round_in_s0[10]}), .a ({y_round_in_s1[2], y_round_in_s0[2]}), .c ({new_AGEMA_signal_898, y_rotated23[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_11_U1 ( .s (round[0]), .b ({y_round_in_s1[11], y_round_in_s0[11]}), .a ({y_round_in_s1[3], y_round_in_s0[3]}), .c ({new_AGEMA_signal_899, y_rotated23[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_12_U1 ( .s (round[0]), .b ({y_round_in_s1[12], y_round_in_s0[12]}), .a ({y_round_in_s1[4], y_round_in_s0[4]}), .c ({new_AGEMA_signal_900, y_rotated23[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_13_U1 ( .s (round[0]), .b ({y_round_in_s1[13], y_round_in_s0[13]}), .a ({y_round_in_s1[5], y_round_in_s0[5]}), .c ({new_AGEMA_signal_901, y_rotated23[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_14_U1 ( .s (round[0]), .b ({y_round_in_s1[14], y_round_in_s0[14]}), .a ({y_round_in_s1[6], y_round_in_s0[6]}), .c ({new_AGEMA_signal_902, y_rotated23[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_15_U1 ( .s (round[0]), .b ({y_round_in_s1[15], y_round_in_s0[15]}), .a ({y_round_in_s1[7], y_round_in_s0[7]}), .c ({new_AGEMA_signal_903, y_rotated23[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_16_U1 ( .s (round[0]), .b ({y_round_in_s1[16], y_round_in_s0[16]}), .a ({y_round_in_s1[8], y_round_in_s0[8]}), .c ({new_AGEMA_signal_904, y_rotated23[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_17_U1 ( .s (round[0]), .b ({y_round_in_s1[17], y_round_in_s0[17]}), .a ({y_round_in_s1[9], y_round_in_s0[9]}), .c ({new_AGEMA_signal_905, y_rotated23[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_18_U1 ( .s (round[0]), .b ({y_round_in_s1[18], y_round_in_s0[18]}), .a ({y_round_in_s1[10], y_round_in_s0[10]}), .c ({new_AGEMA_signal_906, y_rotated23[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_19_U1 ( .s (round[0]), .b ({y_round_in_s1[19], y_round_in_s0[19]}), .a ({y_round_in_s1[11], y_round_in_s0[11]}), .c ({new_AGEMA_signal_907, y_rotated23[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_20_U1 ( .s (round[0]), .b ({y_round_in_s1[20], y_round_in_s0[20]}), .a ({y_round_in_s1[12], y_round_in_s0[12]}), .c ({new_AGEMA_signal_908, y_rotated23[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_21_U1 ( .s (round[0]), .b ({y_round_in_s1[21], y_round_in_s0[21]}), .a ({y_round_in_s1[13], y_round_in_s0[13]}), .c ({new_AGEMA_signal_909, y_rotated23[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_22_U1 ( .s (round[0]), .b ({y_round_in_s1[22], y_round_in_s0[22]}), .a ({y_round_in_s1[14], y_round_in_s0[14]}), .c ({new_AGEMA_signal_910, y_rotated23[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_23_U1 ( .s (round[0]), .b ({y_round_in_s1[23], y_round_in_s0[23]}), .a ({y_round_in_s1[15], y_round_in_s0[15]}), .c ({new_AGEMA_signal_911, y_rotated23[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_24_U1 ( .s (round[0]), .b ({y_round_in_s1[24], y_round_in_s0[24]}), .a ({y_round_in_s1[16], y_round_in_s0[16]}), .c ({new_AGEMA_signal_912, y_rotated23[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_25_U1 ( .s (round[0]), .b ({y_round_in_s1[25], y_round_in_s0[25]}), .a ({y_round_in_s1[17], y_round_in_s0[17]}), .c ({new_AGEMA_signal_913, y_rotated23[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_26_U1 ( .s (round[0]), .b ({y_round_in_s1[26], y_round_in_s0[26]}), .a ({y_round_in_s1[18], y_round_in_s0[18]}), .c ({new_AGEMA_signal_914, y_rotated23[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_27_U1 ( .s (round[0]), .b ({y_round_in_s1[27], y_round_in_s0[27]}), .a ({y_round_in_s1[19], y_round_in_s0[19]}), .c ({new_AGEMA_signal_915, y_rotated23[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_28_U1 ( .s (round[0]), .b ({y_round_in_s1[28], y_round_in_s0[28]}), .a ({y_round_in_s1[20], y_round_in_s0[20]}), .c ({new_AGEMA_signal_916, y_rotated23[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_29_U1 ( .s (round[0]), .b ({y_round_in_s1[29], y_round_in_s0[29]}), .a ({y_round_in_s1[21], y_round_in_s0[21]}), .c ({new_AGEMA_signal_917, y_rotated23[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_30_U1 ( .s (round[0]), .b ({y_round_in_s1[30], y_round_in_s0[30]}), .a ({y_round_in_s1[22], y_round_in_s0[22]}), .c ({new_AGEMA_signal_918, y_rotated23[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M1_mux_inst_31_U1 ( .s (round[0]), .b ({y_round_in_s1[31], y_round_in_s0[31]}), .a ({y_round_in_s1[23], y_round_in_s0[23]}), .c ({new_AGEMA_signal_919, y_rotated23[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_0_U1 ( .s (round[1]), .b ({new_AGEMA_signal_826, y_rotated01[0]}), .a ({new_AGEMA_signal_888, y_rotated23[0]}), .c ({new_AGEMA_signal_920, y_rotated[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_1_U1 ( .s (round[1]), .b ({new_AGEMA_signal_829, y_rotated01[1]}), .a ({new_AGEMA_signal_889, y_rotated23[1]}), .c ({new_AGEMA_signal_921, y_rotated[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_2_U1 ( .s (round[1]), .b ({new_AGEMA_signal_832, y_rotated01[2]}), .a ({new_AGEMA_signal_890, y_rotated23[2]}), .c ({new_AGEMA_signal_922, y_rotated[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_3_U1 ( .s (round[1]), .b ({new_AGEMA_signal_835, y_rotated01[3]}), .a ({new_AGEMA_signal_891, y_rotated23[3]}), .c ({new_AGEMA_signal_923, y_rotated[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_4_U1 ( .s (round[1]), .b ({new_AGEMA_signal_838, y_rotated01[4]}), .a ({new_AGEMA_signal_892, y_rotated23[4]}), .c ({new_AGEMA_signal_924, y_rotated[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_5_U1 ( .s (round[1]), .b ({new_AGEMA_signal_841, y_rotated01[5]}), .a ({new_AGEMA_signal_893, y_rotated23[5]}), .c ({new_AGEMA_signal_925, y_rotated[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_6_U1 ( .s (round[1]), .b ({new_AGEMA_signal_844, y_rotated01[6]}), .a ({new_AGEMA_signal_894, y_rotated23[6]}), .c ({new_AGEMA_signal_926, y_rotated[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_7_U1 ( .s (round[1]), .b ({new_AGEMA_signal_847, y_rotated01[7]}), .a ({new_AGEMA_signal_895, y_rotated23[7]}), .c ({new_AGEMA_signal_927, y_rotated[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_8_U1 ( .s (round[1]), .b ({new_AGEMA_signal_850, y_rotated01[8]}), .a ({new_AGEMA_signal_896, y_rotated23[8]}), .c ({new_AGEMA_signal_928, y_rotated[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_9_U1 ( .s (round[1]), .b ({new_AGEMA_signal_853, y_rotated01[9]}), .a ({new_AGEMA_signal_897, y_rotated23[9]}), .c ({new_AGEMA_signal_929, y_rotated[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_10_U1 ( .s (round[1]), .b ({new_AGEMA_signal_856, y_rotated01[10]}), .a ({new_AGEMA_signal_898, y_rotated23[10]}), .c ({new_AGEMA_signal_930, y_rotated[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_11_U1 ( .s (round[1]), .b ({new_AGEMA_signal_859, y_rotated01[11]}), .a ({new_AGEMA_signal_899, y_rotated23[11]}), .c ({new_AGEMA_signal_931, y_rotated[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_12_U1 ( .s (round[1]), .b ({new_AGEMA_signal_862, y_rotated01[12]}), .a ({new_AGEMA_signal_900, y_rotated23[12]}), .c ({new_AGEMA_signal_932, y_rotated[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_13_U1 ( .s (round[1]), .b ({new_AGEMA_signal_865, y_rotated01[13]}), .a ({new_AGEMA_signal_901, y_rotated23[13]}), .c ({new_AGEMA_signal_933, y_rotated[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_14_U1 ( .s (round[1]), .b ({new_AGEMA_signal_867, y_rotated01[14]}), .a ({new_AGEMA_signal_902, y_rotated23[14]}), .c ({new_AGEMA_signal_934, y_rotated[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_15_U1 ( .s (round[1]), .b ({new_AGEMA_signal_869, y_rotated01[15]}), .a ({new_AGEMA_signal_903, y_rotated23[15]}), .c ({new_AGEMA_signal_935, y_rotated[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_16_U1 ( .s (round[1]), .b ({new_AGEMA_signal_871, y_rotated01[16]}), .a ({new_AGEMA_signal_904, y_rotated23[16]}), .c ({new_AGEMA_signal_936, y_rotated[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_17_U1 ( .s (round[1]), .b ({new_AGEMA_signal_873, y_rotated01[17]}), .a ({new_AGEMA_signal_905, y_rotated23[17]}), .c ({new_AGEMA_signal_937, y_rotated[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_18_U1 ( .s (round[1]), .b ({new_AGEMA_signal_874, y_rotated01[18]}), .a ({new_AGEMA_signal_906, y_rotated23[18]}), .c ({new_AGEMA_signal_938, y_rotated[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_19_U1 ( .s (round[1]), .b ({new_AGEMA_signal_875, y_rotated01[19]}), .a ({new_AGEMA_signal_907, y_rotated23[19]}), .c ({new_AGEMA_signal_939, y_rotated[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_20_U1 ( .s (round[1]), .b ({new_AGEMA_signal_876, y_rotated01[20]}), .a ({new_AGEMA_signal_908, y_rotated23[20]}), .c ({new_AGEMA_signal_940, y_rotated[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_21_U1 ( .s (round[1]), .b ({new_AGEMA_signal_877, y_rotated01[21]}), .a ({new_AGEMA_signal_909, y_rotated23[21]}), .c ({new_AGEMA_signal_941, y_rotated[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_22_U1 ( .s (round[1]), .b ({new_AGEMA_signal_878, y_rotated01[22]}), .a ({new_AGEMA_signal_910, y_rotated23[22]}), .c ({new_AGEMA_signal_942, y_rotated[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_23_U1 ( .s (round[1]), .b ({new_AGEMA_signal_879, y_rotated01[23]}), .a ({new_AGEMA_signal_911, y_rotated23[23]}), .c ({new_AGEMA_signal_943, y_rotated[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_24_U1 ( .s (round[1]), .b ({new_AGEMA_signal_880, y_rotated01[24]}), .a ({new_AGEMA_signal_912, y_rotated23[24]}), .c ({new_AGEMA_signal_944, y_rotated[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_25_U1 ( .s (round[1]), .b ({new_AGEMA_signal_881, y_rotated01[25]}), .a ({new_AGEMA_signal_913, y_rotated23[25]}), .c ({new_AGEMA_signal_945, y_rotated[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_26_U1 ( .s (round[1]), .b ({new_AGEMA_signal_882, y_rotated01[26]}), .a ({new_AGEMA_signal_914, y_rotated23[26]}), .c ({new_AGEMA_signal_946, y_rotated[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_27_U1 ( .s (round[1]), .b ({new_AGEMA_signal_883, y_rotated01[27]}), .a ({new_AGEMA_signal_915, y_rotated23[27]}), .c ({new_AGEMA_signal_947, y_rotated[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_28_U1 ( .s (round[1]), .b ({new_AGEMA_signal_884, y_rotated01[28]}), .a ({new_AGEMA_signal_916, y_rotated23[28]}), .c ({new_AGEMA_signal_948, y_rotated[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_29_U1 ( .s (round[1]), .b ({new_AGEMA_signal_885, y_rotated01[29]}), .a ({new_AGEMA_signal_917, y_rotated23[29]}), .c ({new_AGEMA_signal_949, y_rotated[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_30_U1 ( .s (round[1]), .b ({new_AGEMA_signal_886, y_rotated01[30]}), .a ({new_AGEMA_signal_918, y_rotated23[30]}), .c ({new_AGEMA_signal_950, y_rotated[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M3_mux_inst_31_U1 ( .s (round[1]), .b ({new_AGEMA_signal_887, y_rotated01[31]}), .a ({new_AGEMA_signal_919, y_rotated23[31]}), .c ({new_AGEMA_signal_951, y_rotated[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_0_U1 ( .a ({x_round_in_s1[0], x_round_in_s0[0]}), .b ({new_AGEMA_signal_920, y_rotated[0]}), .c ({new_AGEMA_signal_953, sum[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_1_U1 ( .a ({x_round_in_s1[1], x_round_in_s0[1]}), .b ({new_AGEMA_signal_921, y_rotated[1]}), .c ({new_AGEMA_signal_956, AdderIns_p6[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_2_U1 ( .a ({x_round_in_s1[2], x_round_in_s0[2]}), .b ({new_AGEMA_signal_922, y_rotated[2]}), .c ({new_AGEMA_signal_959, AdderIns_p6[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_3_U1 ( .a ({x_round_in_s1[3], x_round_in_s0[3]}), .b ({new_AGEMA_signal_923, y_rotated[3]}), .c ({new_AGEMA_signal_962, AdderIns_p6[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_4_U1 ( .a ({x_round_in_s1[4], x_round_in_s0[4]}), .b ({new_AGEMA_signal_924, y_rotated[4]}), .c ({new_AGEMA_signal_965, AdderIns_p6[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_5_U1 ( .a ({x_round_in_s1[5], x_round_in_s0[5]}), .b ({new_AGEMA_signal_925, y_rotated[5]}), .c ({new_AGEMA_signal_968, AdderIns_p6[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_6_U1 ( .a ({x_round_in_s1[6], x_round_in_s0[6]}), .b ({new_AGEMA_signal_926, y_rotated[6]}), .c ({new_AGEMA_signal_971, AdderIns_p6[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_7_U1 ( .a ({x_round_in_s1[7], x_round_in_s0[7]}), .b ({new_AGEMA_signal_927, y_rotated[7]}), .c ({new_AGEMA_signal_974, AdderIns_p6[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_8_U1 ( .a ({x_round_in_s1[8], x_round_in_s0[8]}), .b ({new_AGEMA_signal_928, y_rotated[8]}), .c ({new_AGEMA_signal_977, AdderIns_p6[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_9_U1 ( .a ({x_round_in_s1[9], x_round_in_s0[9]}), .b ({new_AGEMA_signal_929, y_rotated[9]}), .c ({new_AGEMA_signal_980, AdderIns_p6[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_10_U1 ( .a ({x_round_in_s1[10], x_round_in_s0[10]}), .b ({new_AGEMA_signal_930, y_rotated[10]}), .c ({new_AGEMA_signal_983, AdderIns_p6[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_11_U1 ( .a ({x_round_in_s1[11], x_round_in_s0[11]}), .b ({new_AGEMA_signal_931, y_rotated[11]}), .c ({new_AGEMA_signal_986, AdderIns_p6[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_12_U1 ( .a ({x_round_in_s1[12], x_round_in_s0[12]}), .b ({new_AGEMA_signal_932, y_rotated[12]}), .c ({new_AGEMA_signal_989, AdderIns_p6[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_13_U1 ( .a ({x_round_in_s1[13], x_round_in_s0[13]}), .b ({new_AGEMA_signal_933, y_rotated[13]}), .c ({new_AGEMA_signal_992, AdderIns_p6[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_14_U1 ( .a ({x_round_in_s1[14], x_round_in_s0[14]}), .b ({new_AGEMA_signal_934, y_rotated[14]}), .c ({new_AGEMA_signal_995, AdderIns_p6[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_15_U1 ( .a ({x_round_in_s1[15], x_round_in_s0[15]}), .b ({new_AGEMA_signal_935, y_rotated[15]}), .c ({new_AGEMA_signal_998, AdderIns_p6[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_16_U1 ( .a ({x_round_in_s1[16], x_round_in_s0[16]}), .b ({new_AGEMA_signal_936, y_rotated[16]}), .c ({new_AGEMA_signal_1001, AdderIns_p6[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_17_U1 ( .a ({x_round_in_s1[17], x_round_in_s0[17]}), .b ({new_AGEMA_signal_937, y_rotated[17]}), .c ({new_AGEMA_signal_1004, AdderIns_p6[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_18_U1 ( .a ({x_round_in_s1[18], x_round_in_s0[18]}), .b ({new_AGEMA_signal_938, y_rotated[18]}), .c ({new_AGEMA_signal_1007, AdderIns_p6[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_19_U1 ( .a ({x_round_in_s1[19], x_round_in_s0[19]}), .b ({new_AGEMA_signal_939, y_rotated[19]}), .c ({new_AGEMA_signal_1010, AdderIns_p6[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_20_U1 ( .a ({x_round_in_s1[20], x_round_in_s0[20]}), .b ({new_AGEMA_signal_940, y_rotated[20]}), .c ({new_AGEMA_signal_1013, AdderIns_p6[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_21_U1 ( .a ({x_round_in_s1[21], x_round_in_s0[21]}), .b ({new_AGEMA_signal_941, y_rotated[21]}), .c ({new_AGEMA_signal_1016, AdderIns_p6[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_22_U1 ( .a ({x_round_in_s1[22], x_round_in_s0[22]}), .b ({new_AGEMA_signal_942, y_rotated[22]}), .c ({new_AGEMA_signal_1019, AdderIns_p6[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_23_U1 ( .a ({x_round_in_s1[23], x_round_in_s0[23]}), .b ({new_AGEMA_signal_943, y_rotated[23]}), .c ({new_AGEMA_signal_1022, AdderIns_p6[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_24_U1 ( .a ({x_round_in_s1[24], x_round_in_s0[24]}), .b ({new_AGEMA_signal_944, y_rotated[24]}), .c ({new_AGEMA_signal_1025, AdderIns_p6[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_25_U1 ( .a ({x_round_in_s1[25], x_round_in_s0[25]}), .b ({new_AGEMA_signal_945, y_rotated[25]}), .c ({new_AGEMA_signal_1028, AdderIns_p6[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_26_U1 ( .a ({x_round_in_s1[26], x_round_in_s0[26]}), .b ({new_AGEMA_signal_946, y_rotated[26]}), .c ({new_AGEMA_signal_1031, AdderIns_p6[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_27_U1 ( .a ({x_round_in_s1[27], x_round_in_s0[27]}), .b ({new_AGEMA_signal_947, y_rotated[27]}), .c ({new_AGEMA_signal_1034, AdderIns_p6[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_28_U1 ( .a ({x_round_in_s1[28], x_round_in_s0[28]}), .b ({new_AGEMA_signal_948, y_rotated[28]}), .c ({new_AGEMA_signal_1037, AdderIns_p6[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_29_U1 ( .a ({x_round_in_s1[29], x_round_in_s0[29]}), .b ({new_AGEMA_signal_949, y_rotated[29]}), .c ({new_AGEMA_signal_1040, AdderIns_p6[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_30_U1 ( .a ({x_round_in_s1[30], x_round_in_s0[30]}), .b ({new_AGEMA_signal_950, y_rotated[30]}), .c ({new_AGEMA_signal_1043, AdderIns_p6[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_31_U1 ( .a ({x_round_in_s1[31], x_round_in_s0[31]}), .b ({new_AGEMA_signal_951, y_rotated[31]}), .c ({new_AGEMA_signal_1046, AdderIns_p6[31]}) ) ;
    //ClockGatingController #(10) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) U140 ( .a ({1'b0, round_constant[1]}), .b ({new_AGEMA_signal_1225, sum[1]}), .c ({x_round_out_s1[1], x_round_out_s0[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_0_a1_U1 ( .a ({x_round_in_s1[0], x_round_in_s0[0]}), .b ({new_AGEMA_signal_920, y_rotated[0]}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_954, AdderIns_g1[0]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_1_a1_U1 ( .a ({x_round_in_s1[1], x_round_in_s0[1]}), .b ({new_AGEMA_signal_921, y_rotated[1]}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_957, AdderIns_g1[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_2_a1_U1 ( .a ({x_round_in_s1[2], x_round_in_s0[2]}), .b ({new_AGEMA_signal_922, y_rotated[2]}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_960, AdderIns_g1[2]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_3_a1_U1 ( .a ({x_round_in_s1[3], x_round_in_s0[3]}), .b ({new_AGEMA_signal_923, y_rotated[3]}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_963, AdderIns_g1[3]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_4_a1_U1 ( .a ({x_round_in_s1[4], x_round_in_s0[4]}), .b ({new_AGEMA_signal_924, y_rotated[4]}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_966, AdderIns_g1[4]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_5_a1_U1 ( .a ({x_round_in_s1[5], x_round_in_s0[5]}), .b ({new_AGEMA_signal_925, y_rotated[5]}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_969, AdderIns_g1[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_6_a1_U1 ( .a ({x_round_in_s1[6], x_round_in_s0[6]}), .b ({new_AGEMA_signal_926, y_rotated[6]}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_972, AdderIns_g1[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_7_a1_U1 ( .a ({x_round_in_s1[7], x_round_in_s0[7]}), .b ({new_AGEMA_signal_927, y_rotated[7]}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_975, AdderIns_g1[7]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_8_a1_U1 ( .a ({x_round_in_s1[8], x_round_in_s0[8]}), .b ({new_AGEMA_signal_928, y_rotated[8]}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_978, AdderIns_g1[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_9_a1_U1 ( .a ({x_round_in_s1[9], x_round_in_s0[9]}), .b ({new_AGEMA_signal_929, y_rotated[9]}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_981, AdderIns_g1[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_10_a1_U1 ( .a ({x_round_in_s1[10], x_round_in_s0[10]}), .b ({new_AGEMA_signal_930, y_rotated[10]}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_984, AdderIns_g1[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_11_a1_U1 ( .a ({x_round_in_s1[11], x_round_in_s0[11]}), .b ({new_AGEMA_signal_931, y_rotated[11]}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_987, AdderIns_g1[11]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_12_a1_U1 ( .a ({x_round_in_s1[12], x_round_in_s0[12]}), .b ({new_AGEMA_signal_932, y_rotated[12]}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_990, AdderIns_g1[12]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_13_a1_U1 ( .a ({x_round_in_s1[13], x_round_in_s0[13]}), .b ({new_AGEMA_signal_933, y_rotated[13]}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_993, AdderIns_g1[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_14_a1_U1 ( .a ({x_round_in_s1[14], x_round_in_s0[14]}), .b ({new_AGEMA_signal_934, y_rotated[14]}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_996, AdderIns_g1[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_15_a1_U1 ( .a ({x_round_in_s1[15], x_round_in_s0[15]}), .b ({new_AGEMA_signal_935, y_rotated[15]}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_999, AdderIns_g1[15]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_16_a1_U1 ( .a ({x_round_in_s1[16], x_round_in_s0[16]}), .b ({new_AGEMA_signal_936, y_rotated[16]}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_1002, AdderIns_g1[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_17_a1_U1 ( .a ({x_round_in_s1[17], x_round_in_s0[17]}), .b ({new_AGEMA_signal_937, y_rotated[17]}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_1005, AdderIns_g1[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_18_a1_U1 ( .a ({x_round_in_s1[18], x_round_in_s0[18]}), .b ({new_AGEMA_signal_938, y_rotated[18]}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_1008, AdderIns_g1[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_19_a1_U1 ( .a ({x_round_in_s1[19], x_round_in_s0[19]}), .b ({new_AGEMA_signal_939, y_rotated[19]}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_1011, AdderIns_g1[19]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_20_a1_U1 ( .a ({x_round_in_s1[20], x_round_in_s0[20]}), .b ({new_AGEMA_signal_940, y_rotated[20]}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_1014, AdderIns_g1[20]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_21_a1_U1 ( .a ({x_round_in_s1[21], x_round_in_s0[21]}), .b ({new_AGEMA_signal_941, y_rotated[21]}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_1017, AdderIns_g1[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_22_a1_U1 ( .a ({x_round_in_s1[22], x_round_in_s0[22]}), .b ({new_AGEMA_signal_942, y_rotated[22]}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_1020, AdderIns_g1[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_23_a1_U1 ( .a ({x_round_in_s1[23], x_round_in_s0[23]}), .b ({new_AGEMA_signal_943, y_rotated[23]}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_1023, AdderIns_g1[23]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_24_a1_U1 ( .a ({x_round_in_s1[24], x_round_in_s0[24]}), .b ({new_AGEMA_signal_944, y_rotated[24]}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_1026, AdderIns_g1[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_25_a1_U1 ( .a ({x_round_in_s1[25], x_round_in_s0[25]}), .b ({new_AGEMA_signal_945, y_rotated[25]}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_1029, AdderIns_g1[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_26_a1_U1 ( .a ({x_round_in_s1[26], x_round_in_s0[26]}), .b ({new_AGEMA_signal_946, y_rotated[26]}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_1032, AdderIns_g1[26]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_27_a1_U1 ( .a ({x_round_in_s1[27], x_round_in_s0[27]}), .b ({new_AGEMA_signal_947, y_rotated[27]}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_1035, AdderIns_g1[27]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_28_a1_U1 ( .a ({x_round_in_s1[28], x_round_in_s0[28]}), .b ({new_AGEMA_signal_948, y_rotated[28]}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_1038, AdderIns_g1[28]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_29_a1_U1 ( .a ({x_round_in_s1[29], x_round_in_s0[29]}), .b ({new_AGEMA_signal_949, y_rotated[29]}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_1041, AdderIns_g1[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s1_pg_30_a1_U1 ( .a ({x_round_in_s1[30], x_round_in_s0[30]}), .b ({new_AGEMA_signal_950, y_rotated[30]}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_1044, AdderIns_g1[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_gc_0_a1_U1 ( .a ({new_AGEMA_signal_954, AdderIns_g1[0]}), .b ({new_AGEMA_signal_1048, AdderIns_s2_gc_0_a1_t}), .c ({new_AGEMA_signal_1109, AdderIns_g6[0]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_953, sum[0]}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_1048, AdderIns_s2_gc_0_a1_t}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_0_a2_U1 ( .a ({new_AGEMA_signal_953, sum[0]}), .b ({new_AGEMA_signal_956, AdderIns_p6[1]}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_1050, AdderIns_p2[0]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_1_a2_U1 ( .a ({new_AGEMA_signal_956, AdderIns_p6[1]}), .b ({new_AGEMA_signal_959, AdderIns_p6[2]}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_1052, AdderIns_p2[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_2_a2_U1 ( .a ({new_AGEMA_signal_959, AdderIns_p6[2]}), .b ({new_AGEMA_signal_962, AdderIns_p6[3]}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_1054, AdderIns_p2[2]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_3_a2_U1 ( .a ({new_AGEMA_signal_962, AdderIns_p6[3]}), .b ({new_AGEMA_signal_965, AdderIns_p6[4]}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_1056, AdderIns_p2[3]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_4_a2_U1 ( .a ({new_AGEMA_signal_965, AdderIns_p6[4]}), .b ({new_AGEMA_signal_968, AdderIns_p6[5]}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_1058, AdderIns_p2[4]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_5_a2_U1 ( .a ({new_AGEMA_signal_968, AdderIns_p6[5]}), .b ({new_AGEMA_signal_971, AdderIns_p6[6]}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_1060, AdderIns_p2[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_6_a2_U1 ( .a ({new_AGEMA_signal_971, AdderIns_p6[6]}), .b ({new_AGEMA_signal_974, AdderIns_p6[7]}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_1062, AdderIns_p2[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_7_a2_U1 ( .a ({new_AGEMA_signal_974, AdderIns_p6[7]}), .b ({new_AGEMA_signal_977, AdderIns_p6[8]}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_1064, AdderIns_p2[7]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_8_a2_U1 ( .a ({new_AGEMA_signal_977, AdderIns_p6[8]}), .b ({new_AGEMA_signal_980, AdderIns_p6[9]}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_1066, AdderIns_p2[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_9_a2_U1 ( .a ({new_AGEMA_signal_980, AdderIns_p6[9]}), .b ({new_AGEMA_signal_983, AdderIns_p6[10]}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_1068, AdderIns_p2[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_10_a2_U1 ( .a ({new_AGEMA_signal_983, AdderIns_p6[10]}), .b ({new_AGEMA_signal_986, AdderIns_p6[11]}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_1070, AdderIns_p2[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_11_a2_U1 ( .a ({new_AGEMA_signal_986, AdderIns_p6[11]}), .b ({new_AGEMA_signal_989, AdderIns_p6[12]}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_1072, AdderIns_p2[11]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_12_a2_U1 ( .a ({new_AGEMA_signal_989, AdderIns_p6[12]}), .b ({new_AGEMA_signal_992, AdderIns_p6[13]}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_1074, AdderIns_p2[12]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_13_a2_U1 ( .a ({new_AGEMA_signal_992, AdderIns_p6[13]}), .b ({new_AGEMA_signal_995, AdderIns_p6[14]}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_1076, AdderIns_p2[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_14_a2_U1 ( .a ({new_AGEMA_signal_995, AdderIns_p6[14]}), .b ({new_AGEMA_signal_998, AdderIns_p6[15]}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_1078, AdderIns_p2[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_15_a2_U1 ( .a ({new_AGEMA_signal_998, AdderIns_p6[15]}), .b ({new_AGEMA_signal_1001, AdderIns_p6[16]}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_1080, AdderIns_p2[15]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_16_a2_U1 ( .a ({new_AGEMA_signal_1001, AdderIns_p6[16]}), .b ({new_AGEMA_signal_1004, AdderIns_p6[17]}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_1082, AdderIns_p2[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_17_a2_U1 ( .a ({new_AGEMA_signal_1004, AdderIns_p6[17]}), .b ({new_AGEMA_signal_1007, AdderIns_p6[18]}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_1084, AdderIns_p2[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_18_a2_U1 ( .a ({new_AGEMA_signal_1007, AdderIns_p6[18]}), .b ({new_AGEMA_signal_1010, AdderIns_p6[19]}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_1086, AdderIns_p2[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_19_a2_U1 ( .a ({new_AGEMA_signal_1010, AdderIns_p6[19]}), .b ({new_AGEMA_signal_1013, AdderIns_p6[20]}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_1088, AdderIns_p2[19]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_20_a2_U1 ( .a ({new_AGEMA_signal_1013, AdderIns_p6[20]}), .b ({new_AGEMA_signal_1016, AdderIns_p6[21]}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_1090, AdderIns_p2[20]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_21_a2_U1 ( .a ({new_AGEMA_signal_1016, AdderIns_p6[21]}), .b ({new_AGEMA_signal_1019, AdderIns_p6[22]}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_1092, AdderIns_p2[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_22_a2_U1 ( .a ({new_AGEMA_signal_1019, AdderIns_p6[22]}), .b ({new_AGEMA_signal_1022, AdderIns_p6[23]}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_1094, AdderIns_p2[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_23_a2_U1 ( .a ({new_AGEMA_signal_1022, AdderIns_p6[23]}), .b ({new_AGEMA_signal_1025, AdderIns_p6[24]}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_1096, AdderIns_p2[23]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_24_a2_U1 ( .a ({new_AGEMA_signal_1025, AdderIns_p6[24]}), .b ({new_AGEMA_signal_1028, AdderIns_p6[25]}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_1098, AdderIns_p2[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_25_a2_U1 ( .a ({new_AGEMA_signal_1028, AdderIns_p6[25]}), .b ({new_AGEMA_signal_1031, AdderIns_p6[26]}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_1100, AdderIns_p2[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_26_a2_U1 ( .a ({new_AGEMA_signal_1031, AdderIns_p6[26]}), .b ({new_AGEMA_signal_1034, AdderIns_p6[27]}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_1102, AdderIns_p2[26]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_27_a2_U1 ( .a ({new_AGEMA_signal_1034, AdderIns_p6[27]}), .b ({new_AGEMA_signal_1037, AdderIns_p6[28]}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_1104, AdderIns_p2[27]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_28_a2_U1 ( .a ({new_AGEMA_signal_1037, AdderIns_p6[28]}), .b ({new_AGEMA_signal_1040, AdderIns_p6[29]}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_1106, AdderIns_p2[28]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_29_a2_U1 ( .a ({new_AGEMA_signal_1040, AdderIns_p6[29]}), .b ({new_AGEMA_signal_1043, AdderIns_p6[30]}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_1108, AdderIns_p2[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U11 ( .a ({new_AGEMA_signal_1109, AdderIns_g6[0]}), .b ({new_AGEMA_signal_956, AdderIns_p6[1]}), .c ({new_AGEMA_signal_1225, sum[1]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) U151 ( .a ({1'b0, round_constant[2]}), .b ({new_AGEMA_signal_1275, sum[2]}), .c ({x_round_out_s1[2], x_round_out_s0[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U154 ( .a ({1'b0, round_constant[3]}), .b ({new_AGEMA_signal_1309, sum[3]}), .c ({x_round_out_s1[3], x_round_out_s0[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_0_a1_U1 ( .a ({new_AGEMA_signal_957, AdderIns_g1[1]}), .b ({new_AGEMA_signal_1049, AdderIns_s2_bc_0_a1_t}), .c ({new_AGEMA_signal_1110, AdderIns_g2[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_954, AdderIns_g1[0]}), .b ({new_AGEMA_signal_956, AdderIns_p6[1]}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_1049, AdderIns_s2_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_1_a1_U1 ( .a ({new_AGEMA_signal_960, AdderIns_g1[2]}), .b ({new_AGEMA_signal_1051, AdderIns_s2_bc_1_a1_t}), .c ({new_AGEMA_signal_1111, AdderIns_g2[2]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_957, AdderIns_g1[1]}), .b ({new_AGEMA_signal_959, AdderIns_p6[2]}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_1051, AdderIns_s2_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_2_a1_U1 ( .a ({new_AGEMA_signal_963, AdderIns_g1[3]}), .b ({new_AGEMA_signal_1053, AdderIns_s2_bc_2_a1_t}), .c ({new_AGEMA_signal_1112, AdderIns_g2[3]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_960, AdderIns_g1[2]}), .b ({new_AGEMA_signal_962, AdderIns_p6[3]}), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_1053, AdderIns_s2_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_3_a1_U1 ( .a ({new_AGEMA_signal_966, AdderIns_g1[4]}), .b ({new_AGEMA_signal_1055, AdderIns_s2_bc_3_a1_t}), .c ({new_AGEMA_signal_1113, AdderIns_g2[4]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_963, AdderIns_g1[3]}), .b ({new_AGEMA_signal_965, AdderIns_p6[4]}), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_1055, AdderIns_s2_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_4_a1_U1 ( .a ({new_AGEMA_signal_969, AdderIns_g1[5]}), .b ({new_AGEMA_signal_1057, AdderIns_s2_bc_4_a1_t}), .c ({new_AGEMA_signal_1114, AdderIns_g2[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_966, AdderIns_g1[4]}), .b ({new_AGEMA_signal_968, AdderIns_p6[5]}), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_1057, AdderIns_s2_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_5_a1_U1 ( .a ({new_AGEMA_signal_972, AdderIns_g1[6]}), .b ({new_AGEMA_signal_1059, AdderIns_s2_bc_5_a1_t}), .c ({new_AGEMA_signal_1115, AdderIns_g2[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_969, AdderIns_g1[5]}), .b ({new_AGEMA_signal_971, AdderIns_p6[6]}), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_1059, AdderIns_s2_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_6_a1_U1 ( .a ({new_AGEMA_signal_975, AdderIns_g1[7]}), .b ({new_AGEMA_signal_1061, AdderIns_s2_bc_6_a1_t}), .c ({new_AGEMA_signal_1116, AdderIns_g2[7]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_972, AdderIns_g1[6]}), .b ({new_AGEMA_signal_974, AdderIns_p6[7]}), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_1061, AdderIns_s2_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_7_a1_U1 ( .a ({new_AGEMA_signal_978, AdderIns_g1[8]}), .b ({new_AGEMA_signal_1063, AdderIns_s2_bc_7_a1_t}), .c ({new_AGEMA_signal_1117, AdderIns_g2[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_975, AdderIns_g1[7]}), .b ({new_AGEMA_signal_977, AdderIns_p6[8]}), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_1063, AdderIns_s2_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_8_a1_U1 ( .a ({new_AGEMA_signal_981, AdderIns_g1[9]}), .b ({new_AGEMA_signal_1065, AdderIns_s2_bc_8_a1_t}), .c ({new_AGEMA_signal_1118, AdderIns_g2[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_978, AdderIns_g1[8]}), .b ({new_AGEMA_signal_980, AdderIns_p6[9]}), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_1065, AdderIns_s2_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_9_a1_U1 ( .a ({new_AGEMA_signal_984, AdderIns_g1[10]}), .b ({new_AGEMA_signal_1067, AdderIns_s2_bc_9_a1_t}), .c ({new_AGEMA_signal_1119, AdderIns_g2[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_981, AdderIns_g1[9]}), .b ({new_AGEMA_signal_983, AdderIns_p6[10]}), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_1067, AdderIns_s2_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_10_a1_U1 ( .a ({new_AGEMA_signal_987, AdderIns_g1[11]}), .b ({new_AGEMA_signal_1069, AdderIns_s2_bc_10_a1_t}), .c ({new_AGEMA_signal_1120, AdderIns_g2[11]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_984, AdderIns_g1[10]}), .b ({new_AGEMA_signal_986, AdderIns_p6[11]}), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_1069, AdderIns_s2_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_11_a1_U1 ( .a ({new_AGEMA_signal_990, AdderIns_g1[12]}), .b ({new_AGEMA_signal_1071, AdderIns_s2_bc_11_a1_t}), .c ({new_AGEMA_signal_1121, AdderIns_g2[12]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_987, AdderIns_g1[11]}), .b ({new_AGEMA_signal_989, AdderIns_p6[12]}), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_1071, AdderIns_s2_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_12_a1_U1 ( .a ({new_AGEMA_signal_993, AdderIns_g1[13]}), .b ({new_AGEMA_signal_1073, AdderIns_s2_bc_12_a1_t}), .c ({new_AGEMA_signal_1122, AdderIns_g2[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_990, AdderIns_g1[12]}), .b ({new_AGEMA_signal_992, AdderIns_p6[13]}), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_1073, AdderIns_s2_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_13_a1_U1 ( .a ({new_AGEMA_signal_996, AdderIns_g1[14]}), .b ({new_AGEMA_signal_1075, AdderIns_s2_bc_13_a1_t}), .c ({new_AGEMA_signal_1123, AdderIns_g2[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_993, AdderIns_g1[13]}), .b ({new_AGEMA_signal_995, AdderIns_p6[14]}), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_1075, AdderIns_s2_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_14_a1_U1 ( .a ({new_AGEMA_signal_999, AdderIns_g1[15]}), .b ({new_AGEMA_signal_1077, AdderIns_s2_bc_14_a1_t}), .c ({new_AGEMA_signal_1124, AdderIns_g2[15]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_996, AdderIns_g1[14]}), .b ({new_AGEMA_signal_998, AdderIns_p6[15]}), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_1077, AdderIns_s2_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_15_a1_U1 ( .a ({new_AGEMA_signal_1002, AdderIns_g1[16]}), .b ({new_AGEMA_signal_1079, AdderIns_s2_bc_15_a1_t}), .c ({new_AGEMA_signal_1125, AdderIns_g2[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_999, AdderIns_g1[15]}), .b ({new_AGEMA_signal_1001, AdderIns_p6[16]}), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_1079, AdderIns_s2_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_16_a1_U1 ( .a ({new_AGEMA_signal_1005, AdderIns_g1[17]}), .b ({new_AGEMA_signal_1081, AdderIns_s2_bc_16_a1_t}), .c ({new_AGEMA_signal_1126, AdderIns_g2[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_16_a1_a1_U1 ( .a ({new_AGEMA_signal_1002, AdderIns_g1[16]}), .b ({new_AGEMA_signal_1004, AdderIns_p6[17]}), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_1081, AdderIns_s2_bc_16_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_17_a1_U1 ( .a ({new_AGEMA_signal_1008, AdderIns_g1[18]}), .b ({new_AGEMA_signal_1083, AdderIns_s2_bc_17_a1_t}), .c ({new_AGEMA_signal_1127, AdderIns_g2[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_17_a1_a1_U1 ( .a ({new_AGEMA_signal_1005, AdderIns_g1[17]}), .b ({new_AGEMA_signal_1007, AdderIns_p6[18]}), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_1083, AdderIns_s2_bc_17_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_18_a1_U1 ( .a ({new_AGEMA_signal_1011, AdderIns_g1[19]}), .b ({new_AGEMA_signal_1085, AdderIns_s2_bc_18_a1_t}), .c ({new_AGEMA_signal_1128, AdderIns_g2[19]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_18_a1_a1_U1 ( .a ({new_AGEMA_signal_1008, AdderIns_g1[18]}), .b ({new_AGEMA_signal_1010, AdderIns_p6[19]}), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_1085, AdderIns_s2_bc_18_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_19_a1_U1 ( .a ({new_AGEMA_signal_1014, AdderIns_g1[20]}), .b ({new_AGEMA_signal_1087, AdderIns_s2_bc_19_a1_t}), .c ({new_AGEMA_signal_1129, AdderIns_g2[20]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_19_a1_a1_U1 ( .a ({new_AGEMA_signal_1011, AdderIns_g1[19]}), .b ({new_AGEMA_signal_1013, AdderIns_p6[20]}), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_1087, AdderIns_s2_bc_19_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_20_a1_U1 ( .a ({new_AGEMA_signal_1017, AdderIns_g1[21]}), .b ({new_AGEMA_signal_1089, AdderIns_s2_bc_20_a1_t}), .c ({new_AGEMA_signal_1130, AdderIns_g2[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_20_a1_a1_U1 ( .a ({new_AGEMA_signal_1014, AdderIns_g1[20]}), .b ({new_AGEMA_signal_1016, AdderIns_p6[21]}), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_1089, AdderIns_s2_bc_20_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_21_a1_U1 ( .a ({new_AGEMA_signal_1020, AdderIns_g1[22]}), .b ({new_AGEMA_signal_1091, AdderIns_s2_bc_21_a1_t}), .c ({new_AGEMA_signal_1131, AdderIns_g2[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_21_a1_a1_U1 ( .a ({new_AGEMA_signal_1017, AdderIns_g1[21]}), .b ({new_AGEMA_signal_1019, AdderIns_p6[22]}), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_1091, AdderIns_s2_bc_21_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_22_a1_U1 ( .a ({new_AGEMA_signal_1023, AdderIns_g1[23]}), .b ({new_AGEMA_signal_1093, AdderIns_s2_bc_22_a1_t}), .c ({new_AGEMA_signal_1132, AdderIns_g2[23]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_22_a1_a1_U1 ( .a ({new_AGEMA_signal_1020, AdderIns_g1[22]}), .b ({new_AGEMA_signal_1022, AdderIns_p6[23]}), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_1093, AdderIns_s2_bc_22_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_23_a1_U1 ( .a ({new_AGEMA_signal_1026, AdderIns_g1[24]}), .b ({new_AGEMA_signal_1095, AdderIns_s2_bc_23_a1_t}), .c ({new_AGEMA_signal_1133, AdderIns_g2[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_23_a1_a1_U1 ( .a ({new_AGEMA_signal_1023, AdderIns_g1[23]}), .b ({new_AGEMA_signal_1025, AdderIns_p6[24]}), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_1095, AdderIns_s2_bc_23_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_24_a1_U1 ( .a ({new_AGEMA_signal_1029, AdderIns_g1[25]}), .b ({new_AGEMA_signal_1097, AdderIns_s2_bc_24_a1_t}), .c ({new_AGEMA_signal_1134, AdderIns_g2[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_24_a1_a1_U1 ( .a ({new_AGEMA_signal_1026, AdderIns_g1[24]}), .b ({new_AGEMA_signal_1028, AdderIns_p6[25]}), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_1097, AdderIns_s2_bc_24_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_25_a1_U1 ( .a ({new_AGEMA_signal_1032, AdderIns_g1[26]}), .b ({new_AGEMA_signal_1099, AdderIns_s2_bc_25_a1_t}), .c ({new_AGEMA_signal_1135, AdderIns_g2[26]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_25_a1_a1_U1 ( .a ({new_AGEMA_signal_1029, AdderIns_g1[25]}), .b ({new_AGEMA_signal_1031, AdderIns_p6[26]}), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_1099, AdderIns_s2_bc_25_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_26_a1_U1 ( .a ({new_AGEMA_signal_1035, AdderIns_g1[27]}), .b ({new_AGEMA_signal_1101, AdderIns_s2_bc_26_a1_t}), .c ({new_AGEMA_signal_1136, AdderIns_g2[27]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_26_a1_a1_U1 ( .a ({new_AGEMA_signal_1032, AdderIns_g1[26]}), .b ({new_AGEMA_signal_1034, AdderIns_p6[27]}), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_1101, AdderIns_s2_bc_26_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_27_a1_U1 ( .a ({new_AGEMA_signal_1038, AdderIns_g1[28]}), .b ({new_AGEMA_signal_1103, AdderIns_s2_bc_27_a1_t}), .c ({new_AGEMA_signal_1137, AdderIns_g2[28]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_27_a1_a1_U1 ( .a ({new_AGEMA_signal_1035, AdderIns_g1[27]}), .b ({new_AGEMA_signal_1037, AdderIns_p6[28]}), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_1103, AdderIns_s2_bc_27_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_28_a1_U1 ( .a ({new_AGEMA_signal_1041, AdderIns_g1[29]}), .b ({new_AGEMA_signal_1105, AdderIns_s2_bc_28_a1_t}), .c ({new_AGEMA_signal_1138, AdderIns_g2[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_28_a1_a1_U1 ( .a ({new_AGEMA_signal_1038, AdderIns_g1[28]}), .b ({new_AGEMA_signal_1040, AdderIns_p6[29]}), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_1105, AdderIns_s2_bc_28_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_29_a1_U1 ( .a ({new_AGEMA_signal_1044, AdderIns_g1[30]}), .b ({new_AGEMA_signal_1107, AdderIns_s2_bc_29_a1_t}), .c ({new_AGEMA_signal_1139, AdderIns_g2[30]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s2_bc_29_a1_a1_U1 ( .a ({new_AGEMA_signal_1041, AdderIns_g1[29]}), .b ({new_AGEMA_signal_1043, AdderIns_p6[30]}), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_1107, AdderIns_s2_bc_29_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_gc_0_a1_U1 ( .a ({new_AGEMA_signal_1110, AdderIns_g2[1]}), .b ({new_AGEMA_signal_1140, AdderIns_s3_gc_0_a1_t}), .c ({new_AGEMA_signal_1169, AdderIns_g6[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1050, AdderIns_p2[0]}), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_1140, AdderIns_s3_gc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_gc_1_a1_U1 ( .a ({new_AGEMA_signal_1111, AdderIns_g2[2]}), .b ({new_AGEMA_signal_1170, AdderIns_s3_gc_1_a1_t}), .c ({new_AGEMA_signal_1227, AdderIns_g6[2]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1109, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1052, AdderIns_p2[1]}), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_1170, AdderIns_s3_gc_1_a1_t}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_0_a2_U1 ( .a ({new_AGEMA_signal_1050, AdderIns_p2[0]}), .b ({new_AGEMA_signal_1054, AdderIns_p2[2]}), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_1141, AdderIns_p3[0]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1052, AdderIns_p2[1]}), .b ({new_AGEMA_signal_1056, AdderIns_p2[3]}), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_1142, AdderIns_p3[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1054, AdderIns_p2[2]}), .b ({new_AGEMA_signal_1058, AdderIns_p2[4]}), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_1143, AdderIns_p3[2]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1056, AdderIns_p2[3]}), .b ({new_AGEMA_signal_1060, AdderIns_p2[5]}), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_1144, AdderIns_p3[3]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1058, AdderIns_p2[4]}), .b ({new_AGEMA_signal_1062, AdderIns_p2[6]}), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_1145, AdderIns_p3[4]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1060, AdderIns_p2[5]}), .b ({new_AGEMA_signal_1064, AdderIns_p2[7]}), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_1146, AdderIns_p3[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1062, AdderIns_p2[6]}), .b ({new_AGEMA_signal_1066, AdderIns_p2[8]}), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_1147, AdderIns_p3[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1064, AdderIns_p2[7]}), .b ({new_AGEMA_signal_1068, AdderIns_p2[9]}), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_1148, AdderIns_p3[7]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1066, AdderIns_p2[8]}), .b ({new_AGEMA_signal_1070, AdderIns_p2[10]}), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_1149, AdderIns_p3[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1068, AdderIns_p2[9]}), .b ({new_AGEMA_signal_1072, AdderIns_p2[11]}), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_1150, AdderIns_p3[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1070, AdderIns_p2[10]}), .b ({new_AGEMA_signal_1074, AdderIns_p2[12]}), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_1151, AdderIns_p3[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1072, AdderIns_p2[11]}), .b ({new_AGEMA_signal_1076, AdderIns_p2[13]}), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_1152, AdderIns_p3[11]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1074, AdderIns_p2[12]}), .b ({new_AGEMA_signal_1078, AdderIns_p2[14]}), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_1153, AdderIns_p3[12]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1076, AdderIns_p2[13]}), .b ({new_AGEMA_signal_1080, AdderIns_p2[15]}), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_1154, AdderIns_p3[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1078, AdderIns_p2[14]}), .b ({new_AGEMA_signal_1082, AdderIns_p2[16]}), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_1155, AdderIns_p3[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_15_a2_U1 ( .a ({new_AGEMA_signal_1080, AdderIns_p2[15]}), .b ({new_AGEMA_signal_1084, AdderIns_p2[17]}), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_1156, AdderIns_p3[15]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_16_a2_U1 ( .a ({new_AGEMA_signal_1082, AdderIns_p2[16]}), .b ({new_AGEMA_signal_1086, AdderIns_p2[18]}), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_1157, AdderIns_p3[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_17_a2_U1 ( .a ({new_AGEMA_signal_1084, AdderIns_p2[17]}), .b ({new_AGEMA_signal_1088, AdderIns_p2[19]}), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_1158, AdderIns_p3[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_18_a2_U1 ( .a ({new_AGEMA_signal_1086, AdderIns_p2[18]}), .b ({new_AGEMA_signal_1090, AdderIns_p2[20]}), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_1159, AdderIns_p3[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_19_a2_U1 ( .a ({new_AGEMA_signal_1088, AdderIns_p2[19]}), .b ({new_AGEMA_signal_1092, AdderIns_p2[21]}), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_1160, AdderIns_p3[19]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_20_a2_U1 ( .a ({new_AGEMA_signal_1090, AdderIns_p2[20]}), .b ({new_AGEMA_signal_1094, AdderIns_p2[22]}), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_1161, AdderIns_p3[20]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_21_a2_U1 ( .a ({new_AGEMA_signal_1092, AdderIns_p2[21]}), .b ({new_AGEMA_signal_1096, AdderIns_p2[23]}), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_1162, AdderIns_p3[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_22_a2_U1 ( .a ({new_AGEMA_signal_1094, AdderIns_p2[22]}), .b ({new_AGEMA_signal_1098, AdderIns_p2[24]}), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_1163, AdderIns_p3[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_23_a2_U1 ( .a ({new_AGEMA_signal_1096, AdderIns_p2[23]}), .b ({new_AGEMA_signal_1100, AdderIns_p2[25]}), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_1164, AdderIns_p3[23]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_24_a2_U1 ( .a ({new_AGEMA_signal_1098, AdderIns_p2[24]}), .b ({new_AGEMA_signal_1102, AdderIns_p2[26]}), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_1165, AdderIns_p3[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_25_a2_U1 ( .a ({new_AGEMA_signal_1100, AdderIns_p2[25]}), .b ({new_AGEMA_signal_1104, AdderIns_p2[27]}), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_1166, AdderIns_p3[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_26_a2_U1 ( .a ({new_AGEMA_signal_1102, AdderIns_p2[26]}), .b ({new_AGEMA_signal_1106, AdderIns_p2[28]}), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_1167, AdderIns_p3[26]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_27_a2_U1 ( .a ({new_AGEMA_signal_1104, AdderIns_p2[27]}), .b ({new_AGEMA_signal_1108, AdderIns_p2[29]}), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_1168, AdderIns_p3[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U25 ( .a ({new_AGEMA_signal_1227, AdderIns_g6[2]}), .b ({new_AGEMA_signal_962, AdderIns_p6[3]}), .c ({new_AGEMA_signal_1309, sum[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U22 ( .a ({new_AGEMA_signal_1169, AdderIns_g6[1]}), .b ({new_AGEMA_signal_959, AdderIns_p6[2]}), .c ({new_AGEMA_signal_1275, sum[2]}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) U155 ( .a ({1'b0, round_constant[4]}), .b ({new_AGEMA_signal_1344, sum[4]}), .c ({x_round_out_s1[4], x_round_out_s0[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U156 ( .a ({1'b0, round_constant[5]}), .b ({new_AGEMA_signal_1343, sum[5]}), .c ({x_round_out_s1[5], x_round_out_s0[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U157 ( .a ({1'b0, round_constant[6]}), .b ({new_AGEMA_signal_1342, sum[6]}), .c ({x_round_out_s1[6], x_round_out_s0[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U158 ( .a ({1'b0, round_constant[7]}), .b ({new_AGEMA_signal_1373, sum[7]}), .c ({x_round_out_s1[7], x_round_out_s0[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_0_a1_U1 ( .a ({new_AGEMA_signal_1112, AdderIns_g2[3]}), .b ({new_AGEMA_signal_1171, AdderIns_s3_bc_0_a1_t}), .c ({new_AGEMA_signal_1228, AdderIns_g3[3]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_1110, AdderIns_g2[1]}), .b ({new_AGEMA_signal_1054, AdderIns_p2[2]}), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_1171, AdderIns_s3_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_1_a1_U1 ( .a ({new_AGEMA_signal_1113, AdderIns_g2[4]}), .b ({new_AGEMA_signal_1172, AdderIns_s3_bc_1_a1_t}), .c ({new_AGEMA_signal_1229, AdderIns_g3[4]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1111, AdderIns_g2[2]}), .b ({new_AGEMA_signal_1056, AdderIns_p2[3]}), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_1172, AdderIns_s3_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_2_a1_U1 ( .a ({new_AGEMA_signal_1114, AdderIns_g2[5]}), .b ({new_AGEMA_signal_1173, AdderIns_s3_bc_2_a1_t}), .c ({new_AGEMA_signal_1230, AdderIns_g3[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1112, AdderIns_g2[3]}), .b ({new_AGEMA_signal_1058, AdderIns_p2[4]}), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_1173, AdderIns_s3_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_3_a1_U1 ( .a ({new_AGEMA_signal_1115, AdderIns_g2[6]}), .b ({new_AGEMA_signal_1174, AdderIns_s3_bc_3_a1_t}), .c ({new_AGEMA_signal_1231, AdderIns_g3[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1113, AdderIns_g2[4]}), .b ({new_AGEMA_signal_1060, AdderIns_p2[5]}), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_1174, AdderIns_s3_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_4_a1_U1 ( .a ({new_AGEMA_signal_1116, AdderIns_g2[7]}), .b ({new_AGEMA_signal_1175, AdderIns_s3_bc_4_a1_t}), .c ({new_AGEMA_signal_1232, AdderIns_g3[7]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1114, AdderIns_g2[5]}), .b ({new_AGEMA_signal_1062, AdderIns_p2[6]}), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_1175, AdderIns_s3_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_5_a1_U1 ( .a ({new_AGEMA_signal_1117, AdderIns_g2[8]}), .b ({new_AGEMA_signal_1176, AdderIns_s3_bc_5_a1_t}), .c ({new_AGEMA_signal_1233, AdderIns_g3[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1115, AdderIns_g2[6]}), .b ({new_AGEMA_signal_1064, AdderIns_p2[7]}), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_1176, AdderIns_s3_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_6_a1_U1 ( .a ({new_AGEMA_signal_1118, AdderIns_g2[9]}), .b ({new_AGEMA_signal_1177, AdderIns_s3_bc_6_a1_t}), .c ({new_AGEMA_signal_1234, AdderIns_g3[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1116, AdderIns_g2[7]}), .b ({new_AGEMA_signal_1066, AdderIns_p2[8]}), .clk (clk), .r (Fresh[128]), .c ({new_AGEMA_signal_1177, AdderIns_s3_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_7_a1_U1 ( .a ({new_AGEMA_signal_1119, AdderIns_g2[10]}), .b ({new_AGEMA_signal_1178, AdderIns_s3_bc_7_a1_t}), .c ({new_AGEMA_signal_1235, AdderIns_g3[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1117, AdderIns_g2[8]}), .b ({new_AGEMA_signal_1068, AdderIns_p2[9]}), .clk (clk), .r (Fresh[129]), .c ({new_AGEMA_signal_1178, AdderIns_s3_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_8_a1_U1 ( .a ({new_AGEMA_signal_1120, AdderIns_g2[11]}), .b ({new_AGEMA_signal_1179, AdderIns_s3_bc_8_a1_t}), .c ({new_AGEMA_signal_1236, AdderIns_g3[11]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1118, AdderIns_g2[9]}), .b ({new_AGEMA_signal_1070, AdderIns_p2[10]}), .clk (clk), .r (Fresh[130]), .c ({new_AGEMA_signal_1179, AdderIns_s3_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_9_a1_U1 ( .a ({new_AGEMA_signal_1121, AdderIns_g2[12]}), .b ({new_AGEMA_signal_1180, AdderIns_s3_bc_9_a1_t}), .c ({new_AGEMA_signal_1237, AdderIns_g3[12]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1119, AdderIns_g2[10]}), .b ({new_AGEMA_signal_1072, AdderIns_p2[11]}), .clk (clk), .r (Fresh[131]), .c ({new_AGEMA_signal_1180, AdderIns_s3_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_10_a1_U1 ( .a ({new_AGEMA_signal_1122, AdderIns_g2[13]}), .b ({new_AGEMA_signal_1181, AdderIns_s3_bc_10_a1_t}), .c ({new_AGEMA_signal_1238, AdderIns_g3[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1120, AdderIns_g2[11]}), .b ({new_AGEMA_signal_1074, AdderIns_p2[12]}), .clk (clk), .r (Fresh[132]), .c ({new_AGEMA_signal_1181, AdderIns_s3_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_11_a1_U1 ( .a ({new_AGEMA_signal_1123, AdderIns_g2[14]}), .b ({new_AGEMA_signal_1182, AdderIns_s3_bc_11_a1_t}), .c ({new_AGEMA_signal_1239, AdderIns_g3[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1121, AdderIns_g2[12]}), .b ({new_AGEMA_signal_1076, AdderIns_p2[13]}), .clk (clk), .r (Fresh[133]), .c ({new_AGEMA_signal_1182, AdderIns_s3_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_12_a1_U1 ( .a ({new_AGEMA_signal_1124, AdderIns_g2[15]}), .b ({new_AGEMA_signal_1183, AdderIns_s3_bc_12_a1_t}), .c ({new_AGEMA_signal_1240, AdderIns_g3[15]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1122, AdderIns_g2[13]}), .b ({new_AGEMA_signal_1078, AdderIns_p2[14]}), .clk (clk), .r (Fresh[134]), .c ({new_AGEMA_signal_1183, AdderIns_s3_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_13_a1_U1 ( .a ({new_AGEMA_signal_1125, AdderIns_g2[16]}), .b ({new_AGEMA_signal_1184, AdderIns_s3_bc_13_a1_t}), .c ({new_AGEMA_signal_1241, AdderIns_g3[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1123, AdderIns_g2[14]}), .b ({new_AGEMA_signal_1080, AdderIns_p2[15]}), .clk (clk), .r (Fresh[135]), .c ({new_AGEMA_signal_1184, AdderIns_s3_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_14_a1_U1 ( .a ({new_AGEMA_signal_1126, AdderIns_g2[17]}), .b ({new_AGEMA_signal_1185, AdderIns_s3_bc_14_a1_t}), .c ({new_AGEMA_signal_1242, AdderIns_g3[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1124, AdderIns_g2[15]}), .b ({new_AGEMA_signal_1082, AdderIns_p2[16]}), .clk (clk), .r (Fresh[136]), .c ({new_AGEMA_signal_1185, AdderIns_s3_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_15_a1_U1 ( .a ({new_AGEMA_signal_1127, AdderIns_g2[18]}), .b ({new_AGEMA_signal_1186, AdderIns_s3_bc_15_a1_t}), .c ({new_AGEMA_signal_1243, AdderIns_g3[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1125, AdderIns_g2[16]}), .b ({new_AGEMA_signal_1084, AdderIns_p2[17]}), .clk (clk), .r (Fresh[137]), .c ({new_AGEMA_signal_1186, AdderIns_s3_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_16_a1_U1 ( .a ({new_AGEMA_signal_1128, AdderIns_g2[19]}), .b ({new_AGEMA_signal_1187, AdderIns_s3_bc_16_a1_t}), .c ({new_AGEMA_signal_1244, AdderIns_g3[19]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_16_a1_a1_U1 ( .a ({new_AGEMA_signal_1126, AdderIns_g2[17]}), .b ({new_AGEMA_signal_1086, AdderIns_p2[18]}), .clk (clk), .r (Fresh[138]), .c ({new_AGEMA_signal_1187, AdderIns_s3_bc_16_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_17_a1_U1 ( .a ({new_AGEMA_signal_1129, AdderIns_g2[20]}), .b ({new_AGEMA_signal_1188, AdderIns_s3_bc_17_a1_t}), .c ({new_AGEMA_signal_1245, AdderIns_g3[20]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_17_a1_a1_U1 ( .a ({new_AGEMA_signal_1127, AdderIns_g2[18]}), .b ({new_AGEMA_signal_1088, AdderIns_p2[19]}), .clk (clk), .r (Fresh[139]), .c ({new_AGEMA_signal_1188, AdderIns_s3_bc_17_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_18_a1_U1 ( .a ({new_AGEMA_signal_1130, AdderIns_g2[21]}), .b ({new_AGEMA_signal_1189, AdderIns_s3_bc_18_a1_t}), .c ({new_AGEMA_signal_1246, AdderIns_g3[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_18_a1_a1_U1 ( .a ({new_AGEMA_signal_1128, AdderIns_g2[19]}), .b ({new_AGEMA_signal_1090, AdderIns_p2[20]}), .clk (clk), .r (Fresh[140]), .c ({new_AGEMA_signal_1189, AdderIns_s3_bc_18_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_19_a1_U1 ( .a ({new_AGEMA_signal_1131, AdderIns_g2[22]}), .b ({new_AGEMA_signal_1190, AdderIns_s3_bc_19_a1_t}), .c ({new_AGEMA_signal_1247, AdderIns_g3[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_19_a1_a1_U1 ( .a ({new_AGEMA_signal_1129, AdderIns_g2[20]}), .b ({new_AGEMA_signal_1092, AdderIns_p2[21]}), .clk (clk), .r (Fresh[141]), .c ({new_AGEMA_signal_1190, AdderIns_s3_bc_19_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_20_a1_U1 ( .a ({new_AGEMA_signal_1132, AdderIns_g2[23]}), .b ({new_AGEMA_signal_1191, AdderIns_s3_bc_20_a1_t}), .c ({new_AGEMA_signal_1248, AdderIns_g3[23]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_20_a1_a1_U1 ( .a ({new_AGEMA_signal_1130, AdderIns_g2[21]}), .b ({new_AGEMA_signal_1094, AdderIns_p2[22]}), .clk (clk), .r (Fresh[142]), .c ({new_AGEMA_signal_1191, AdderIns_s3_bc_20_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_21_a1_U1 ( .a ({new_AGEMA_signal_1133, AdderIns_g2[24]}), .b ({new_AGEMA_signal_1192, AdderIns_s3_bc_21_a1_t}), .c ({new_AGEMA_signal_1249, AdderIns_g3[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_21_a1_a1_U1 ( .a ({new_AGEMA_signal_1131, AdderIns_g2[22]}), .b ({new_AGEMA_signal_1096, AdderIns_p2[23]}), .clk (clk), .r (Fresh[143]), .c ({new_AGEMA_signal_1192, AdderIns_s3_bc_21_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_22_a1_U1 ( .a ({new_AGEMA_signal_1134, AdderIns_g2[25]}), .b ({new_AGEMA_signal_1193, AdderIns_s3_bc_22_a1_t}), .c ({new_AGEMA_signal_1250, AdderIns_g3[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_22_a1_a1_U1 ( .a ({new_AGEMA_signal_1132, AdderIns_g2[23]}), .b ({new_AGEMA_signal_1098, AdderIns_p2[24]}), .clk (clk), .r (Fresh[144]), .c ({new_AGEMA_signal_1193, AdderIns_s3_bc_22_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_23_a1_U1 ( .a ({new_AGEMA_signal_1135, AdderIns_g2[26]}), .b ({new_AGEMA_signal_1194, AdderIns_s3_bc_23_a1_t}), .c ({new_AGEMA_signal_1251, AdderIns_g3[26]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_23_a1_a1_U1 ( .a ({new_AGEMA_signal_1133, AdderIns_g2[24]}), .b ({new_AGEMA_signal_1100, AdderIns_p2[25]}), .clk (clk), .r (Fresh[145]), .c ({new_AGEMA_signal_1194, AdderIns_s3_bc_23_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_24_a1_U1 ( .a ({new_AGEMA_signal_1136, AdderIns_g2[27]}), .b ({new_AGEMA_signal_1195, AdderIns_s3_bc_24_a1_t}), .c ({new_AGEMA_signal_1252, AdderIns_g3[27]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_24_a1_a1_U1 ( .a ({new_AGEMA_signal_1134, AdderIns_g2[25]}), .b ({new_AGEMA_signal_1102, AdderIns_p2[26]}), .clk (clk), .r (Fresh[146]), .c ({new_AGEMA_signal_1195, AdderIns_s3_bc_24_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_25_a1_U1 ( .a ({new_AGEMA_signal_1137, AdderIns_g2[28]}), .b ({new_AGEMA_signal_1196, AdderIns_s3_bc_25_a1_t}), .c ({new_AGEMA_signal_1253, AdderIns_g3[28]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_25_a1_a1_U1 ( .a ({new_AGEMA_signal_1135, AdderIns_g2[26]}), .b ({new_AGEMA_signal_1104, AdderIns_p2[27]}), .clk (clk), .r (Fresh[147]), .c ({new_AGEMA_signal_1196, AdderIns_s3_bc_25_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_26_a1_U1 ( .a ({new_AGEMA_signal_1138, AdderIns_g2[29]}), .b ({new_AGEMA_signal_1197, AdderIns_s3_bc_26_a1_t}), .c ({new_AGEMA_signal_1254, AdderIns_g3[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_26_a1_a1_U1 ( .a ({new_AGEMA_signal_1136, AdderIns_g2[27]}), .b ({new_AGEMA_signal_1106, AdderIns_p2[28]}), .clk (clk), .r (Fresh[148]), .c ({new_AGEMA_signal_1197, AdderIns_s3_bc_26_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_27_a1_U1 ( .a ({new_AGEMA_signal_1139, AdderIns_g2[30]}), .b ({new_AGEMA_signal_1198, AdderIns_s3_bc_27_a1_t}), .c ({new_AGEMA_signal_1255, AdderIns_g3[30]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s3_bc_27_a1_a1_U1 ( .a ({new_AGEMA_signal_1137, AdderIns_g2[28]}), .b ({new_AGEMA_signal_1108, AdderIns_p2[29]}), .clk (clk), .r (Fresh[149]), .c ({new_AGEMA_signal_1198, AdderIns_s3_bc_27_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_gc_0_a1_U1 ( .a ({new_AGEMA_signal_1228, AdderIns_g3[3]}), .b ({new_AGEMA_signal_1199, AdderIns_s4_gc_0_a1_t}), .c ({new_AGEMA_signal_1277, AdderIns_g6[3]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1141, AdderIns_p3[0]}), .clk (clk), .r (Fresh[150]), .c ({new_AGEMA_signal_1199, AdderIns_s4_gc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_gc_1_a1_U1 ( .a ({new_AGEMA_signal_1229, AdderIns_g3[4]}), .b ({new_AGEMA_signal_1200, AdderIns_s4_gc_1_a1_t}), .c ({new_AGEMA_signal_1278, AdderIns_g6[4]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1109, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1142, AdderIns_p3[1]}), .clk (clk), .r (Fresh[151]), .c ({new_AGEMA_signal_1200, AdderIns_s4_gc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_gc_2_a1_U1 ( .a ({new_AGEMA_signal_1230, AdderIns_g3[5]}), .b ({new_AGEMA_signal_1256, AdderIns_s4_gc_2_a1_t}), .c ({new_AGEMA_signal_1279, AdderIns_g6[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_gc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1169, AdderIns_g6[1]}), .b ({new_AGEMA_signal_1143, AdderIns_p3[2]}), .clk (clk), .r (Fresh[152]), .c ({new_AGEMA_signal_1256, AdderIns_s4_gc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_gc_3_a1_U1 ( .a ({new_AGEMA_signal_1231, AdderIns_g3[6]}), .b ({new_AGEMA_signal_1280, AdderIns_s4_gc_3_a1_t}), .c ({new_AGEMA_signal_1311, AdderIns_g6[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_gc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1227, AdderIns_g6[2]}), .b ({new_AGEMA_signal_1144, AdderIns_p3[3]}), .clk (clk), .r (Fresh[153]), .c ({new_AGEMA_signal_1280, AdderIns_s4_gc_3_a1_t}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_0_a2_U1 ( .a ({new_AGEMA_signal_1141, AdderIns_p3[0]}), .b ({new_AGEMA_signal_1145, AdderIns_p3[4]}), .clk (clk), .r (Fresh[154]), .c ({new_AGEMA_signal_1201, AdderIns_p4[0]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1142, AdderIns_p3[1]}), .b ({new_AGEMA_signal_1146, AdderIns_p3[5]}), .clk (clk), .r (Fresh[155]), .c ({new_AGEMA_signal_1202, AdderIns_p4[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1143, AdderIns_p3[2]}), .b ({new_AGEMA_signal_1147, AdderIns_p3[6]}), .clk (clk), .r (Fresh[156]), .c ({new_AGEMA_signal_1203, AdderIns_p4[2]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1144, AdderIns_p3[3]}), .b ({new_AGEMA_signal_1148, AdderIns_p3[7]}), .clk (clk), .r (Fresh[157]), .c ({new_AGEMA_signal_1204, AdderIns_p4[3]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1145, AdderIns_p3[4]}), .b ({new_AGEMA_signal_1149, AdderIns_p3[8]}), .clk (clk), .r (Fresh[158]), .c ({new_AGEMA_signal_1205, AdderIns_p4[4]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1146, AdderIns_p3[5]}), .b ({new_AGEMA_signal_1150, AdderIns_p3[9]}), .clk (clk), .r (Fresh[159]), .c ({new_AGEMA_signal_1206, AdderIns_p4[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1147, AdderIns_p3[6]}), .b ({new_AGEMA_signal_1151, AdderIns_p3[10]}), .clk (clk), .r (Fresh[160]), .c ({new_AGEMA_signal_1207, AdderIns_p4[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1148, AdderIns_p3[7]}), .b ({new_AGEMA_signal_1152, AdderIns_p3[11]}), .clk (clk), .r (Fresh[161]), .c ({new_AGEMA_signal_1208, AdderIns_p4[7]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1149, AdderIns_p3[8]}), .b ({new_AGEMA_signal_1153, AdderIns_p3[12]}), .clk (clk), .r (Fresh[162]), .c ({new_AGEMA_signal_1209, AdderIns_p4[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1150, AdderIns_p3[9]}), .b ({new_AGEMA_signal_1154, AdderIns_p3[13]}), .clk (clk), .r (Fresh[163]), .c ({new_AGEMA_signal_1210, AdderIns_p4[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1151, AdderIns_p3[10]}), .b ({new_AGEMA_signal_1155, AdderIns_p3[14]}), .clk (clk), .r (Fresh[164]), .c ({new_AGEMA_signal_1211, AdderIns_p4[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1152, AdderIns_p3[11]}), .b ({new_AGEMA_signal_1156, AdderIns_p3[15]}), .clk (clk), .r (Fresh[165]), .c ({new_AGEMA_signal_1212, AdderIns_p4[11]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1153, AdderIns_p3[12]}), .b ({new_AGEMA_signal_1157, AdderIns_p3[16]}), .clk (clk), .r (Fresh[166]), .c ({new_AGEMA_signal_1213, AdderIns_p4[12]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1154, AdderIns_p3[13]}), .b ({new_AGEMA_signal_1158, AdderIns_p3[17]}), .clk (clk), .r (Fresh[167]), .c ({new_AGEMA_signal_1214, AdderIns_p4[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1155, AdderIns_p3[14]}), .b ({new_AGEMA_signal_1159, AdderIns_p3[18]}), .clk (clk), .r (Fresh[168]), .c ({new_AGEMA_signal_1215, AdderIns_p4[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_15_a2_U1 ( .a ({new_AGEMA_signal_1156, AdderIns_p3[15]}), .b ({new_AGEMA_signal_1160, AdderIns_p3[19]}), .clk (clk), .r (Fresh[169]), .c ({new_AGEMA_signal_1216, AdderIns_p4[15]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_16_a2_U1 ( .a ({new_AGEMA_signal_1157, AdderIns_p3[16]}), .b ({new_AGEMA_signal_1161, AdderIns_p3[20]}), .clk (clk), .r (Fresh[170]), .c ({new_AGEMA_signal_1217, AdderIns_p4[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_17_a2_U1 ( .a ({new_AGEMA_signal_1158, AdderIns_p3[17]}), .b ({new_AGEMA_signal_1162, AdderIns_p3[21]}), .clk (clk), .r (Fresh[171]), .c ({new_AGEMA_signal_1218, AdderIns_p4[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_18_a2_U1 ( .a ({new_AGEMA_signal_1159, AdderIns_p3[18]}), .b ({new_AGEMA_signal_1163, AdderIns_p3[22]}), .clk (clk), .r (Fresh[172]), .c ({new_AGEMA_signal_1219, AdderIns_p4[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_19_a2_U1 ( .a ({new_AGEMA_signal_1160, AdderIns_p3[19]}), .b ({new_AGEMA_signal_1164, AdderIns_p3[23]}), .clk (clk), .r (Fresh[173]), .c ({new_AGEMA_signal_1220, AdderIns_p4[19]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_20_a2_U1 ( .a ({new_AGEMA_signal_1161, AdderIns_p3[20]}), .b ({new_AGEMA_signal_1165, AdderIns_p3[24]}), .clk (clk), .r (Fresh[174]), .c ({new_AGEMA_signal_1221, AdderIns_p4[20]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_21_a2_U1 ( .a ({new_AGEMA_signal_1162, AdderIns_p3[21]}), .b ({new_AGEMA_signal_1166, AdderIns_p3[25]}), .clk (clk), .r (Fresh[175]), .c ({new_AGEMA_signal_1222, AdderIns_p4[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_22_a2_U1 ( .a ({new_AGEMA_signal_1163, AdderIns_p3[22]}), .b ({new_AGEMA_signal_1167, AdderIns_p3[26]}), .clk (clk), .r (Fresh[176]), .c ({new_AGEMA_signal_1223, AdderIns_p4[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_23_a2_U1 ( .a ({new_AGEMA_signal_1164, AdderIns_p3[23]}), .b ({new_AGEMA_signal_1168, AdderIns_p3[27]}), .clk (clk), .r (Fresh[177]), .c ({new_AGEMA_signal_1224, AdderIns_p4[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U29 ( .a ({new_AGEMA_signal_1311, AdderIns_g6[6]}), .b ({new_AGEMA_signal_974, AdderIns_p6[7]}), .c ({new_AGEMA_signal_1373, sum[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U28 ( .a ({new_AGEMA_signal_1279, AdderIns_g6[5]}), .b ({new_AGEMA_signal_971, AdderIns_p6[6]}), .c ({new_AGEMA_signal_1342, sum[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U27 ( .a ({new_AGEMA_signal_1278, AdderIns_g6[4]}), .b ({new_AGEMA_signal_968, AdderIns_p6[5]}), .c ({new_AGEMA_signal_1343, sum[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U26 ( .a ({new_AGEMA_signal_1277, AdderIns_g6[3]}), .b ({new_AGEMA_signal_965, AdderIns_p6[4]}), .c ({new_AGEMA_signal_1344, sum[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_15_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1373, sum[7]}), .a ({new_AGEMA_signal_953, sum[0]}), .c ({new_AGEMA_signal_1406, sum_rotated01[15]}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) U130 ( .a ({1'b0, round_constant[10]}), .b ({new_AGEMA_signal_1405, sum[10]}), .c ({x_round_out_s1[10], x_round_out_s0[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U131 ( .a ({1'b0, round_constant[11]}), .b ({new_AGEMA_signal_1404, sum[11]}), .c ({x_round_out_s1[11], x_round_out_s0[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U132 ( .a ({1'b0, round_constant[12]}), .b ({new_AGEMA_signal_1403, sum[12]}), .c ({x_round_out_s1[12], x_round_out_s0[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U133 ( .a ({1'b0, round_constant[13]}), .b ({new_AGEMA_signal_1402, sum[13]}), .c ({x_round_out_s1[13], x_round_out_s0[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U134 ( .a ({1'b0, round_constant[14]}), .b ({new_AGEMA_signal_1401, sum[14]}), .c ({x_round_out_s1[14], x_round_out_s0[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U135 ( .a ({1'b0, round_constant[15]}), .b ({new_AGEMA_signal_1430, sum[15]}), .c ({x_round_out_s1[15], x_round_out_s0[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U159 ( .a ({1'b0, round_constant[8]}), .b ({new_AGEMA_signal_1400, sum[8]}), .c ({x_round_out_s1[8], x_round_out_s0[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U160 ( .a ({1'b0, round_constant[9]}), .b ({new_AGEMA_signal_1399, sum[9]}), .c ({x_round_out_s1[9], x_round_out_s0[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U168 ( .a ({new_AGEMA_signal_1522, sum_rotated[16]}), .b ({y_round_in_s1[16], y_round_in_s0[16]}), .c ({y_round_out_s1[16], y_round_out_s0[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_0_a1_U1 ( .a ({new_AGEMA_signal_1232, AdderIns_g3[7]}), .b ({new_AGEMA_signal_1281, AdderIns_s4_bc_0_a1_t}), .c ({new_AGEMA_signal_1312, AdderIns_g4[7]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_1228, AdderIns_g3[3]}), .b ({new_AGEMA_signal_1145, AdderIns_p3[4]}), .clk (clk), .r (Fresh[178]), .c ({new_AGEMA_signal_1281, AdderIns_s4_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_1_a1_U1 ( .a ({new_AGEMA_signal_1233, AdderIns_g3[8]}), .b ({new_AGEMA_signal_1282, AdderIns_s4_bc_1_a1_t}), .c ({new_AGEMA_signal_1313, AdderIns_g4[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1229, AdderIns_g3[4]}), .b ({new_AGEMA_signal_1146, AdderIns_p3[5]}), .clk (clk), .r (Fresh[179]), .c ({new_AGEMA_signal_1282, AdderIns_s4_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_2_a1_U1 ( .a ({new_AGEMA_signal_1234, AdderIns_g3[9]}), .b ({new_AGEMA_signal_1283, AdderIns_s4_bc_2_a1_t}), .c ({new_AGEMA_signal_1314, AdderIns_g4[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1230, AdderIns_g3[5]}), .b ({new_AGEMA_signal_1147, AdderIns_p3[6]}), .clk (clk), .r (Fresh[180]), .c ({new_AGEMA_signal_1283, AdderIns_s4_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_3_a1_U1 ( .a ({new_AGEMA_signal_1235, AdderIns_g3[10]}), .b ({new_AGEMA_signal_1284, AdderIns_s4_bc_3_a1_t}), .c ({new_AGEMA_signal_1315, AdderIns_g4[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1231, AdderIns_g3[6]}), .b ({new_AGEMA_signal_1148, AdderIns_p3[7]}), .clk (clk), .r (Fresh[181]), .c ({new_AGEMA_signal_1284, AdderIns_s4_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_4_a1_U1 ( .a ({new_AGEMA_signal_1236, AdderIns_g3[11]}), .b ({new_AGEMA_signal_1285, AdderIns_s4_bc_4_a1_t}), .c ({new_AGEMA_signal_1316, AdderIns_g4[11]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1232, AdderIns_g3[7]}), .b ({new_AGEMA_signal_1149, AdderIns_p3[8]}), .clk (clk), .r (Fresh[182]), .c ({new_AGEMA_signal_1285, AdderIns_s4_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_5_a1_U1 ( .a ({new_AGEMA_signal_1237, AdderIns_g3[12]}), .b ({new_AGEMA_signal_1286, AdderIns_s4_bc_5_a1_t}), .c ({new_AGEMA_signal_1317, AdderIns_g4[12]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1233, AdderIns_g3[8]}), .b ({new_AGEMA_signal_1150, AdderIns_p3[9]}), .clk (clk), .r (Fresh[183]), .c ({new_AGEMA_signal_1286, AdderIns_s4_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_6_a1_U1 ( .a ({new_AGEMA_signal_1238, AdderIns_g3[13]}), .b ({new_AGEMA_signal_1287, AdderIns_s4_bc_6_a1_t}), .c ({new_AGEMA_signal_1318, AdderIns_g4[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1234, AdderIns_g3[9]}), .b ({new_AGEMA_signal_1151, AdderIns_p3[10]}), .clk (clk), .r (Fresh[184]), .c ({new_AGEMA_signal_1287, AdderIns_s4_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_7_a1_U1 ( .a ({new_AGEMA_signal_1239, AdderIns_g3[14]}), .b ({new_AGEMA_signal_1288, AdderIns_s4_bc_7_a1_t}), .c ({new_AGEMA_signal_1319, AdderIns_g4[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1235, AdderIns_g3[10]}), .b ({new_AGEMA_signal_1152, AdderIns_p3[11]}), .clk (clk), .r (Fresh[185]), .c ({new_AGEMA_signal_1288, AdderIns_s4_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_8_a1_U1 ( .a ({new_AGEMA_signal_1240, AdderIns_g3[15]}), .b ({new_AGEMA_signal_1289, AdderIns_s4_bc_8_a1_t}), .c ({new_AGEMA_signal_1320, AdderIns_g4[15]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1236, AdderIns_g3[11]}), .b ({new_AGEMA_signal_1153, AdderIns_p3[12]}), .clk (clk), .r (Fresh[186]), .c ({new_AGEMA_signal_1289, AdderIns_s4_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_9_a1_U1 ( .a ({new_AGEMA_signal_1241, AdderIns_g3[16]}), .b ({new_AGEMA_signal_1290, AdderIns_s4_bc_9_a1_t}), .c ({new_AGEMA_signal_1321, AdderIns_g4[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1237, AdderIns_g3[12]}), .b ({new_AGEMA_signal_1154, AdderIns_p3[13]}), .clk (clk), .r (Fresh[187]), .c ({new_AGEMA_signal_1290, AdderIns_s4_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_10_a1_U1 ( .a ({new_AGEMA_signal_1242, AdderIns_g3[17]}), .b ({new_AGEMA_signal_1291, AdderIns_s4_bc_10_a1_t}), .c ({new_AGEMA_signal_1322, AdderIns_g4[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1238, AdderIns_g3[13]}), .b ({new_AGEMA_signal_1155, AdderIns_p3[14]}), .clk (clk), .r (Fresh[188]), .c ({new_AGEMA_signal_1291, AdderIns_s4_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_11_a1_U1 ( .a ({new_AGEMA_signal_1243, AdderIns_g3[18]}), .b ({new_AGEMA_signal_1292, AdderIns_s4_bc_11_a1_t}), .c ({new_AGEMA_signal_1323, AdderIns_g4[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1239, AdderIns_g3[14]}), .b ({new_AGEMA_signal_1156, AdderIns_p3[15]}), .clk (clk), .r (Fresh[189]), .c ({new_AGEMA_signal_1292, AdderIns_s4_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_12_a1_U1 ( .a ({new_AGEMA_signal_1244, AdderIns_g3[19]}), .b ({new_AGEMA_signal_1293, AdderIns_s4_bc_12_a1_t}), .c ({new_AGEMA_signal_1324, AdderIns_g4[19]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1240, AdderIns_g3[15]}), .b ({new_AGEMA_signal_1157, AdderIns_p3[16]}), .clk (clk), .r (Fresh[190]), .c ({new_AGEMA_signal_1293, AdderIns_s4_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_13_a1_U1 ( .a ({new_AGEMA_signal_1245, AdderIns_g3[20]}), .b ({new_AGEMA_signal_1294, AdderIns_s4_bc_13_a1_t}), .c ({new_AGEMA_signal_1325, AdderIns_g4[20]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1241, AdderIns_g3[16]}), .b ({new_AGEMA_signal_1158, AdderIns_p3[17]}), .clk (clk), .r (Fresh[191]), .c ({new_AGEMA_signal_1294, AdderIns_s4_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_14_a1_U1 ( .a ({new_AGEMA_signal_1246, AdderIns_g3[21]}), .b ({new_AGEMA_signal_1295, AdderIns_s4_bc_14_a1_t}), .c ({new_AGEMA_signal_1326, AdderIns_g4[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1242, AdderIns_g3[17]}), .b ({new_AGEMA_signal_1159, AdderIns_p3[18]}), .clk (clk), .r (Fresh[192]), .c ({new_AGEMA_signal_1295, AdderIns_s4_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_15_a1_U1 ( .a ({new_AGEMA_signal_1247, AdderIns_g3[22]}), .b ({new_AGEMA_signal_1296, AdderIns_s4_bc_15_a1_t}), .c ({new_AGEMA_signal_1327, AdderIns_g4[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1243, AdderIns_g3[18]}), .b ({new_AGEMA_signal_1160, AdderIns_p3[19]}), .clk (clk), .r (Fresh[193]), .c ({new_AGEMA_signal_1296, AdderIns_s4_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_16_a1_U1 ( .a ({new_AGEMA_signal_1248, AdderIns_g3[23]}), .b ({new_AGEMA_signal_1297, AdderIns_s4_bc_16_a1_t}), .c ({new_AGEMA_signal_1328, AdderIns_g4[23]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_16_a1_a1_U1 ( .a ({new_AGEMA_signal_1244, AdderIns_g3[19]}), .b ({new_AGEMA_signal_1161, AdderIns_p3[20]}), .clk (clk), .r (Fresh[194]), .c ({new_AGEMA_signal_1297, AdderIns_s4_bc_16_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_17_a1_U1 ( .a ({new_AGEMA_signal_1249, AdderIns_g3[24]}), .b ({new_AGEMA_signal_1298, AdderIns_s4_bc_17_a1_t}), .c ({new_AGEMA_signal_1329, AdderIns_g4[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_17_a1_a1_U1 ( .a ({new_AGEMA_signal_1245, AdderIns_g3[20]}), .b ({new_AGEMA_signal_1162, AdderIns_p3[21]}), .clk (clk), .r (Fresh[195]), .c ({new_AGEMA_signal_1298, AdderIns_s4_bc_17_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_18_a1_U1 ( .a ({new_AGEMA_signal_1250, AdderIns_g3[25]}), .b ({new_AGEMA_signal_1299, AdderIns_s4_bc_18_a1_t}), .c ({new_AGEMA_signal_1330, AdderIns_g4[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_18_a1_a1_U1 ( .a ({new_AGEMA_signal_1246, AdderIns_g3[21]}), .b ({new_AGEMA_signal_1163, AdderIns_p3[22]}), .clk (clk), .r (Fresh[196]), .c ({new_AGEMA_signal_1299, AdderIns_s4_bc_18_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_19_a1_U1 ( .a ({new_AGEMA_signal_1251, AdderIns_g3[26]}), .b ({new_AGEMA_signal_1300, AdderIns_s4_bc_19_a1_t}), .c ({new_AGEMA_signal_1331, AdderIns_g4[26]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_19_a1_a1_U1 ( .a ({new_AGEMA_signal_1247, AdderIns_g3[22]}), .b ({new_AGEMA_signal_1164, AdderIns_p3[23]}), .clk (clk), .r (Fresh[197]), .c ({new_AGEMA_signal_1300, AdderIns_s4_bc_19_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_20_a1_U1 ( .a ({new_AGEMA_signal_1252, AdderIns_g3[27]}), .b ({new_AGEMA_signal_1301, AdderIns_s4_bc_20_a1_t}), .c ({new_AGEMA_signal_1332, AdderIns_g4[27]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_20_a1_a1_U1 ( .a ({new_AGEMA_signal_1248, AdderIns_g3[23]}), .b ({new_AGEMA_signal_1165, AdderIns_p3[24]}), .clk (clk), .r (Fresh[198]), .c ({new_AGEMA_signal_1301, AdderIns_s4_bc_20_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_21_a1_U1 ( .a ({new_AGEMA_signal_1253, AdderIns_g3[28]}), .b ({new_AGEMA_signal_1302, AdderIns_s4_bc_21_a1_t}), .c ({new_AGEMA_signal_1333, AdderIns_g4[28]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_21_a1_a1_U1 ( .a ({new_AGEMA_signal_1249, AdderIns_g3[24]}), .b ({new_AGEMA_signal_1166, AdderIns_p3[25]}), .clk (clk), .r (Fresh[199]), .c ({new_AGEMA_signal_1302, AdderIns_s4_bc_21_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_22_a1_U1 ( .a ({new_AGEMA_signal_1254, AdderIns_g3[29]}), .b ({new_AGEMA_signal_1303, AdderIns_s4_bc_22_a1_t}), .c ({new_AGEMA_signal_1334, AdderIns_g4[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_22_a1_a1_U1 ( .a ({new_AGEMA_signal_1250, AdderIns_g3[25]}), .b ({new_AGEMA_signal_1167, AdderIns_p3[26]}), .clk (clk), .r (Fresh[200]), .c ({new_AGEMA_signal_1303, AdderIns_s4_bc_22_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_23_a1_U1 ( .a ({new_AGEMA_signal_1255, AdderIns_g3[30]}), .b ({new_AGEMA_signal_1304, AdderIns_s4_bc_23_a1_t}), .c ({new_AGEMA_signal_1335, AdderIns_g4[30]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s4_bc_23_a1_a1_U1 ( .a ({new_AGEMA_signal_1251, AdderIns_g3[26]}), .b ({new_AGEMA_signal_1168, AdderIns_p3[27]}), .clk (clk), .r (Fresh[201]), .c ({new_AGEMA_signal_1304, AdderIns_s4_bc_23_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_0_a1_U1 ( .a ({new_AGEMA_signal_1312, AdderIns_g4[7]}), .b ({new_AGEMA_signal_1257, AdderIns_s5_gc_0_a1_t}), .c ({new_AGEMA_signal_1348, AdderIns_g6[7]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1201, AdderIns_p4[0]}), .clk (clk), .r (Fresh[202]), .c ({new_AGEMA_signal_1257, AdderIns_s5_gc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_1_a1_U1 ( .a ({new_AGEMA_signal_1313, AdderIns_g4[8]}), .b ({new_AGEMA_signal_1258, AdderIns_s5_gc_1_a1_t}), .c ({new_AGEMA_signal_1349, AdderIns_g6[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1109, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1202, AdderIns_p4[1]}), .clk (clk), .r (Fresh[203]), .c ({new_AGEMA_signal_1258, AdderIns_s5_gc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_2_a1_U1 ( .a ({new_AGEMA_signal_1314, AdderIns_g4[9]}), .b ({new_AGEMA_signal_1259, AdderIns_s5_gc_2_a1_t}), .c ({new_AGEMA_signal_1350, AdderIns_g6[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1169, AdderIns_g6[1]}), .b ({new_AGEMA_signal_1203, AdderIns_p4[2]}), .clk (clk), .r (Fresh[204]), .c ({new_AGEMA_signal_1259, AdderIns_s5_gc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_3_a1_U1 ( .a ({new_AGEMA_signal_1315, AdderIns_g4[10]}), .b ({new_AGEMA_signal_1305, AdderIns_s5_gc_3_a1_t}), .c ({new_AGEMA_signal_1351, AdderIns_g6[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1227, AdderIns_g6[2]}), .b ({new_AGEMA_signal_1204, AdderIns_p4[3]}), .clk (clk), .r (Fresh[205]), .c ({new_AGEMA_signal_1305, AdderIns_s5_gc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_4_a1_U1 ( .a ({new_AGEMA_signal_1316, AdderIns_g4[11]}), .b ({new_AGEMA_signal_1336, AdderIns_s5_gc_4_a1_t}), .c ({new_AGEMA_signal_1352, AdderIns_g6[11]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1277, AdderIns_g6[3]}), .b ({new_AGEMA_signal_1205, AdderIns_p4[4]}), .clk (clk), .r (Fresh[206]), .c ({new_AGEMA_signal_1336, AdderIns_s5_gc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_5_a1_U1 ( .a ({new_AGEMA_signal_1317, AdderIns_g4[12]}), .b ({new_AGEMA_signal_1337, AdderIns_s5_gc_5_a1_t}), .c ({new_AGEMA_signal_1353, AdderIns_g6[12]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1278, AdderIns_g6[4]}), .b ({new_AGEMA_signal_1206, AdderIns_p4[5]}), .clk (clk), .r (Fresh[207]), .c ({new_AGEMA_signal_1337, AdderIns_s5_gc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_6_a1_U1 ( .a ({new_AGEMA_signal_1318, AdderIns_g4[13]}), .b ({new_AGEMA_signal_1338, AdderIns_s5_gc_6_a1_t}), .c ({new_AGEMA_signal_1354, AdderIns_g6[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1279, AdderIns_g6[5]}), .b ({new_AGEMA_signal_1207, AdderIns_p4[6]}), .clk (clk), .r (Fresh[208]), .c ({new_AGEMA_signal_1338, AdderIns_s5_gc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_7_a1_U1 ( .a ({new_AGEMA_signal_1319, AdderIns_g4[14]}), .b ({new_AGEMA_signal_1355, AdderIns_s5_gc_7_a1_t}), .c ({new_AGEMA_signal_1375, AdderIns_g6[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_gc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1311, AdderIns_g6[6]}), .b ({new_AGEMA_signal_1208, AdderIns_p4[7]}), .clk (clk), .r (Fresh[209]), .c ({new_AGEMA_signal_1355, AdderIns_s5_gc_7_a1_t}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1202, AdderIns_p4[1]}), .b ({new_AGEMA_signal_1210, AdderIns_p4[9]}), .clk (clk), .r (Fresh[210]), .c ({new_AGEMA_signal_1260, AdderIns_p5[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1203, AdderIns_p4[2]}), .b ({new_AGEMA_signal_1211, AdderIns_p4[10]}), .clk (clk), .r (Fresh[211]), .c ({new_AGEMA_signal_1261, AdderIns_p5[2]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1204, AdderIns_p4[3]}), .b ({new_AGEMA_signal_1212, AdderIns_p4[11]}), .clk (clk), .r (Fresh[212]), .c ({new_AGEMA_signal_1262, AdderIns_p5[3]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1205, AdderIns_p4[4]}), .b ({new_AGEMA_signal_1213, AdderIns_p4[12]}), .clk (clk), .r (Fresh[213]), .c ({new_AGEMA_signal_1263, AdderIns_p5[4]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1206, AdderIns_p4[5]}), .b ({new_AGEMA_signal_1214, AdderIns_p4[13]}), .clk (clk), .r (Fresh[214]), .c ({new_AGEMA_signal_1264, AdderIns_p5[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1207, AdderIns_p4[6]}), .b ({new_AGEMA_signal_1215, AdderIns_p4[14]}), .clk (clk), .r (Fresh[215]), .c ({new_AGEMA_signal_1265, AdderIns_p5[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1208, AdderIns_p4[7]}), .b ({new_AGEMA_signal_1216, AdderIns_p4[15]}), .clk (clk), .r (Fresh[216]), .c ({new_AGEMA_signal_1266, AdderIns_p5[7]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1209, AdderIns_p4[8]}), .b ({new_AGEMA_signal_1217, AdderIns_p4[16]}), .clk (clk), .r (Fresh[217]), .c ({new_AGEMA_signal_1267, AdderIns_p5[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1210, AdderIns_p4[9]}), .b ({new_AGEMA_signal_1218, AdderIns_p4[17]}), .clk (clk), .r (Fresh[218]), .c ({new_AGEMA_signal_1268, AdderIns_p5[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1211, AdderIns_p4[10]}), .b ({new_AGEMA_signal_1219, AdderIns_p4[18]}), .clk (clk), .r (Fresh[219]), .c ({new_AGEMA_signal_1269, AdderIns_p5[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1212, AdderIns_p4[11]}), .b ({new_AGEMA_signal_1220, AdderIns_p4[19]}), .clk (clk), .r (Fresh[220]), .c ({new_AGEMA_signal_1270, AdderIns_p5[11]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1213, AdderIns_p4[12]}), .b ({new_AGEMA_signal_1221, AdderIns_p4[20]}), .clk (clk), .r (Fresh[221]), .c ({new_AGEMA_signal_1271, AdderIns_p5[12]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1214, AdderIns_p4[13]}), .b ({new_AGEMA_signal_1222, AdderIns_p4[21]}), .clk (clk), .r (Fresh[222]), .c ({new_AGEMA_signal_1272, AdderIns_p5[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1215, AdderIns_p4[14]}), .b ({new_AGEMA_signal_1223, AdderIns_p4[22]}), .clk (clk), .r (Fresh[223]), .c ({new_AGEMA_signal_1273, AdderIns_p5[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_15_a2_U1 ( .a ({new_AGEMA_signal_1216, AdderIns_p4[15]}), .b ({new_AGEMA_signal_1224, AdderIns_p4[23]}), .clk (clk), .r (Fresh[224]), .c ({new_AGEMA_signal_1274, AdderIns_p5[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U31 ( .a ({new_AGEMA_signal_1349, AdderIns_g6[8]}), .b ({new_AGEMA_signal_980, AdderIns_p6[9]}), .c ({new_AGEMA_signal_1399, sum[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U30 ( .a ({new_AGEMA_signal_1348, AdderIns_g6[7]}), .b ({new_AGEMA_signal_977, AdderIns_p6[8]}), .c ({new_AGEMA_signal_1400, sum[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U6 ( .a ({new_AGEMA_signal_1375, AdderIns_g6[14]}), .b ({new_AGEMA_signal_998, AdderIns_p6[15]}), .c ({new_AGEMA_signal_1430, sum[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U5 ( .a ({new_AGEMA_signal_1354, AdderIns_g6[13]}), .b ({new_AGEMA_signal_995, AdderIns_p6[14]}), .c ({new_AGEMA_signal_1401, sum[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U4 ( .a ({new_AGEMA_signal_1353, AdderIns_g6[12]}), .b ({new_AGEMA_signal_992, AdderIns_p6[13]}), .c ({new_AGEMA_signal_1402, sum[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U3 ( .a ({new_AGEMA_signal_1352, AdderIns_g6[11]}), .b ({new_AGEMA_signal_989, AdderIns_p6[12]}), .c ({new_AGEMA_signal_1403, sum[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U2 ( .a ({new_AGEMA_signal_1351, AdderIns_g6[10]}), .b ({new_AGEMA_signal_986, AdderIns_p6[11]}), .c ({new_AGEMA_signal_1404, sum[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U1 ( .a ({new_AGEMA_signal_1350, AdderIns_g6[9]}), .b ({new_AGEMA_signal_983, AdderIns_p6[10]}), .c ({new_AGEMA_signal_1405, sum[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_16_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1400, sum[8]}), .a ({new_AGEMA_signal_1225, sum[1]}), .c ({new_AGEMA_signal_1431, sum_rotated01[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_17_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1399, sum[9]}), .a ({new_AGEMA_signal_1275, sum[2]}), .c ({new_AGEMA_signal_1432, sum_rotated01[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_18_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1405, sum[10]}), .a ({new_AGEMA_signal_1309, sum[3]}), .c ({new_AGEMA_signal_1433, sum_rotated01[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_19_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1404, sum[11]}), .a ({new_AGEMA_signal_1344, sum[4]}), .c ({new_AGEMA_signal_1434, sum_rotated01[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_20_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1403, sum[12]}), .a ({new_AGEMA_signal_1343, sum[5]}), .c ({new_AGEMA_signal_1435, sum_rotated01[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_21_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1402, sum[13]}), .a ({new_AGEMA_signal_1342, sum[6]}), .c ({new_AGEMA_signal_1436, sum_rotated01[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_22_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1401, sum[14]}), .a ({new_AGEMA_signal_1373, sum[7]}), .c ({new_AGEMA_signal_1437, sum_rotated01[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_23_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1430, sum[15]}), .a ({new_AGEMA_signal_1400, sum[8]}), .c ({new_AGEMA_signal_1455, sum_rotated01[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_16_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1430, sum[15]}), .a ({new_AGEMA_signal_953, sum[0]}), .c ({new_AGEMA_signal_1457, sum_rotated23[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_16_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1431, sum_rotated01[16]}), .a ({new_AGEMA_signal_1457, sum_rotated23[16]}), .c ({new_AGEMA_signal_1522, sum_rotated[16]}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) U136 ( .a ({1'b0, round_constant[16]}), .b ({new_AGEMA_signal_1429, sum[16]}), .c ({x_round_out_s1[16], x_round_out_s0[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U137 ( .a ({1'b0, round_constant[17]}), .b ({new_AGEMA_signal_1454, sum[17]}), .c ({x_round_out_s1[17], x_round_out_s0[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U138 ( .a ({1'b0, round_constant[18]}), .b ({new_AGEMA_signal_1453, sum[18]}), .c ({x_round_out_s1[18], x_round_out_s0[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U139 ( .a ({1'b0, round_constant[19]}), .b ({new_AGEMA_signal_1452, sum[19]}), .c ({x_round_out_s1[19], x_round_out_s0[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U141 ( .a ({1'b0, round_constant[20]}), .b ({new_AGEMA_signal_1451, sum[20]}), .c ({x_round_out_s1[20], x_round_out_s0[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U142 ( .a ({1'b0, round_constant[21]}), .b ({new_AGEMA_signal_1450, sum[21]}), .c ({x_round_out_s1[21], x_round_out_s0[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U143 ( .a ({1'b0, round_constant[22]}), .b ({new_AGEMA_signal_1449, sum[22]}), .c ({x_round_out_s1[22], x_round_out_s0[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U144 ( .a ({1'b0, round_constant[23]}), .b ({new_AGEMA_signal_1448, sum[23]}), .c ({x_round_out_s1[23], x_round_out_s0[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U145 ( .a ({1'b0, round_constant[24]}), .b ({new_AGEMA_signal_1447, sum[24]}), .c ({x_round_out_s1[24], x_round_out_s0[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U146 ( .a ({1'b0, round_constant[25]}), .b ({new_AGEMA_signal_1446, sum[25]}), .c ({x_round_out_s1[25], x_round_out_s0[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U147 ( .a ({1'b0, round_constant[26]}), .b ({new_AGEMA_signal_1445, sum[26]}), .c ({x_round_out_s1[26], x_round_out_s0[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U148 ( .a ({1'b0, round_constant[27]}), .b ({new_AGEMA_signal_1444, sum[27]}), .c ({x_round_out_s1[27], x_round_out_s0[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U149 ( .a ({1'b0, round_constant[28]}), .b ({new_AGEMA_signal_1443, sum[28]}), .c ({x_round_out_s1[28], x_round_out_s0[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U150 ( .a ({1'b0, round_constant[29]}), .b ({new_AGEMA_signal_1442, sum[29]}), .c ({x_round_out_s1[29], x_round_out_s0[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U152 ( .a ({1'b0, round_constant[30]}), .b ({new_AGEMA_signal_1441, sum[30]}), .c ({x_round_out_s1[30], x_round_out_s0[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U153 ( .a ({1'b0, round_constant[31]}), .b ({new_AGEMA_signal_1473, sum[31]}), .c ({x_round_out_s1[31], x_round_out_s0[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U161 ( .a ({new_AGEMA_signal_1583, sum_rotated[0]}), .b ({y_round_in_s1[0], y_round_in_s0[0]}), .c ({y_round_out_s1[0], y_round_out_s0[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U162 ( .a ({new_AGEMA_signal_1539, sum_rotated[10]}), .b ({y_round_in_s1[10], y_round_in_s0[10]}), .c ({y_round_out_s1[10], y_round_out_s0[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U163 ( .a ({new_AGEMA_signal_1540, sum_rotated[11]}), .b ({y_round_in_s1[11], y_round_in_s0[11]}), .c ({y_round_out_s1[11], y_round_out_s0[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U164 ( .a ({new_AGEMA_signal_1541, sum_rotated[12]}), .b ({y_round_in_s1[12], y_round_in_s0[12]}), .c ({y_round_out_s1[12], y_round_out_s0[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U165 ( .a ({new_AGEMA_signal_1542, sum_rotated[13]}), .b ({y_round_in_s1[13], y_round_in_s0[13]}), .c ({y_round_out_s1[13], y_round_out_s0[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U166 ( .a ({new_AGEMA_signal_1585, sum_rotated[14]}), .b ({y_round_in_s1[14], y_round_in_s0[14]}), .c ({y_round_out_s1[14], y_round_out_s0[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U167 ( .a ({new_AGEMA_signal_1586, sum_rotated[15]}), .b ({y_round_in_s1[15], y_round_in_s0[15]}), .c ({y_round_out_s1[15], y_round_out_s0[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U169 ( .a ({new_AGEMA_signal_1523, sum_rotated[17]}), .b ({y_round_in_s1[17], y_round_in_s0[17]}), .c ({y_round_out_s1[17], y_round_out_s0[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U170 ( .a ({new_AGEMA_signal_1543, sum_rotated[18]}), .b ({y_round_in_s1[18], y_round_in_s0[18]}), .c ({y_round_out_s1[18], y_round_out_s0[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U171 ( .a ({new_AGEMA_signal_1544, sum_rotated[19]}), .b ({y_round_in_s1[19], y_round_in_s0[19]}), .c ({y_round_out_s1[19], y_round_out_s0[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U172 ( .a ({new_AGEMA_signal_1531, sum_rotated[1]}), .b ({y_round_in_s1[1], y_round_in_s0[1]}), .c ({y_round_out_s1[1], y_round_out_s0[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U173 ( .a ({new_AGEMA_signal_1545, sum_rotated[20]}), .b ({y_round_in_s1[20], y_round_in_s0[20]}), .c ({y_round_out_s1[20], y_round_out_s0[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U174 ( .a ({new_AGEMA_signal_1546, sum_rotated[21]}), .b ({y_round_in_s1[21], y_round_in_s0[21]}), .c ({y_round_out_s1[21], y_round_out_s0[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U175 ( .a ({new_AGEMA_signal_1547, sum_rotated[22]}), .b ({y_round_in_s1[22], y_round_in_s0[22]}), .c ({y_round_out_s1[22], y_round_out_s0[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U176 ( .a ({new_AGEMA_signal_1548, sum_rotated[23]}), .b ({y_round_in_s1[23], y_round_in_s0[23]}), .c ({y_round_out_s1[23], y_round_out_s0[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U177 ( .a ({new_AGEMA_signal_1549, sum_rotated[24]}), .b ({y_round_in_s1[24], y_round_in_s0[24]}), .c ({y_round_out_s1[24], y_round_out_s0[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U178 ( .a ({new_AGEMA_signal_1550, sum_rotated[25]}), .b ({y_round_in_s1[25], y_round_in_s0[25]}), .c ({y_round_out_s1[25], y_round_out_s0[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U179 ( .a ({new_AGEMA_signal_1551, sum_rotated[26]}), .b ({y_round_in_s1[26], y_round_in_s0[26]}), .c ({y_round_out_s1[26], y_round_out_s0[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U180 ( .a ({new_AGEMA_signal_1552, sum_rotated[27]}), .b ({y_round_in_s1[27], y_round_in_s0[27]}), .c ({y_round_out_s1[27], y_round_out_s0[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U181 ( .a ({new_AGEMA_signal_1553, sum_rotated[28]}), .b ({y_round_in_s1[28], y_round_in_s0[28]}), .c ({y_round_out_s1[28], y_round_out_s0[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U182 ( .a ({new_AGEMA_signal_1554, sum_rotated[29]}), .b ({y_round_in_s1[29], y_round_in_s0[29]}), .c ({y_round_out_s1[29], y_round_out_s0[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U183 ( .a ({new_AGEMA_signal_1532, sum_rotated[2]}), .b ({y_round_in_s1[2], y_round_in_s0[2]}), .c ({y_round_out_s1[2], y_round_out_s0[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U184 ( .a ({new_AGEMA_signal_1555, sum_rotated[30]}), .b ({y_round_in_s1[30], y_round_in_s0[30]}), .c ({y_round_out_s1[30], y_round_out_s0[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U185 ( .a ({new_AGEMA_signal_1556, sum_rotated[31]}), .b ({y_round_in_s1[31], y_round_in_s0[31]}), .c ({y_round_out_s1[31], y_round_out_s0[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U186 ( .a ({new_AGEMA_signal_1533, sum_rotated[3]}), .b ({y_round_in_s1[3], y_round_in_s0[3]}), .c ({y_round_out_s1[3], y_round_out_s0[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U187 ( .a ({new_AGEMA_signal_1534, sum_rotated[4]}), .b ({y_round_in_s1[4], y_round_in_s0[4]}), .c ({y_round_out_s1[4], y_round_out_s0[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U188 ( .a ({new_AGEMA_signal_1535, sum_rotated[5]}), .b ({y_round_in_s1[5], y_round_in_s0[5]}), .c ({y_round_out_s1[5], y_round_out_s0[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U189 ( .a ({new_AGEMA_signal_1536, sum_rotated[6]}), .b ({y_round_in_s1[6], y_round_in_s0[6]}), .c ({y_round_out_s1[6], y_round_out_s0[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U190 ( .a ({new_AGEMA_signal_1584, sum_rotated[7]}), .b ({y_round_in_s1[7], y_round_in_s0[7]}), .c ({y_round_out_s1[7], y_round_out_s0[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U191 ( .a ({new_AGEMA_signal_1537, sum_rotated[8]}), .b ({y_round_in_s1[8], y_round_in_s0[8]}), .c ({y_round_out_s1[8], y_round_out_s0[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U192 ( .a ({new_AGEMA_signal_1538, sum_rotated[9]}), .b ({y_round_in_s1[9], y_round_in_s0[9]}), .c ({y_round_out_s1[9], y_round_out_s0[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_0_a1_U1 ( .a ({new_AGEMA_signal_1320, AdderIns_g4[15]}), .b ({new_AGEMA_signal_1356, AdderIns_s5_bc_0_a1_t}), .c ({new_AGEMA_signal_1376, AdderIns_g6[15]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_1312, AdderIns_g4[7]}), .b ({new_AGEMA_signal_1209, AdderIns_p4[8]}), .clk (clk), .r (Fresh[225]), .c ({new_AGEMA_signal_1356, AdderIns_s5_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_1_a1_U1 ( .a ({new_AGEMA_signal_1321, AdderIns_g4[16]}), .b ({new_AGEMA_signal_1357, AdderIns_s5_bc_1_a1_t}), .c ({new_AGEMA_signal_1377, AdderIns_g5[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1313, AdderIns_g4[8]}), .b ({new_AGEMA_signal_1210, AdderIns_p4[9]}), .clk (clk), .r (Fresh[226]), .c ({new_AGEMA_signal_1357, AdderIns_s5_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_2_a1_U1 ( .a ({new_AGEMA_signal_1322, AdderIns_g4[17]}), .b ({new_AGEMA_signal_1358, AdderIns_s5_bc_2_a1_t}), .c ({new_AGEMA_signal_1378, AdderIns_g5[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1314, AdderIns_g4[9]}), .b ({new_AGEMA_signal_1211, AdderIns_p4[10]}), .clk (clk), .r (Fresh[227]), .c ({new_AGEMA_signal_1358, AdderIns_s5_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_3_a1_U1 ( .a ({new_AGEMA_signal_1323, AdderIns_g4[18]}), .b ({new_AGEMA_signal_1359, AdderIns_s5_bc_3_a1_t}), .c ({new_AGEMA_signal_1379, AdderIns_g5[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1315, AdderIns_g4[10]}), .b ({new_AGEMA_signal_1212, AdderIns_p4[11]}), .clk (clk), .r (Fresh[228]), .c ({new_AGEMA_signal_1359, AdderIns_s5_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_4_a1_U1 ( .a ({new_AGEMA_signal_1324, AdderIns_g4[19]}), .b ({new_AGEMA_signal_1360, AdderIns_s5_bc_4_a1_t}), .c ({new_AGEMA_signal_1380, AdderIns_g5[19]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1316, AdderIns_g4[11]}), .b ({new_AGEMA_signal_1213, AdderIns_p4[12]}), .clk (clk), .r (Fresh[229]), .c ({new_AGEMA_signal_1360, AdderIns_s5_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_5_a1_U1 ( .a ({new_AGEMA_signal_1325, AdderIns_g4[20]}), .b ({new_AGEMA_signal_1361, AdderIns_s5_bc_5_a1_t}), .c ({new_AGEMA_signal_1381, AdderIns_g5[20]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1317, AdderIns_g4[12]}), .b ({new_AGEMA_signal_1214, AdderIns_p4[13]}), .clk (clk), .r (Fresh[230]), .c ({new_AGEMA_signal_1361, AdderIns_s5_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_6_a1_U1 ( .a ({new_AGEMA_signal_1326, AdderIns_g4[21]}), .b ({new_AGEMA_signal_1362, AdderIns_s5_bc_6_a1_t}), .c ({new_AGEMA_signal_1382, AdderIns_g5[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1318, AdderIns_g4[13]}), .b ({new_AGEMA_signal_1215, AdderIns_p4[14]}), .clk (clk), .r (Fresh[231]), .c ({new_AGEMA_signal_1362, AdderIns_s5_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_7_a1_U1 ( .a ({new_AGEMA_signal_1327, AdderIns_g4[22]}), .b ({new_AGEMA_signal_1363, AdderIns_s5_bc_7_a1_t}), .c ({new_AGEMA_signal_1383, AdderIns_g5[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1319, AdderIns_g4[14]}), .b ({new_AGEMA_signal_1216, AdderIns_p4[15]}), .clk (clk), .r (Fresh[232]), .c ({new_AGEMA_signal_1363, AdderIns_s5_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_8_a1_U1 ( .a ({new_AGEMA_signal_1328, AdderIns_g4[23]}), .b ({new_AGEMA_signal_1364, AdderIns_s5_bc_8_a1_t}), .c ({new_AGEMA_signal_1384, AdderIns_g5[23]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1320, AdderIns_g4[15]}), .b ({new_AGEMA_signal_1217, AdderIns_p4[16]}), .clk (clk), .r (Fresh[233]), .c ({new_AGEMA_signal_1364, AdderIns_s5_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_9_a1_U1 ( .a ({new_AGEMA_signal_1329, AdderIns_g4[24]}), .b ({new_AGEMA_signal_1365, AdderIns_s5_bc_9_a1_t}), .c ({new_AGEMA_signal_1385, AdderIns_g5[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1321, AdderIns_g4[16]}), .b ({new_AGEMA_signal_1218, AdderIns_p4[17]}), .clk (clk), .r (Fresh[234]), .c ({new_AGEMA_signal_1365, AdderIns_s5_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_10_a1_U1 ( .a ({new_AGEMA_signal_1330, AdderIns_g4[25]}), .b ({new_AGEMA_signal_1366, AdderIns_s5_bc_10_a1_t}), .c ({new_AGEMA_signal_1386, AdderIns_g5[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1322, AdderIns_g4[17]}), .b ({new_AGEMA_signal_1219, AdderIns_p4[18]}), .clk (clk), .r (Fresh[235]), .c ({new_AGEMA_signal_1366, AdderIns_s5_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_11_a1_U1 ( .a ({new_AGEMA_signal_1331, AdderIns_g4[26]}), .b ({new_AGEMA_signal_1367, AdderIns_s5_bc_11_a1_t}), .c ({new_AGEMA_signal_1387, AdderIns_g5[26]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1323, AdderIns_g4[18]}), .b ({new_AGEMA_signal_1220, AdderIns_p4[19]}), .clk (clk), .r (Fresh[236]), .c ({new_AGEMA_signal_1367, AdderIns_s5_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_12_a1_U1 ( .a ({new_AGEMA_signal_1332, AdderIns_g4[27]}), .b ({new_AGEMA_signal_1368, AdderIns_s5_bc_12_a1_t}), .c ({new_AGEMA_signal_1388, AdderIns_g5[27]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1324, AdderIns_g4[19]}), .b ({new_AGEMA_signal_1221, AdderIns_p4[20]}), .clk (clk), .r (Fresh[237]), .c ({new_AGEMA_signal_1368, AdderIns_s5_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_13_a1_U1 ( .a ({new_AGEMA_signal_1333, AdderIns_g4[28]}), .b ({new_AGEMA_signal_1369, AdderIns_s5_bc_13_a1_t}), .c ({new_AGEMA_signal_1389, AdderIns_g5[28]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1325, AdderIns_g4[20]}), .b ({new_AGEMA_signal_1222, AdderIns_p4[21]}), .clk (clk), .r (Fresh[238]), .c ({new_AGEMA_signal_1369, AdderIns_s5_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_14_a1_U1 ( .a ({new_AGEMA_signal_1334, AdderIns_g4[29]}), .b ({new_AGEMA_signal_1370, AdderIns_s5_bc_14_a1_t}), .c ({new_AGEMA_signal_1390, AdderIns_g5[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1326, AdderIns_g4[21]}), .b ({new_AGEMA_signal_1223, AdderIns_p4[22]}), .clk (clk), .r (Fresh[239]), .c ({new_AGEMA_signal_1370, AdderIns_s5_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_15_a1_U1 ( .a ({new_AGEMA_signal_1335, AdderIns_g4[30]}), .b ({new_AGEMA_signal_1371, AdderIns_s5_bc_15_a1_t}), .c ({new_AGEMA_signal_1391, AdderIns_g5[30]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s5_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1327, AdderIns_g4[22]}), .b ({new_AGEMA_signal_1224, AdderIns_p4[23]}), .clk (clk), .r (Fresh[240]), .c ({new_AGEMA_signal_1371, AdderIns_s5_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_1_a1_U1 ( .a ({new_AGEMA_signal_1377, AdderIns_g5[16]}), .b ({new_AGEMA_signal_1306, AdderIns_s6_gc_1_a1_t}), .c ({new_AGEMA_signal_1414, AdderIns_g6[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1109, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1260, AdderIns_p5[1]}), .clk (clk), .r (Fresh[241]), .c ({new_AGEMA_signal_1306, AdderIns_s6_gc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_2_a1_U1 ( .a ({new_AGEMA_signal_1378, AdderIns_g5[17]}), .b ({new_AGEMA_signal_1307, AdderIns_s6_gc_2_a1_t}), .c ({new_AGEMA_signal_1415, AdderIns_g6[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1169, AdderIns_g6[1]}), .b ({new_AGEMA_signal_1261, AdderIns_p5[2]}), .clk (clk), .r (Fresh[242]), .c ({new_AGEMA_signal_1307, AdderIns_s6_gc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_3_a1_U1 ( .a ({new_AGEMA_signal_1379, AdderIns_g5[18]}), .b ({new_AGEMA_signal_1308, AdderIns_s6_gc_3_a1_t}), .c ({new_AGEMA_signal_1416, AdderIns_g6[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1227, AdderIns_g6[2]}), .b ({new_AGEMA_signal_1262, AdderIns_p5[3]}), .clk (clk), .r (Fresh[243]), .c ({new_AGEMA_signal_1308, AdderIns_s6_gc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_4_a1_U1 ( .a ({new_AGEMA_signal_1380, AdderIns_g5[19]}), .b ({new_AGEMA_signal_1339, AdderIns_s6_gc_4_a1_t}), .c ({new_AGEMA_signal_1417, AdderIns_g6[19]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1277, AdderIns_g6[3]}), .b ({new_AGEMA_signal_1263, AdderIns_p5[4]}), .clk (clk), .r (Fresh[244]), .c ({new_AGEMA_signal_1339, AdderIns_s6_gc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_5_a1_U1 ( .a ({new_AGEMA_signal_1381, AdderIns_g5[20]}), .b ({new_AGEMA_signal_1340, AdderIns_s6_gc_5_a1_t}), .c ({new_AGEMA_signal_1418, AdderIns_g6[20]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1278, AdderIns_g6[4]}), .b ({new_AGEMA_signal_1264, AdderIns_p5[5]}), .clk (clk), .r (Fresh[245]), .c ({new_AGEMA_signal_1340, AdderIns_s6_gc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_6_a1_U1 ( .a ({new_AGEMA_signal_1382, AdderIns_g5[21]}), .b ({new_AGEMA_signal_1341, AdderIns_s6_gc_6_a1_t}), .c ({new_AGEMA_signal_1419, AdderIns_g6[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1279, AdderIns_g6[5]}), .b ({new_AGEMA_signal_1265, AdderIns_p5[6]}), .clk (clk), .r (Fresh[246]), .c ({new_AGEMA_signal_1341, AdderIns_s6_gc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_7_a1_U1 ( .a ({new_AGEMA_signal_1383, AdderIns_g5[22]}), .b ({new_AGEMA_signal_1372, AdderIns_s6_gc_7_a1_t}), .c ({new_AGEMA_signal_1420, AdderIns_g6[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1311, AdderIns_g6[6]}), .b ({new_AGEMA_signal_1266, AdderIns_p5[7]}), .clk (clk), .r (Fresh[247]), .c ({new_AGEMA_signal_1372, AdderIns_s6_gc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_8_a1_U1 ( .a ({new_AGEMA_signal_1384, AdderIns_g5[23]}), .b ({new_AGEMA_signal_1392, AdderIns_s6_gc_8_a1_t}), .c ({new_AGEMA_signal_1421, AdderIns_g6[23]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1348, AdderIns_g6[7]}), .b ({new_AGEMA_signal_1267, AdderIns_p5[8]}), .clk (clk), .r (Fresh[248]), .c ({new_AGEMA_signal_1392, AdderIns_s6_gc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_9_a1_U1 ( .a ({new_AGEMA_signal_1385, AdderIns_g5[24]}), .b ({new_AGEMA_signal_1393, AdderIns_s6_gc_9_a1_t}), .c ({new_AGEMA_signal_1422, AdderIns_g6[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1349, AdderIns_g6[8]}), .b ({new_AGEMA_signal_1268, AdderIns_p5[9]}), .clk (clk), .r (Fresh[249]), .c ({new_AGEMA_signal_1393, AdderIns_s6_gc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_10_a1_U1 ( .a ({new_AGEMA_signal_1386, AdderIns_g5[25]}), .b ({new_AGEMA_signal_1394, AdderIns_s6_gc_10_a1_t}), .c ({new_AGEMA_signal_1423, AdderIns_g6[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1350, AdderIns_g6[9]}), .b ({new_AGEMA_signal_1269, AdderIns_p5[10]}), .clk (clk), .r (Fresh[250]), .c ({new_AGEMA_signal_1394, AdderIns_s6_gc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_11_a1_U1 ( .a ({new_AGEMA_signal_1387, AdderIns_g5[26]}), .b ({new_AGEMA_signal_1395, AdderIns_s6_gc_11_a1_t}), .c ({new_AGEMA_signal_1424, AdderIns_g6[26]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1351, AdderIns_g6[10]}), .b ({new_AGEMA_signal_1270, AdderIns_p5[11]}), .clk (clk), .r (Fresh[251]), .c ({new_AGEMA_signal_1395, AdderIns_s6_gc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_12_a1_U1 ( .a ({new_AGEMA_signal_1388, AdderIns_g5[27]}), .b ({new_AGEMA_signal_1396, AdderIns_s6_gc_12_a1_t}), .c ({new_AGEMA_signal_1425, AdderIns_g6[27]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1352, AdderIns_g6[11]}), .b ({new_AGEMA_signal_1271, AdderIns_p5[12]}), .clk (clk), .r (Fresh[252]), .c ({new_AGEMA_signal_1396, AdderIns_s6_gc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_13_a1_U1 ( .a ({new_AGEMA_signal_1389, AdderIns_g5[28]}), .b ({new_AGEMA_signal_1397, AdderIns_s6_gc_13_a1_t}), .c ({new_AGEMA_signal_1426, AdderIns_g6[28]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1353, AdderIns_g6[12]}), .b ({new_AGEMA_signal_1272, AdderIns_p5[13]}), .clk (clk), .r (Fresh[253]), .c ({new_AGEMA_signal_1397, AdderIns_s6_gc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_14_a1_U1 ( .a ({new_AGEMA_signal_1390, AdderIns_g5[29]}), .b ({new_AGEMA_signal_1398, AdderIns_s6_gc_14_a1_t}), .c ({new_AGEMA_signal_1427, AdderIns_g6[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1354, AdderIns_g6[13]}), .b ({new_AGEMA_signal_1273, AdderIns_p5[14]}), .clk (clk), .r (Fresh[254]), .c ({new_AGEMA_signal_1398, AdderIns_s6_gc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_15_a1_U1 ( .a ({new_AGEMA_signal_1391, AdderIns_g5[30]}), .b ({new_AGEMA_signal_1428, AdderIns_s6_gc_15_a1_t}), .c ({new_AGEMA_signal_1440, AdderIns_g6[30]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s6_gc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1375, AdderIns_g6[14]}), .b ({new_AGEMA_signal_1274, AdderIns_p5[15]}), .clk (clk), .r (Fresh[255]), .c ({new_AGEMA_signal_1428, AdderIns_s6_gc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U24 ( .a ({new_AGEMA_signal_1440, AdderIns_g6[30]}), .b ({new_AGEMA_signal_1046, AdderIns_p6[31]}), .c ({new_AGEMA_signal_1473, sum[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U23 ( .a ({new_AGEMA_signal_1427, AdderIns_g6[29]}), .b ({new_AGEMA_signal_1043, AdderIns_p6[30]}), .c ({new_AGEMA_signal_1441, sum[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U21 ( .a ({new_AGEMA_signal_1426, AdderIns_g6[28]}), .b ({new_AGEMA_signal_1040, AdderIns_p6[29]}), .c ({new_AGEMA_signal_1442, sum[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U20 ( .a ({new_AGEMA_signal_1425, AdderIns_g6[27]}), .b ({new_AGEMA_signal_1037, AdderIns_p6[28]}), .c ({new_AGEMA_signal_1443, sum[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U19 ( .a ({new_AGEMA_signal_1424, AdderIns_g6[26]}), .b ({new_AGEMA_signal_1034, AdderIns_p6[27]}), .c ({new_AGEMA_signal_1444, sum[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U18 ( .a ({new_AGEMA_signal_1423, AdderIns_g6[25]}), .b ({new_AGEMA_signal_1031, AdderIns_p6[26]}), .c ({new_AGEMA_signal_1445, sum[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U17 ( .a ({new_AGEMA_signal_1422, AdderIns_g6[24]}), .b ({new_AGEMA_signal_1028, AdderIns_p6[25]}), .c ({new_AGEMA_signal_1446, sum[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U16 ( .a ({new_AGEMA_signal_1421, AdderIns_g6[23]}), .b ({new_AGEMA_signal_1025, AdderIns_p6[24]}), .c ({new_AGEMA_signal_1447, sum[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U15 ( .a ({new_AGEMA_signal_1420, AdderIns_g6[22]}), .b ({new_AGEMA_signal_1022, AdderIns_p6[23]}), .c ({new_AGEMA_signal_1448, sum[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U14 ( .a ({new_AGEMA_signal_1419, AdderIns_g6[21]}), .b ({new_AGEMA_signal_1019, AdderIns_p6[22]}), .c ({new_AGEMA_signal_1449, sum[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U13 ( .a ({new_AGEMA_signal_1418, AdderIns_g6[20]}), .b ({new_AGEMA_signal_1016, AdderIns_p6[21]}), .c ({new_AGEMA_signal_1450, sum[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U12 ( .a ({new_AGEMA_signal_1417, AdderIns_g6[19]}), .b ({new_AGEMA_signal_1013, AdderIns_p6[20]}), .c ({new_AGEMA_signal_1451, sum[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U10 ( .a ({new_AGEMA_signal_1416, AdderIns_g6[18]}), .b ({new_AGEMA_signal_1010, AdderIns_p6[19]}), .c ({new_AGEMA_signal_1452, sum[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U9 ( .a ({new_AGEMA_signal_1415, AdderIns_g6[17]}), .b ({new_AGEMA_signal_1007, AdderIns_p6[18]}), .c ({new_AGEMA_signal_1453, sum[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U8 ( .a ({new_AGEMA_signal_1414, AdderIns_g6[16]}), .b ({new_AGEMA_signal_1004, AdderIns_p6[17]}), .c ({new_AGEMA_signal_1454, sum[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) AdderIns_s7_U7 ( .a ({new_AGEMA_signal_1376, AdderIns_g6[15]}), .b ({new_AGEMA_signal_1001, AdderIns_p6[16]}), .c ({new_AGEMA_signal_1429, sum[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_0_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1447, sum[24]}), .a ({new_AGEMA_signal_1454, sum[17]}), .c ({new_AGEMA_signal_1474, sum_rotated01[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_1_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1446, sum[25]}), .a ({new_AGEMA_signal_1453, sum[18]}), .c ({new_AGEMA_signal_1475, sum_rotated01[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_2_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1445, sum[26]}), .a ({new_AGEMA_signal_1452, sum[19]}), .c ({new_AGEMA_signal_1476, sum_rotated01[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_3_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1444, sum[27]}), .a ({new_AGEMA_signal_1451, sum[20]}), .c ({new_AGEMA_signal_1477, sum_rotated01[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_4_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1443, sum[28]}), .a ({new_AGEMA_signal_1450, sum[21]}), .c ({new_AGEMA_signal_1478, sum_rotated01[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_5_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1442, sum[29]}), .a ({new_AGEMA_signal_1449, sum[22]}), .c ({new_AGEMA_signal_1479, sum_rotated01[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_6_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1441, sum[30]}), .a ({new_AGEMA_signal_1448, sum[23]}), .c ({new_AGEMA_signal_1480, sum_rotated01[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_7_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1473, sum[31]}), .a ({new_AGEMA_signal_1447, sum[24]}), .c ({new_AGEMA_signal_1527, sum_rotated01[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_8_U1 ( .s (round[0]), .b ({new_AGEMA_signal_953, sum[0]}), .a ({new_AGEMA_signal_1446, sum[25]}), .c ({new_AGEMA_signal_1481, sum_rotated01[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_9_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1225, sum[1]}), .a ({new_AGEMA_signal_1445, sum[26]}), .c ({new_AGEMA_signal_1482, sum_rotated01[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_10_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1275, sum[2]}), .a ({new_AGEMA_signal_1444, sum[27]}), .c ({new_AGEMA_signal_1483, sum_rotated01[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_11_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1309, sum[3]}), .a ({new_AGEMA_signal_1443, sum[28]}), .c ({new_AGEMA_signal_1484, sum_rotated01[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_12_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1344, sum[4]}), .a ({new_AGEMA_signal_1442, sum[29]}), .c ({new_AGEMA_signal_1485, sum_rotated01[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_13_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1343, sum[5]}), .a ({new_AGEMA_signal_1441, sum[30]}), .c ({new_AGEMA_signal_1486, sum_rotated01[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_14_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1342, sum[6]}), .a ({new_AGEMA_signal_1473, sum[31]}), .c ({new_AGEMA_signal_1528, sum_rotated01[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_24_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1429, sum[16]}), .a ({new_AGEMA_signal_1399, sum[9]}), .c ({new_AGEMA_signal_1456, sum_rotated01[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_25_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1454, sum[17]}), .a ({new_AGEMA_signal_1405, sum[10]}), .c ({new_AGEMA_signal_1487, sum_rotated01[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_26_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1453, sum[18]}), .a ({new_AGEMA_signal_1404, sum[11]}), .c ({new_AGEMA_signal_1488, sum_rotated01[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_27_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1452, sum[19]}), .a ({new_AGEMA_signal_1403, sum[12]}), .c ({new_AGEMA_signal_1489, sum_rotated01[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_28_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1451, sum[20]}), .a ({new_AGEMA_signal_1402, sum[13]}), .c ({new_AGEMA_signal_1490, sum_rotated01[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_29_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1450, sum[21]}), .a ({new_AGEMA_signal_1401, sum[14]}), .c ({new_AGEMA_signal_1491, sum_rotated01[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_30_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1449, sum[22]}), .a ({new_AGEMA_signal_1430, sum[15]}), .c ({new_AGEMA_signal_1492, sum_rotated01[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M4_mux_inst_31_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1448, sum[23]}), .a ({new_AGEMA_signal_1429, sum[16]}), .c ({new_AGEMA_signal_1493, sum_rotated01[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_0_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1473, sum[31]}), .a ({new_AGEMA_signal_1429, sum[16]}), .c ({new_AGEMA_signal_1529, sum_rotated23[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_1_U1 ( .s (round[0]), .b ({new_AGEMA_signal_953, sum[0]}), .a ({new_AGEMA_signal_1454, sum[17]}), .c ({new_AGEMA_signal_1494, sum_rotated23[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_2_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1225, sum[1]}), .a ({new_AGEMA_signal_1453, sum[18]}), .c ({new_AGEMA_signal_1495, sum_rotated23[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_3_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1275, sum[2]}), .a ({new_AGEMA_signal_1452, sum[19]}), .c ({new_AGEMA_signal_1496, sum_rotated23[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_4_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1309, sum[3]}), .a ({new_AGEMA_signal_1451, sum[20]}), .c ({new_AGEMA_signal_1497, sum_rotated23[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_5_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1344, sum[4]}), .a ({new_AGEMA_signal_1450, sum[21]}), .c ({new_AGEMA_signal_1498, sum_rotated23[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_6_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1343, sum[5]}), .a ({new_AGEMA_signal_1449, sum[22]}), .c ({new_AGEMA_signal_1499, sum_rotated23[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_7_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1342, sum[6]}), .a ({new_AGEMA_signal_1448, sum[23]}), .c ({new_AGEMA_signal_1500, sum_rotated23[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_8_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1373, sum[7]}), .a ({new_AGEMA_signal_1447, sum[24]}), .c ({new_AGEMA_signal_1501, sum_rotated23[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_9_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1400, sum[8]}), .a ({new_AGEMA_signal_1446, sum[25]}), .c ({new_AGEMA_signal_1502, sum_rotated23[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_10_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1399, sum[9]}), .a ({new_AGEMA_signal_1445, sum[26]}), .c ({new_AGEMA_signal_1503, sum_rotated23[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_11_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1405, sum[10]}), .a ({new_AGEMA_signal_1444, sum[27]}), .c ({new_AGEMA_signal_1504, sum_rotated23[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_12_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1404, sum[11]}), .a ({new_AGEMA_signal_1443, sum[28]}), .c ({new_AGEMA_signal_1505, sum_rotated23[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_13_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1403, sum[12]}), .a ({new_AGEMA_signal_1442, sum[29]}), .c ({new_AGEMA_signal_1506, sum_rotated23[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_14_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1402, sum[13]}), .a ({new_AGEMA_signal_1441, sum[30]}), .c ({new_AGEMA_signal_1507, sum_rotated23[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_15_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1401, sum[14]}), .a ({new_AGEMA_signal_1473, sum[31]}), .c ({new_AGEMA_signal_1530, sum_rotated23[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_17_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1429, sum[16]}), .a ({new_AGEMA_signal_1225, sum[1]}), .c ({new_AGEMA_signal_1458, sum_rotated23[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_18_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1454, sum[17]}), .a ({new_AGEMA_signal_1275, sum[2]}), .c ({new_AGEMA_signal_1508, sum_rotated23[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_19_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1453, sum[18]}), .a ({new_AGEMA_signal_1309, sum[3]}), .c ({new_AGEMA_signal_1509, sum_rotated23[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_20_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1452, sum[19]}), .a ({new_AGEMA_signal_1344, sum[4]}), .c ({new_AGEMA_signal_1510, sum_rotated23[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_21_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1451, sum[20]}), .a ({new_AGEMA_signal_1343, sum[5]}), .c ({new_AGEMA_signal_1511, sum_rotated23[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_22_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1450, sum[21]}), .a ({new_AGEMA_signal_1342, sum[6]}), .c ({new_AGEMA_signal_1512, sum_rotated23[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_23_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1449, sum[22]}), .a ({new_AGEMA_signal_1373, sum[7]}), .c ({new_AGEMA_signal_1513, sum_rotated23[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_24_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1448, sum[23]}), .a ({new_AGEMA_signal_1400, sum[8]}), .c ({new_AGEMA_signal_1514, sum_rotated23[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_25_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1447, sum[24]}), .a ({new_AGEMA_signal_1399, sum[9]}), .c ({new_AGEMA_signal_1515, sum_rotated23[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_26_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1446, sum[25]}), .a ({new_AGEMA_signal_1405, sum[10]}), .c ({new_AGEMA_signal_1516, sum_rotated23[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_27_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1445, sum[26]}), .a ({new_AGEMA_signal_1404, sum[11]}), .c ({new_AGEMA_signal_1517, sum_rotated23[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_28_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1444, sum[27]}), .a ({new_AGEMA_signal_1403, sum[12]}), .c ({new_AGEMA_signal_1518, sum_rotated23[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_29_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1443, sum[28]}), .a ({new_AGEMA_signal_1402, sum[13]}), .c ({new_AGEMA_signal_1519, sum_rotated23[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_30_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1442, sum[29]}), .a ({new_AGEMA_signal_1401, sum[14]}), .c ({new_AGEMA_signal_1520, sum_rotated23[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M5_mux_inst_31_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1441, sum[30]}), .a ({new_AGEMA_signal_1430, sum[15]}), .c ({new_AGEMA_signal_1521, sum_rotated23[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_0_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1474, sum_rotated01[0]}), .a ({new_AGEMA_signal_1529, sum_rotated23[0]}), .c ({new_AGEMA_signal_1583, sum_rotated[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_1_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1475, sum_rotated01[1]}), .a ({new_AGEMA_signal_1494, sum_rotated23[1]}), .c ({new_AGEMA_signal_1531, sum_rotated[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_2_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1476, sum_rotated01[2]}), .a ({new_AGEMA_signal_1495, sum_rotated23[2]}), .c ({new_AGEMA_signal_1532, sum_rotated[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_3_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1477, sum_rotated01[3]}), .a ({new_AGEMA_signal_1496, sum_rotated23[3]}), .c ({new_AGEMA_signal_1533, sum_rotated[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_4_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1478, sum_rotated01[4]}), .a ({new_AGEMA_signal_1497, sum_rotated23[4]}), .c ({new_AGEMA_signal_1534, sum_rotated[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_5_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1479, sum_rotated01[5]}), .a ({new_AGEMA_signal_1498, sum_rotated23[5]}), .c ({new_AGEMA_signal_1535, sum_rotated[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_6_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1480, sum_rotated01[6]}), .a ({new_AGEMA_signal_1499, sum_rotated23[6]}), .c ({new_AGEMA_signal_1536, sum_rotated[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_7_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1527, sum_rotated01[7]}), .a ({new_AGEMA_signal_1500, sum_rotated23[7]}), .c ({new_AGEMA_signal_1584, sum_rotated[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_8_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1481, sum_rotated01[8]}), .a ({new_AGEMA_signal_1501, sum_rotated23[8]}), .c ({new_AGEMA_signal_1537, sum_rotated[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_9_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1482, sum_rotated01[9]}), .a ({new_AGEMA_signal_1502, sum_rotated23[9]}), .c ({new_AGEMA_signal_1538, sum_rotated[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_10_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1483, sum_rotated01[10]}), .a ({new_AGEMA_signal_1503, sum_rotated23[10]}), .c ({new_AGEMA_signal_1539, sum_rotated[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_11_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1484, sum_rotated01[11]}), .a ({new_AGEMA_signal_1504, sum_rotated23[11]}), .c ({new_AGEMA_signal_1540, sum_rotated[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_12_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1485, sum_rotated01[12]}), .a ({new_AGEMA_signal_1505, sum_rotated23[12]}), .c ({new_AGEMA_signal_1541, sum_rotated[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_13_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1486, sum_rotated01[13]}), .a ({new_AGEMA_signal_1506, sum_rotated23[13]}), .c ({new_AGEMA_signal_1542, sum_rotated[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_14_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1528, sum_rotated01[14]}), .a ({new_AGEMA_signal_1507, sum_rotated23[14]}), .c ({new_AGEMA_signal_1585, sum_rotated[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_15_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1406, sum_rotated01[15]}), .a ({new_AGEMA_signal_1530, sum_rotated23[15]}), .c ({new_AGEMA_signal_1586, sum_rotated[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_17_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1432, sum_rotated01[17]}), .a ({new_AGEMA_signal_1458, sum_rotated23[17]}), .c ({new_AGEMA_signal_1523, sum_rotated[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_18_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1433, sum_rotated01[18]}), .a ({new_AGEMA_signal_1508, sum_rotated23[18]}), .c ({new_AGEMA_signal_1543, sum_rotated[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_19_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1434, sum_rotated01[19]}), .a ({new_AGEMA_signal_1509, sum_rotated23[19]}), .c ({new_AGEMA_signal_1544, sum_rotated[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_20_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1435, sum_rotated01[20]}), .a ({new_AGEMA_signal_1510, sum_rotated23[20]}), .c ({new_AGEMA_signal_1545, sum_rotated[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_21_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1436, sum_rotated01[21]}), .a ({new_AGEMA_signal_1511, sum_rotated23[21]}), .c ({new_AGEMA_signal_1546, sum_rotated[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_22_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1437, sum_rotated01[22]}), .a ({new_AGEMA_signal_1512, sum_rotated23[22]}), .c ({new_AGEMA_signal_1547, sum_rotated[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_23_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1455, sum_rotated01[23]}), .a ({new_AGEMA_signal_1513, sum_rotated23[23]}), .c ({new_AGEMA_signal_1548, sum_rotated[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_24_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1456, sum_rotated01[24]}), .a ({new_AGEMA_signal_1514, sum_rotated23[24]}), .c ({new_AGEMA_signal_1549, sum_rotated[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_25_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1487, sum_rotated01[25]}), .a ({new_AGEMA_signal_1515, sum_rotated23[25]}), .c ({new_AGEMA_signal_1550, sum_rotated[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_26_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1488, sum_rotated01[26]}), .a ({new_AGEMA_signal_1516, sum_rotated23[26]}), .c ({new_AGEMA_signal_1551, sum_rotated[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_27_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1489, sum_rotated01[27]}), .a ({new_AGEMA_signal_1517, sum_rotated23[27]}), .c ({new_AGEMA_signal_1552, sum_rotated[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_28_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1490, sum_rotated01[28]}), .a ({new_AGEMA_signal_1518, sum_rotated23[28]}), .c ({new_AGEMA_signal_1553, sum_rotated[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_29_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1491, sum_rotated01[29]}), .a ({new_AGEMA_signal_1519, sum_rotated23[29]}), .c ({new_AGEMA_signal_1554, sum_rotated[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_30_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1492, sum_rotated01[30]}), .a ({new_AGEMA_signal_1520, sum_rotated23[30]}), .c ({new_AGEMA_signal_1555, sum_rotated[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) M6_mux_inst_31_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1493, sum_rotated01[31]}), .a ({new_AGEMA_signal_1521, sum_rotated23[31]}), .c ({new_AGEMA_signal_1556, sum_rotated[31]}) ) ;

endmodule
