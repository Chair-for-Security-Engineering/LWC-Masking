/* modified netlist. Source: module SubCells in file ./test/SubCells.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module SubCells_HPC2_ClockGating_d3 (SubC_in_s0, clk, SubC_in_s1, SubC_in_s2, SubC_in_s3, Fresh, /*rst,*/ SubC_out_s0, SubC_out_s1, SubC_out_s2, SubC_out_s3/*, Synch*/);
    input [127:0] SubC_in_s0 ;
    input clk ;
    input [127:0] SubC_in_s1 ;
    input [127:0] SubC_in_s2 ;
    input [127:0] SubC_in_s3 ;
    //input rst ;
    input [1151:0] Fresh ;
    output [127:0] SubC_out_s0 ;
    output [127:0] SubC_out_s1 ;
    output [127:0] SubC_out_s2 ;
    output [127:0] SubC_out_s3 ;
    //output Synch ;
    wire SB_31_n15 ;
    wire SB_31_n14 ;
    wire SB_31_n13 ;
    wire SB_31_n12 ;
    wire SB_31_n11 ;
    wire SB_31_n10 ;
    wire SB_31_n9 ;
    wire SB_31_T5 ;
    wire SB_31_T4 ;
    wire SB_31_T3 ;
    wire SB_31_T2 ;
    wire SB_31_T1 ;
    wire SB_31_T0 ;
    wire SB_30_n15 ;
    wire SB_30_n14 ;
    wire SB_30_n13 ;
    wire SB_30_n12 ;
    wire SB_30_n11 ;
    wire SB_30_n10 ;
    wire SB_30_n9 ;
    wire SB_30_T5 ;
    wire SB_30_T4 ;
    wire SB_30_T3 ;
    wire SB_30_T2 ;
    wire SB_30_T1 ;
    wire SB_30_T0 ;
    wire SB_29_n15 ;
    wire SB_29_n14 ;
    wire SB_29_n13 ;
    wire SB_29_n12 ;
    wire SB_29_n11 ;
    wire SB_29_n10 ;
    wire SB_29_n9 ;
    wire SB_29_T5 ;
    wire SB_29_T4 ;
    wire SB_29_T3 ;
    wire SB_29_T2 ;
    wire SB_29_T1 ;
    wire SB_29_T0 ;
    wire SB_28_n15 ;
    wire SB_28_n14 ;
    wire SB_28_n13 ;
    wire SB_28_n12 ;
    wire SB_28_n11 ;
    wire SB_28_n10 ;
    wire SB_28_n9 ;
    wire SB_28_T5 ;
    wire SB_28_T4 ;
    wire SB_28_T3 ;
    wire SB_28_T2 ;
    wire SB_28_T1 ;
    wire SB_28_T0 ;
    wire SB_27_n15 ;
    wire SB_27_n14 ;
    wire SB_27_n13 ;
    wire SB_27_n12 ;
    wire SB_27_n11 ;
    wire SB_27_n10 ;
    wire SB_27_n9 ;
    wire SB_27_T5 ;
    wire SB_27_T4 ;
    wire SB_27_T3 ;
    wire SB_27_T2 ;
    wire SB_27_T1 ;
    wire SB_27_T0 ;
    wire SB_26_n15 ;
    wire SB_26_n14 ;
    wire SB_26_n13 ;
    wire SB_26_n12 ;
    wire SB_26_n11 ;
    wire SB_26_n10 ;
    wire SB_26_n9 ;
    wire SB_26_T5 ;
    wire SB_26_T4 ;
    wire SB_26_T3 ;
    wire SB_26_T2 ;
    wire SB_26_T1 ;
    wire SB_26_T0 ;
    wire SB_25_n15 ;
    wire SB_25_n14 ;
    wire SB_25_n13 ;
    wire SB_25_n12 ;
    wire SB_25_n11 ;
    wire SB_25_n10 ;
    wire SB_25_n9 ;
    wire SB_25_T5 ;
    wire SB_25_T4 ;
    wire SB_25_T3 ;
    wire SB_25_T2 ;
    wire SB_25_T1 ;
    wire SB_25_T0 ;
    wire SB_24_n15 ;
    wire SB_24_n14 ;
    wire SB_24_n13 ;
    wire SB_24_n12 ;
    wire SB_24_n11 ;
    wire SB_24_n10 ;
    wire SB_24_n9 ;
    wire SB_24_T5 ;
    wire SB_24_T4 ;
    wire SB_24_T3 ;
    wire SB_24_T2 ;
    wire SB_24_T1 ;
    wire SB_24_T0 ;
    wire SB_23_n15 ;
    wire SB_23_n14 ;
    wire SB_23_n13 ;
    wire SB_23_n12 ;
    wire SB_23_n11 ;
    wire SB_23_n10 ;
    wire SB_23_n9 ;
    wire SB_23_T5 ;
    wire SB_23_T4 ;
    wire SB_23_T3 ;
    wire SB_23_T2 ;
    wire SB_23_T1 ;
    wire SB_23_T0 ;
    wire SB_22_n15 ;
    wire SB_22_n14 ;
    wire SB_22_n13 ;
    wire SB_22_n12 ;
    wire SB_22_n11 ;
    wire SB_22_n10 ;
    wire SB_22_n9 ;
    wire SB_22_T5 ;
    wire SB_22_T4 ;
    wire SB_22_T3 ;
    wire SB_22_T2 ;
    wire SB_22_T1 ;
    wire SB_22_T0 ;
    wire SB_21_n15 ;
    wire SB_21_n14 ;
    wire SB_21_n13 ;
    wire SB_21_n12 ;
    wire SB_21_n11 ;
    wire SB_21_n10 ;
    wire SB_21_n9 ;
    wire SB_21_T5 ;
    wire SB_21_T4 ;
    wire SB_21_T3 ;
    wire SB_21_T2 ;
    wire SB_21_T1 ;
    wire SB_21_T0 ;
    wire SB_20_n15 ;
    wire SB_20_n14 ;
    wire SB_20_n13 ;
    wire SB_20_n12 ;
    wire SB_20_n11 ;
    wire SB_20_n10 ;
    wire SB_20_n9 ;
    wire SB_20_T5 ;
    wire SB_20_T4 ;
    wire SB_20_T3 ;
    wire SB_20_T2 ;
    wire SB_20_T1 ;
    wire SB_20_T0 ;
    wire SB_19_n15 ;
    wire SB_19_n14 ;
    wire SB_19_n13 ;
    wire SB_19_n12 ;
    wire SB_19_n11 ;
    wire SB_19_n10 ;
    wire SB_19_n9 ;
    wire SB_19_T5 ;
    wire SB_19_T4 ;
    wire SB_19_T3 ;
    wire SB_19_T2 ;
    wire SB_19_T1 ;
    wire SB_19_T0 ;
    wire SB_18_n15 ;
    wire SB_18_n14 ;
    wire SB_18_n13 ;
    wire SB_18_n12 ;
    wire SB_18_n11 ;
    wire SB_18_n10 ;
    wire SB_18_n9 ;
    wire SB_18_T5 ;
    wire SB_18_T4 ;
    wire SB_18_T3 ;
    wire SB_18_T2 ;
    wire SB_18_T1 ;
    wire SB_18_T0 ;
    wire SB_17_n15 ;
    wire SB_17_n14 ;
    wire SB_17_n13 ;
    wire SB_17_n12 ;
    wire SB_17_n11 ;
    wire SB_17_n10 ;
    wire SB_17_n9 ;
    wire SB_17_T5 ;
    wire SB_17_T4 ;
    wire SB_17_T3 ;
    wire SB_17_T2 ;
    wire SB_17_T1 ;
    wire SB_17_T0 ;
    wire SB_16_n15 ;
    wire SB_16_n14 ;
    wire SB_16_n13 ;
    wire SB_16_n12 ;
    wire SB_16_n11 ;
    wire SB_16_n10 ;
    wire SB_16_n9 ;
    wire SB_16_T5 ;
    wire SB_16_T4 ;
    wire SB_16_T3 ;
    wire SB_16_T2 ;
    wire SB_16_T1 ;
    wire SB_16_T0 ;
    wire SB_15_n15 ;
    wire SB_15_n14 ;
    wire SB_15_n13 ;
    wire SB_15_n12 ;
    wire SB_15_n11 ;
    wire SB_15_n10 ;
    wire SB_15_n9 ;
    wire SB_15_T5 ;
    wire SB_15_T4 ;
    wire SB_15_T3 ;
    wire SB_15_T2 ;
    wire SB_15_T1 ;
    wire SB_15_T0 ;
    wire SB_14_n15 ;
    wire SB_14_n14 ;
    wire SB_14_n13 ;
    wire SB_14_n12 ;
    wire SB_14_n11 ;
    wire SB_14_n10 ;
    wire SB_14_n9 ;
    wire SB_14_T5 ;
    wire SB_14_T4 ;
    wire SB_14_T3 ;
    wire SB_14_T2 ;
    wire SB_14_T1 ;
    wire SB_14_T0 ;
    wire SB_13_n15 ;
    wire SB_13_n14 ;
    wire SB_13_n13 ;
    wire SB_13_n12 ;
    wire SB_13_n11 ;
    wire SB_13_n10 ;
    wire SB_13_n9 ;
    wire SB_13_T5 ;
    wire SB_13_T4 ;
    wire SB_13_T3 ;
    wire SB_13_T2 ;
    wire SB_13_T1 ;
    wire SB_13_T0 ;
    wire SB_12_n15 ;
    wire SB_12_n14 ;
    wire SB_12_n13 ;
    wire SB_12_n12 ;
    wire SB_12_n11 ;
    wire SB_12_n10 ;
    wire SB_12_n9 ;
    wire SB_12_T5 ;
    wire SB_12_T4 ;
    wire SB_12_T3 ;
    wire SB_12_T2 ;
    wire SB_12_T1 ;
    wire SB_12_T0 ;
    wire SB_11_n15 ;
    wire SB_11_n14 ;
    wire SB_11_n13 ;
    wire SB_11_n12 ;
    wire SB_11_n11 ;
    wire SB_11_n10 ;
    wire SB_11_n9 ;
    wire SB_11_T5 ;
    wire SB_11_T4 ;
    wire SB_11_T3 ;
    wire SB_11_T2 ;
    wire SB_11_T1 ;
    wire SB_11_T0 ;
    wire SB_10_n15 ;
    wire SB_10_n14 ;
    wire SB_10_n13 ;
    wire SB_10_n12 ;
    wire SB_10_n11 ;
    wire SB_10_n10 ;
    wire SB_10_n9 ;
    wire SB_10_T5 ;
    wire SB_10_T4 ;
    wire SB_10_T3 ;
    wire SB_10_T2 ;
    wire SB_10_T1 ;
    wire SB_10_T0 ;
    wire SB_9_n15 ;
    wire SB_9_n14 ;
    wire SB_9_n13 ;
    wire SB_9_n12 ;
    wire SB_9_n11 ;
    wire SB_9_n10 ;
    wire SB_9_n9 ;
    wire SB_9_T5 ;
    wire SB_9_T4 ;
    wire SB_9_T3 ;
    wire SB_9_T2 ;
    wire SB_9_T1 ;
    wire SB_9_T0 ;
    wire SB_8_n15 ;
    wire SB_8_n14 ;
    wire SB_8_n13 ;
    wire SB_8_n12 ;
    wire SB_8_n11 ;
    wire SB_8_n10 ;
    wire SB_8_n9 ;
    wire SB_8_T5 ;
    wire SB_8_T4 ;
    wire SB_8_T3 ;
    wire SB_8_T2 ;
    wire SB_8_T1 ;
    wire SB_8_T0 ;
    wire SB_7_n15 ;
    wire SB_7_n14 ;
    wire SB_7_n13 ;
    wire SB_7_n12 ;
    wire SB_7_n11 ;
    wire SB_7_n10 ;
    wire SB_7_n9 ;
    wire SB_7_T5 ;
    wire SB_7_T4 ;
    wire SB_7_T3 ;
    wire SB_7_T2 ;
    wire SB_7_T1 ;
    wire SB_7_T0 ;
    wire SB_6_n15 ;
    wire SB_6_n14 ;
    wire SB_6_n13 ;
    wire SB_6_n12 ;
    wire SB_6_n11 ;
    wire SB_6_n10 ;
    wire SB_6_n9 ;
    wire SB_6_T5 ;
    wire SB_6_T4 ;
    wire SB_6_T3 ;
    wire SB_6_T2 ;
    wire SB_6_T1 ;
    wire SB_6_T0 ;
    wire SB_5_n15 ;
    wire SB_5_n14 ;
    wire SB_5_n13 ;
    wire SB_5_n12 ;
    wire SB_5_n11 ;
    wire SB_5_n10 ;
    wire SB_5_n9 ;
    wire SB_5_T5 ;
    wire SB_5_T4 ;
    wire SB_5_T3 ;
    wire SB_5_T2 ;
    wire SB_5_T1 ;
    wire SB_5_T0 ;
    wire SB_4_n15 ;
    wire SB_4_n14 ;
    wire SB_4_n13 ;
    wire SB_4_n12 ;
    wire SB_4_n11 ;
    wire SB_4_n10 ;
    wire SB_4_n9 ;
    wire SB_4_T5 ;
    wire SB_4_T4 ;
    wire SB_4_T3 ;
    wire SB_4_T2 ;
    wire SB_4_T1 ;
    wire SB_4_T0 ;
    wire SB_3_n15 ;
    wire SB_3_n14 ;
    wire SB_3_n13 ;
    wire SB_3_n12 ;
    wire SB_3_n11 ;
    wire SB_3_n10 ;
    wire SB_3_n9 ;
    wire SB_3_T5 ;
    wire SB_3_T4 ;
    wire SB_3_T3 ;
    wire SB_3_T2 ;
    wire SB_3_T1 ;
    wire SB_3_T0 ;
    wire SB_2_n15 ;
    wire SB_2_n14 ;
    wire SB_2_n13 ;
    wire SB_2_n12 ;
    wire SB_2_n11 ;
    wire SB_2_n10 ;
    wire SB_2_n9 ;
    wire SB_2_T5 ;
    wire SB_2_T4 ;
    wire SB_2_T3 ;
    wire SB_2_T2 ;
    wire SB_2_T1 ;
    wire SB_2_T0 ;
    wire SB_1_n15 ;
    wire SB_1_n14 ;
    wire SB_1_n13 ;
    wire SB_1_n12 ;
    wire SB_1_n11 ;
    wire SB_1_n10 ;
    wire SB_1_n9 ;
    wire SB_1_T5 ;
    wire SB_1_T4 ;
    wire SB_1_T3 ;
    wire SB_1_T2 ;
    wire SB_1_T1 ;
    wire SB_1_T0 ;
    wire SB_0_n15 ;
    wire SB_0_n14 ;
    wire SB_0_n13 ;
    wire SB_0_n12 ;
    wire SB_0_n11 ;
    wire SB_0_n10 ;
    wire SB_0_n9 ;
    wire SB_0_T5 ;
    wire SB_0_T4 ;
    wire SB_0_T3 ;
    wire SB_0_T2 ;
    wire SB_0_T1 ;
    wire SB_0_T0 ;
    wire new_AGEMA_signal_685 ;
    wire new_AGEMA_signal_686 ;
    wire new_AGEMA_signal_687 ;
    wire new_AGEMA_signal_694 ;
    wire new_AGEMA_signal_695 ;
    wire new_AGEMA_signal_696 ;
    wire new_AGEMA_signal_697 ;
    wire new_AGEMA_signal_698 ;
    wire new_AGEMA_signal_699 ;
    wire new_AGEMA_signal_700 ;
    wire new_AGEMA_signal_701 ;
    wire new_AGEMA_signal_702 ;
    wire new_AGEMA_signal_703 ;
    wire new_AGEMA_signal_704 ;
    wire new_AGEMA_signal_705 ;
    wire new_AGEMA_signal_706 ;
    wire new_AGEMA_signal_707 ;
    wire new_AGEMA_signal_708 ;
    wire new_AGEMA_signal_715 ;
    wire new_AGEMA_signal_716 ;
    wire new_AGEMA_signal_717 ;
    wire new_AGEMA_signal_724 ;
    wire new_AGEMA_signal_725 ;
    wire new_AGEMA_signal_726 ;
    wire new_AGEMA_signal_727 ;
    wire new_AGEMA_signal_728 ;
    wire new_AGEMA_signal_729 ;
    wire new_AGEMA_signal_730 ;
    wire new_AGEMA_signal_731 ;
    wire new_AGEMA_signal_732 ;
    wire new_AGEMA_signal_733 ;
    wire new_AGEMA_signal_734 ;
    wire new_AGEMA_signal_735 ;
    wire new_AGEMA_signal_736 ;
    wire new_AGEMA_signal_737 ;
    wire new_AGEMA_signal_738 ;
    wire new_AGEMA_signal_745 ;
    wire new_AGEMA_signal_746 ;
    wire new_AGEMA_signal_747 ;
    wire new_AGEMA_signal_754 ;
    wire new_AGEMA_signal_755 ;
    wire new_AGEMA_signal_756 ;
    wire new_AGEMA_signal_757 ;
    wire new_AGEMA_signal_758 ;
    wire new_AGEMA_signal_759 ;
    wire new_AGEMA_signal_760 ;
    wire new_AGEMA_signal_761 ;
    wire new_AGEMA_signal_762 ;
    wire new_AGEMA_signal_763 ;
    wire new_AGEMA_signal_764 ;
    wire new_AGEMA_signal_765 ;
    wire new_AGEMA_signal_766 ;
    wire new_AGEMA_signal_767 ;
    wire new_AGEMA_signal_768 ;
    wire new_AGEMA_signal_775 ;
    wire new_AGEMA_signal_776 ;
    wire new_AGEMA_signal_777 ;
    wire new_AGEMA_signal_784 ;
    wire new_AGEMA_signal_785 ;
    wire new_AGEMA_signal_786 ;
    wire new_AGEMA_signal_787 ;
    wire new_AGEMA_signal_788 ;
    wire new_AGEMA_signal_789 ;
    wire new_AGEMA_signal_790 ;
    wire new_AGEMA_signal_791 ;
    wire new_AGEMA_signal_792 ;
    wire new_AGEMA_signal_793 ;
    wire new_AGEMA_signal_794 ;
    wire new_AGEMA_signal_795 ;
    wire new_AGEMA_signal_796 ;
    wire new_AGEMA_signal_797 ;
    wire new_AGEMA_signal_798 ;
    wire new_AGEMA_signal_805 ;
    wire new_AGEMA_signal_806 ;
    wire new_AGEMA_signal_807 ;
    wire new_AGEMA_signal_814 ;
    wire new_AGEMA_signal_815 ;
    wire new_AGEMA_signal_816 ;
    wire new_AGEMA_signal_817 ;
    wire new_AGEMA_signal_818 ;
    wire new_AGEMA_signal_819 ;
    wire new_AGEMA_signal_820 ;
    wire new_AGEMA_signal_821 ;
    wire new_AGEMA_signal_822 ;
    wire new_AGEMA_signal_823 ;
    wire new_AGEMA_signal_824 ;
    wire new_AGEMA_signal_825 ;
    wire new_AGEMA_signal_826 ;
    wire new_AGEMA_signal_827 ;
    wire new_AGEMA_signal_828 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_836 ;
    wire new_AGEMA_signal_837 ;
    wire new_AGEMA_signal_844 ;
    wire new_AGEMA_signal_845 ;
    wire new_AGEMA_signal_846 ;
    wire new_AGEMA_signal_847 ;
    wire new_AGEMA_signal_848 ;
    wire new_AGEMA_signal_849 ;
    wire new_AGEMA_signal_850 ;
    wire new_AGEMA_signal_851 ;
    wire new_AGEMA_signal_852 ;
    wire new_AGEMA_signal_853 ;
    wire new_AGEMA_signal_854 ;
    wire new_AGEMA_signal_855 ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_857 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_874 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_878 ;
    wire new_AGEMA_signal_879 ;
    wire new_AGEMA_signal_880 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_886 ;
    wire new_AGEMA_signal_887 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_896 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_904 ;
    wire new_AGEMA_signal_905 ;
    wire new_AGEMA_signal_906 ;
    wire new_AGEMA_signal_907 ;
    wire new_AGEMA_signal_908 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_910 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_912 ;
    wire new_AGEMA_signal_913 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_915 ;
    wire new_AGEMA_signal_916 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_934 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_939 ;
    wire new_AGEMA_signal_940 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_942 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U8 ( .a ({SubC_in_s3[63], SubC_in_s2[63], SubC_in_s1[63], SubC_in_s0[63]}), .b ({SubC_in_s3[95], SubC_in_s2[95], SubC_in_s1[95], SubC_in_s0[95]}), .c ({new_AGEMA_signal_687, new_AGEMA_signal_686, new_AGEMA_signal_685, SB_31_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U3 ( .a ({SubC_in_s3[31], SubC_in_s2[31], SubC_in_s1[31], SubC_in_s0[31]}), .b ({SubC_in_s3[127], SubC_in_s2[127], SubC_in_s1[127], SubC_in_s0[127]}), .c ({new_AGEMA_signal_696, new_AGEMA_signal_695, new_AGEMA_signal_694, SB_31_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U8 ( .a ({SubC_in_s3[62], SubC_in_s2[62], SubC_in_s1[62], SubC_in_s0[62]}), .b ({SubC_in_s3[94], SubC_in_s2[94], SubC_in_s1[94], SubC_in_s0[94]}), .c ({new_AGEMA_signal_717, new_AGEMA_signal_716, new_AGEMA_signal_715, SB_30_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U3 ( .a ({SubC_in_s3[30], SubC_in_s2[30], SubC_in_s1[30], SubC_in_s0[30]}), .b ({SubC_in_s3[126], SubC_in_s2[126], SubC_in_s1[126], SubC_in_s0[126]}), .c ({new_AGEMA_signal_726, new_AGEMA_signal_725, new_AGEMA_signal_724, SB_30_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U8 ( .a ({SubC_in_s3[61], SubC_in_s2[61], SubC_in_s1[61], SubC_in_s0[61]}), .b ({SubC_in_s3[93], SubC_in_s2[93], SubC_in_s1[93], SubC_in_s0[93]}), .c ({new_AGEMA_signal_747, new_AGEMA_signal_746, new_AGEMA_signal_745, SB_29_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U3 ( .a ({SubC_in_s3[29], SubC_in_s2[29], SubC_in_s1[29], SubC_in_s0[29]}), .b ({SubC_in_s3[125], SubC_in_s2[125], SubC_in_s1[125], SubC_in_s0[125]}), .c ({new_AGEMA_signal_756, new_AGEMA_signal_755, new_AGEMA_signal_754, SB_29_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U8 ( .a ({SubC_in_s3[60], SubC_in_s2[60], SubC_in_s1[60], SubC_in_s0[60]}), .b ({SubC_in_s3[92], SubC_in_s2[92], SubC_in_s1[92], SubC_in_s0[92]}), .c ({new_AGEMA_signal_777, new_AGEMA_signal_776, new_AGEMA_signal_775, SB_28_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U3 ( .a ({SubC_in_s3[28], SubC_in_s2[28], SubC_in_s1[28], SubC_in_s0[28]}), .b ({SubC_in_s3[124], SubC_in_s2[124], SubC_in_s1[124], SubC_in_s0[124]}), .c ({new_AGEMA_signal_786, new_AGEMA_signal_785, new_AGEMA_signal_784, SB_28_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U8 ( .a ({SubC_in_s3[59], SubC_in_s2[59], SubC_in_s1[59], SubC_in_s0[59]}), .b ({SubC_in_s3[91], SubC_in_s2[91], SubC_in_s1[91], SubC_in_s0[91]}), .c ({new_AGEMA_signal_807, new_AGEMA_signal_806, new_AGEMA_signal_805, SB_27_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U3 ( .a ({SubC_in_s3[27], SubC_in_s2[27], SubC_in_s1[27], SubC_in_s0[27]}), .b ({SubC_in_s3[123], SubC_in_s2[123], SubC_in_s1[123], SubC_in_s0[123]}), .c ({new_AGEMA_signal_816, new_AGEMA_signal_815, new_AGEMA_signal_814, SB_27_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U8 ( .a ({SubC_in_s3[58], SubC_in_s2[58], SubC_in_s1[58], SubC_in_s0[58]}), .b ({SubC_in_s3[90], SubC_in_s2[90], SubC_in_s1[90], SubC_in_s0[90]}), .c ({new_AGEMA_signal_837, new_AGEMA_signal_836, new_AGEMA_signal_835, SB_26_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U3 ( .a ({SubC_in_s3[26], SubC_in_s2[26], SubC_in_s1[26], SubC_in_s0[26]}), .b ({SubC_in_s3[122], SubC_in_s2[122], SubC_in_s1[122], SubC_in_s0[122]}), .c ({new_AGEMA_signal_846, new_AGEMA_signal_845, new_AGEMA_signal_844, SB_26_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U8 ( .a ({SubC_in_s3[57], SubC_in_s2[57], SubC_in_s1[57], SubC_in_s0[57]}), .b ({SubC_in_s3[89], SubC_in_s2[89], SubC_in_s1[89], SubC_in_s0[89]}), .c ({new_AGEMA_signal_867, new_AGEMA_signal_866, new_AGEMA_signal_865, SB_25_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U3 ( .a ({SubC_in_s3[25], SubC_in_s2[25], SubC_in_s1[25], SubC_in_s0[25]}), .b ({SubC_in_s3[121], SubC_in_s2[121], SubC_in_s1[121], SubC_in_s0[121]}), .c ({new_AGEMA_signal_876, new_AGEMA_signal_875, new_AGEMA_signal_874, SB_25_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U8 ( .a ({SubC_in_s3[56], SubC_in_s2[56], SubC_in_s1[56], SubC_in_s0[56]}), .b ({SubC_in_s3[88], SubC_in_s2[88], SubC_in_s1[88], SubC_in_s0[88]}), .c ({new_AGEMA_signal_897, new_AGEMA_signal_896, new_AGEMA_signal_895, SB_24_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U3 ( .a ({SubC_in_s3[24], SubC_in_s2[24], SubC_in_s1[24], SubC_in_s0[24]}), .b ({SubC_in_s3[120], SubC_in_s2[120], SubC_in_s1[120], SubC_in_s0[120]}), .c ({new_AGEMA_signal_906, new_AGEMA_signal_905, new_AGEMA_signal_904, SB_24_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U8 ( .a ({SubC_in_s3[55], SubC_in_s2[55], SubC_in_s1[55], SubC_in_s0[55]}), .b ({SubC_in_s3[87], SubC_in_s2[87], SubC_in_s1[87], SubC_in_s0[87]}), .c ({new_AGEMA_signal_927, new_AGEMA_signal_926, new_AGEMA_signal_925, SB_23_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U3 ( .a ({SubC_in_s3[23], SubC_in_s2[23], SubC_in_s1[23], SubC_in_s0[23]}), .b ({SubC_in_s3[119], SubC_in_s2[119], SubC_in_s1[119], SubC_in_s0[119]}), .c ({new_AGEMA_signal_936, new_AGEMA_signal_935, new_AGEMA_signal_934, SB_23_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U8 ( .a ({SubC_in_s3[54], SubC_in_s2[54], SubC_in_s1[54], SubC_in_s0[54]}), .b ({SubC_in_s3[86], SubC_in_s2[86], SubC_in_s1[86], SubC_in_s0[86]}), .c ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, SB_22_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U3 ( .a ({SubC_in_s3[22], SubC_in_s2[22], SubC_in_s1[22], SubC_in_s0[22]}), .b ({SubC_in_s3[118], SubC_in_s2[118], SubC_in_s1[118], SubC_in_s0[118]}), .c ({new_AGEMA_signal_966, new_AGEMA_signal_965, new_AGEMA_signal_964, SB_22_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U8 ( .a ({SubC_in_s3[53], SubC_in_s2[53], SubC_in_s1[53], SubC_in_s0[53]}), .b ({SubC_in_s3[85], SubC_in_s2[85], SubC_in_s1[85], SubC_in_s0[85]}), .c ({new_AGEMA_signal_987, new_AGEMA_signal_986, new_AGEMA_signal_985, SB_21_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U3 ( .a ({SubC_in_s3[21], SubC_in_s2[21], SubC_in_s1[21], SubC_in_s0[21]}), .b ({SubC_in_s3[117], SubC_in_s2[117], SubC_in_s1[117], SubC_in_s0[117]}), .c ({new_AGEMA_signal_996, new_AGEMA_signal_995, new_AGEMA_signal_994, SB_21_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U8 ( .a ({SubC_in_s3[52], SubC_in_s2[52], SubC_in_s1[52], SubC_in_s0[52]}), .b ({SubC_in_s3[84], SubC_in_s2[84], SubC_in_s1[84], SubC_in_s0[84]}), .c ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, SB_20_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U3 ( .a ({SubC_in_s3[20], SubC_in_s2[20], SubC_in_s1[20], SubC_in_s0[20]}), .b ({SubC_in_s3[116], SubC_in_s2[116], SubC_in_s1[116], SubC_in_s0[116]}), .c ({new_AGEMA_signal_1026, new_AGEMA_signal_1025, new_AGEMA_signal_1024, SB_20_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U8 ( .a ({SubC_in_s3[51], SubC_in_s2[51], SubC_in_s1[51], SubC_in_s0[51]}), .b ({SubC_in_s3[83], SubC_in_s2[83], SubC_in_s1[83], SubC_in_s0[83]}), .c ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, new_AGEMA_signal_1045, SB_19_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U3 ( .a ({SubC_in_s3[19], SubC_in_s2[19], SubC_in_s1[19], SubC_in_s0[19]}), .b ({SubC_in_s3[115], SubC_in_s2[115], SubC_in_s1[115], SubC_in_s0[115]}), .c ({new_AGEMA_signal_1056, new_AGEMA_signal_1055, new_AGEMA_signal_1054, SB_19_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U8 ( .a ({SubC_in_s3[50], SubC_in_s2[50], SubC_in_s1[50], SubC_in_s0[50]}), .b ({SubC_in_s3[82], SubC_in_s2[82], SubC_in_s1[82], SubC_in_s0[82]}), .c ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, SB_18_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U3 ( .a ({SubC_in_s3[18], SubC_in_s2[18], SubC_in_s1[18], SubC_in_s0[18]}), .b ({SubC_in_s3[114], SubC_in_s2[114], SubC_in_s1[114], SubC_in_s0[114]}), .c ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, SB_18_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U8 ( .a ({SubC_in_s3[49], SubC_in_s2[49], SubC_in_s1[49], SubC_in_s0[49]}), .b ({SubC_in_s3[81], SubC_in_s2[81], SubC_in_s1[81], SubC_in_s0[81]}), .c ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, new_AGEMA_signal_1105, SB_17_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U3 ( .a ({SubC_in_s3[17], SubC_in_s2[17], SubC_in_s1[17], SubC_in_s0[17]}), .b ({SubC_in_s3[113], SubC_in_s2[113], SubC_in_s1[113], SubC_in_s0[113]}), .c ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, new_AGEMA_signal_1114, SB_17_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U8 ( .a ({SubC_in_s3[48], SubC_in_s2[48], SubC_in_s1[48], SubC_in_s0[48]}), .b ({SubC_in_s3[80], SubC_in_s2[80], SubC_in_s1[80], SubC_in_s0[80]}), .c ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, new_AGEMA_signal_1135, SB_16_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U3 ( .a ({SubC_in_s3[16], SubC_in_s2[16], SubC_in_s1[16], SubC_in_s0[16]}), .b ({SubC_in_s3[112], SubC_in_s2[112], SubC_in_s1[112], SubC_in_s0[112]}), .c ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, new_AGEMA_signal_1144, SB_16_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U8 ( .a ({SubC_in_s3[47], SubC_in_s2[47], SubC_in_s1[47], SubC_in_s0[47]}), .b ({SubC_in_s3[79], SubC_in_s2[79], SubC_in_s1[79], SubC_in_s0[79]}), .c ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, new_AGEMA_signal_1165, SB_15_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U3 ( .a ({SubC_in_s3[15], SubC_in_s2[15], SubC_in_s1[15], SubC_in_s0[15]}), .b ({SubC_in_s3[111], SubC_in_s2[111], SubC_in_s1[111], SubC_in_s0[111]}), .c ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, new_AGEMA_signal_1174, SB_15_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U8 ( .a ({SubC_in_s3[46], SubC_in_s2[46], SubC_in_s1[46], SubC_in_s0[46]}), .b ({SubC_in_s3[78], SubC_in_s2[78], SubC_in_s1[78], SubC_in_s0[78]}), .c ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, SB_14_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U3 ( .a ({SubC_in_s3[14], SubC_in_s2[14], SubC_in_s1[14], SubC_in_s0[14]}), .b ({SubC_in_s3[110], SubC_in_s2[110], SubC_in_s1[110], SubC_in_s0[110]}), .c ({new_AGEMA_signal_1206, new_AGEMA_signal_1205, new_AGEMA_signal_1204, SB_14_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U8 ( .a ({SubC_in_s3[45], SubC_in_s2[45], SubC_in_s1[45], SubC_in_s0[45]}), .b ({SubC_in_s3[77], SubC_in_s2[77], SubC_in_s1[77], SubC_in_s0[77]}), .c ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, new_AGEMA_signal_1225, SB_13_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U3 ( .a ({SubC_in_s3[13], SubC_in_s2[13], SubC_in_s1[13], SubC_in_s0[13]}), .b ({SubC_in_s3[109], SubC_in_s2[109], SubC_in_s1[109], SubC_in_s0[109]}), .c ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, new_AGEMA_signal_1234, SB_13_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U8 ( .a ({SubC_in_s3[44], SubC_in_s2[44], SubC_in_s1[44], SubC_in_s0[44]}), .b ({SubC_in_s3[76], SubC_in_s2[76], SubC_in_s1[76], SubC_in_s0[76]}), .c ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, new_AGEMA_signal_1255, SB_12_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U3 ( .a ({SubC_in_s3[12], SubC_in_s2[12], SubC_in_s1[12], SubC_in_s0[12]}), .b ({SubC_in_s3[108], SubC_in_s2[108], SubC_in_s1[108], SubC_in_s0[108]}), .c ({new_AGEMA_signal_1266, new_AGEMA_signal_1265, new_AGEMA_signal_1264, SB_12_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U8 ( .a ({SubC_in_s3[43], SubC_in_s2[43], SubC_in_s1[43], SubC_in_s0[43]}), .b ({SubC_in_s3[75], SubC_in_s2[75], SubC_in_s1[75], SubC_in_s0[75]}), .c ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, new_AGEMA_signal_1285, SB_11_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U3 ( .a ({SubC_in_s3[11], SubC_in_s2[11], SubC_in_s1[11], SubC_in_s0[11]}), .b ({SubC_in_s3[107], SubC_in_s2[107], SubC_in_s1[107], SubC_in_s0[107]}), .c ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, new_AGEMA_signal_1294, SB_11_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U8 ( .a ({SubC_in_s3[42], SubC_in_s2[42], SubC_in_s1[42], SubC_in_s0[42]}), .b ({SubC_in_s3[74], SubC_in_s2[74], SubC_in_s1[74], SubC_in_s0[74]}), .c ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, SB_10_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U3 ( .a ({SubC_in_s3[10], SubC_in_s2[10], SubC_in_s1[10], SubC_in_s0[10]}), .b ({SubC_in_s3[106], SubC_in_s2[106], SubC_in_s1[106], SubC_in_s0[106]}), .c ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, new_AGEMA_signal_1324, SB_10_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U8 ( .a ({SubC_in_s3[41], SubC_in_s2[41], SubC_in_s1[41], SubC_in_s0[41]}), .b ({SubC_in_s3[73], SubC_in_s2[73], SubC_in_s1[73], SubC_in_s0[73]}), .c ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, new_AGEMA_signal_1345, SB_9_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U3 ( .a ({SubC_in_s3[9], SubC_in_s2[9], SubC_in_s1[9], SubC_in_s0[9]}), .b ({SubC_in_s3[105], SubC_in_s2[105], SubC_in_s1[105], SubC_in_s0[105]}), .c ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, new_AGEMA_signal_1354, SB_9_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U8 ( .a ({SubC_in_s3[40], SubC_in_s2[40], SubC_in_s1[40], SubC_in_s0[40]}), .b ({SubC_in_s3[72], SubC_in_s2[72], SubC_in_s1[72], SubC_in_s0[72]}), .c ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, SB_8_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U3 ( .a ({SubC_in_s3[8], SubC_in_s2[8], SubC_in_s1[8], SubC_in_s0[8]}), .b ({SubC_in_s3[104], SubC_in_s2[104], SubC_in_s1[104], SubC_in_s0[104]}), .c ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, new_AGEMA_signal_1384, SB_8_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U8 ( .a ({SubC_in_s3[39], SubC_in_s2[39], SubC_in_s1[39], SubC_in_s0[39]}), .b ({SubC_in_s3[71], SubC_in_s2[71], SubC_in_s1[71], SubC_in_s0[71]}), .c ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, new_AGEMA_signal_1405, SB_7_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U3 ( .a ({SubC_in_s3[7], SubC_in_s2[7], SubC_in_s1[7], SubC_in_s0[7]}), .b ({SubC_in_s3[103], SubC_in_s2[103], SubC_in_s1[103], SubC_in_s0[103]}), .c ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, new_AGEMA_signal_1414, SB_7_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U8 ( .a ({SubC_in_s3[38], SubC_in_s2[38], SubC_in_s1[38], SubC_in_s0[38]}), .b ({SubC_in_s3[70], SubC_in_s2[70], SubC_in_s1[70], SubC_in_s0[70]}), .c ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, new_AGEMA_signal_1435, SB_6_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U3 ( .a ({SubC_in_s3[6], SubC_in_s2[6], SubC_in_s1[6], SubC_in_s0[6]}), .b ({SubC_in_s3[102], SubC_in_s2[102], SubC_in_s1[102], SubC_in_s0[102]}), .c ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, new_AGEMA_signal_1444, SB_6_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U8 ( .a ({SubC_in_s3[37], SubC_in_s2[37], SubC_in_s1[37], SubC_in_s0[37]}), .b ({SubC_in_s3[69], SubC_in_s2[69], SubC_in_s1[69], SubC_in_s0[69]}), .c ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, new_AGEMA_signal_1465, SB_5_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U3 ( .a ({SubC_in_s3[5], SubC_in_s2[5], SubC_in_s1[5], SubC_in_s0[5]}), .b ({SubC_in_s3[101], SubC_in_s2[101], SubC_in_s1[101], SubC_in_s0[101]}), .c ({new_AGEMA_signal_1476, new_AGEMA_signal_1475, new_AGEMA_signal_1474, SB_5_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U8 ( .a ({SubC_in_s3[36], SubC_in_s2[36], SubC_in_s1[36], SubC_in_s0[36]}), .b ({SubC_in_s3[68], SubC_in_s2[68], SubC_in_s1[68], SubC_in_s0[68]}), .c ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, new_AGEMA_signal_1495, SB_4_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U3 ( .a ({SubC_in_s3[4], SubC_in_s2[4], SubC_in_s1[4], SubC_in_s0[4]}), .b ({SubC_in_s3[100], SubC_in_s2[100], SubC_in_s1[100], SubC_in_s0[100]}), .c ({new_AGEMA_signal_1506, new_AGEMA_signal_1505, new_AGEMA_signal_1504, SB_4_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U8 ( .a ({SubC_in_s3[35], SubC_in_s2[35], SubC_in_s1[35], SubC_in_s0[35]}), .b ({SubC_in_s3[67], SubC_in_s2[67], SubC_in_s1[67], SubC_in_s0[67]}), .c ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, SB_3_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U3 ( .a ({SubC_in_s3[3], SubC_in_s2[3], SubC_in_s1[3], SubC_in_s0[3]}), .b ({SubC_in_s3[99], SubC_in_s2[99], SubC_in_s1[99], SubC_in_s0[99]}), .c ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, new_AGEMA_signal_1534, SB_3_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U8 ( .a ({SubC_in_s3[34], SubC_in_s2[34], SubC_in_s1[34], SubC_in_s0[34]}), .b ({SubC_in_s3[66], SubC_in_s2[66], SubC_in_s1[66], SubC_in_s0[66]}), .c ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, new_AGEMA_signal_1555, SB_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U3 ( .a ({SubC_in_s3[2], SubC_in_s2[2], SubC_in_s1[2], SubC_in_s0[2]}), .b ({SubC_in_s3[98], SubC_in_s2[98], SubC_in_s1[98], SubC_in_s0[98]}), .c ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, new_AGEMA_signal_1564, SB_2_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U8 ( .a ({SubC_in_s3[33], SubC_in_s2[33], SubC_in_s1[33], SubC_in_s0[33]}), .b ({SubC_in_s3[65], SubC_in_s2[65], SubC_in_s1[65], SubC_in_s0[65]}), .c ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, new_AGEMA_signal_1585, SB_1_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U3 ( .a ({SubC_in_s3[1], SubC_in_s2[1], SubC_in_s1[1], SubC_in_s0[1]}), .b ({SubC_in_s3[97], SubC_in_s2[97], SubC_in_s1[97], SubC_in_s0[97]}), .c ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, new_AGEMA_signal_1594, SB_1_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U8 ( .a ({SubC_in_s3[32], SubC_in_s2[32], SubC_in_s1[32], SubC_in_s0[32]}), .b ({SubC_in_s3[64], SubC_in_s2[64], SubC_in_s1[64], SubC_in_s0[64]}), .c ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, SB_0_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U3 ( .a ({SubC_in_s3[0], SubC_in_s2[0], SubC_in_s1[0], SubC_in_s0[0]}), .b ({SubC_in_s3[96], SubC_in_s2[96], SubC_in_s1[96], SubC_in_s0[96]}), .c ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, new_AGEMA_signal_1624, SB_0_n10}) ) ;
    //ClockGatingController #(4) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U11 ( .a ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, SB_31_n15}), .b ({new_AGEMA_signal_687, new_AGEMA_signal_686, new_AGEMA_signal_685, SB_31_n14}), .c ({SubC_out_s3[127], SubC_out_s2[127], SubC_out_s1[127], SubC_out_s0[127]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U9 ( .a ({new_AGEMA_signal_687, new_AGEMA_signal_686, new_AGEMA_signal_685, SB_31_n14}), .b ({new_AGEMA_signal_705, new_AGEMA_signal_704, new_AGEMA_signal_703, SB_31_T2}), .c ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, new_AGEMA_signal_1639, SB_31_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U6 ( .a ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, new_AGEMA_signal_2125, SB_31_n11}), .b ({new_AGEMA_signal_702, new_AGEMA_signal_701, new_AGEMA_signal_700, SB_31_T1}), .c ({SubC_out_s3[95], SubC_out_s2[95], SubC_out_s1[95], SubC_out_s0[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U5 ( .a ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, SB_31_n15}), .b ({SubC_in_s3[63], SubC_in_s2[63], SubC_in_s1[63], SubC_in_s0[63]}), .c ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, new_AGEMA_signal_2125, SB_31_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U4 ( .a ({new_AGEMA_signal_696, new_AGEMA_signal_695, new_AGEMA_signal_694, SB_31_n10}), .b ({new_AGEMA_signal_699, new_AGEMA_signal_698, new_AGEMA_signal_697, SB_31_T0}), .c ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, new_AGEMA_signal_1642, SB_31_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U1 ( .a ({SubC_in_s3[127], SubC_in_s2[127], SubC_in_s1[127], SubC_in_s0[127]}), .b ({new_AGEMA_signal_708, new_AGEMA_signal_707, new_AGEMA_signal_706, SB_31_T3}), .c ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, new_AGEMA_signal_1645, SB_31_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_31_t0_AND_U1 ( .a ({SubC_in_s3[127], SubC_in_s2[127], SubC_in_s1[127], SubC_in_s0[127]}), .b ({SubC_in_s3[95], SubC_in_s2[95], SubC_in_s1[95], SubC_in_s0[95]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_699, new_AGEMA_signal_698, new_AGEMA_signal_697, SB_31_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_31_t1_AND_U1 ( .a ({SubC_in_s3[127], SubC_in_s2[127], SubC_in_s1[127], SubC_in_s0[127]}), .b ({SubC_in_s3[63], SubC_in_s2[63], SubC_in_s1[63], SubC_in_s0[63]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_702, new_AGEMA_signal_701, new_AGEMA_signal_700, SB_31_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_31_t2_AND_U1 ( .a ({SubC_in_s3[127], SubC_in_s2[127], SubC_in_s1[127], SubC_in_s0[127]}), .b ({SubC_in_s3[31], SubC_in_s2[31], SubC_in_s1[31], SubC_in_s0[31]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_705, new_AGEMA_signal_704, new_AGEMA_signal_703, SB_31_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_31_t3_AND_U1 ( .a ({SubC_in_s3[95], SubC_in_s2[95], SubC_in_s1[95], SubC_in_s0[95]}), .b ({SubC_in_s3[31], SubC_in_s2[31], SubC_in_s1[31], SubC_in_s0[31]}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_708, new_AGEMA_signal_707, new_AGEMA_signal_706, SB_31_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U11 ( .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, new_AGEMA_signal_1657, SB_30_n15}), .b ({new_AGEMA_signal_717, new_AGEMA_signal_716, new_AGEMA_signal_715, SB_30_n14}), .c ({SubC_out_s3[126], SubC_out_s2[126], SubC_out_s1[126], SubC_out_s0[126]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U9 ( .a ({new_AGEMA_signal_717, new_AGEMA_signal_716, new_AGEMA_signal_715, SB_30_n14}), .b ({new_AGEMA_signal_735, new_AGEMA_signal_734, new_AGEMA_signal_733, SB_30_T2}), .c ({new_AGEMA_signal_1656, new_AGEMA_signal_1655, new_AGEMA_signal_1654, SB_30_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U6 ( .a ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, SB_30_n11}), .b ({new_AGEMA_signal_732, new_AGEMA_signal_731, new_AGEMA_signal_730, SB_30_T1}), .c ({SubC_out_s3[94], SubC_out_s2[94], SubC_out_s1[94], SubC_out_s0[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U5 ( .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, new_AGEMA_signal_1657, SB_30_n15}), .b ({SubC_in_s3[62], SubC_in_s2[62], SubC_in_s1[62], SubC_in_s0[62]}), .c ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, SB_30_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U4 ( .a ({new_AGEMA_signal_726, new_AGEMA_signal_725, new_AGEMA_signal_724, SB_30_n10}), .b ({new_AGEMA_signal_729, new_AGEMA_signal_728, new_AGEMA_signal_727, SB_30_T0}), .c ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, new_AGEMA_signal_1657, SB_30_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U1 ( .a ({SubC_in_s3[126], SubC_in_s2[126], SubC_in_s1[126], SubC_in_s0[126]}), .b ({new_AGEMA_signal_738, new_AGEMA_signal_737, new_AGEMA_signal_736, SB_30_T3}), .c ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, SB_30_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_30_t0_AND_U1 ( .a ({SubC_in_s3[126], SubC_in_s2[126], SubC_in_s1[126], SubC_in_s0[126]}), .b ({SubC_in_s3[94], SubC_in_s2[94], SubC_in_s1[94], SubC_in_s0[94]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_729, new_AGEMA_signal_728, new_AGEMA_signal_727, SB_30_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_30_t1_AND_U1 ( .a ({SubC_in_s3[126], SubC_in_s2[126], SubC_in_s1[126], SubC_in_s0[126]}), .b ({SubC_in_s3[62], SubC_in_s2[62], SubC_in_s1[62], SubC_in_s0[62]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_732, new_AGEMA_signal_731, new_AGEMA_signal_730, SB_30_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_30_t2_AND_U1 ( .a ({SubC_in_s3[126], SubC_in_s2[126], SubC_in_s1[126], SubC_in_s0[126]}), .b ({SubC_in_s3[30], SubC_in_s2[30], SubC_in_s1[30], SubC_in_s0[30]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_735, new_AGEMA_signal_734, new_AGEMA_signal_733, SB_30_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_30_t3_AND_U1 ( .a ({SubC_in_s3[94], SubC_in_s2[94], SubC_in_s1[94], SubC_in_s0[94]}), .b ({SubC_in_s3[30], SubC_in_s2[30], SubC_in_s1[30], SubC_in_s0[30]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_738, new_AGEMA_signal_737, new_AGEMA_signal_736, SB_30_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U11 ( .a ({new_AGEMA_signal_1674, new_AGEMA_signal_1673, new_AGEMA_signal_1672, SB_29_n15}), .b ({new_AGEMA_signal_747, new_AGEMA_signal_746, new_AGEMA_signal_745, SB_29_n14}), .c ({SubC_out_s3[125], SubC_out_s2[125], SubC_out_s1[125], SubC_out_s0[125]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U9 ( .a ({new_AGEMA_signal_747, new_AGEMA_signal_746, new_AGEMA_signal_745, SB_29_n14}), .b ({new_AGEMA_signal_765, new_AGEMA_signal_764, new_AGEMA_signal_763, SB_29_T2}), .c ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, new_AGEMA_signal_1669, SB_29_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U6 ( .a ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, new_AGEMA_signal_2149, SB_29_n11}), .b ({new_AGEMA_signal_762, new_AGEMA_signal_761, new_AGEMA_signal_760, SB_29_T1}), .c ({SubC_out_s3[93], SubC_out_s2[93], SubC_out_s1[93], SubC_out_s0[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U5 ( .a ({new_AGEMA_signal_1674, new_AGEMA_signal_1673, new_AGEMA_signal_1672, SB_29_n15}), .b ({SubC_in_s3[61], SubC_in_s2[61], SubC_in_s1[61], SubC_in_s0[61]}), .c ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, new_AGEMA_signal_2149, SB_29_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U4 ( .a ({new_AGEMA_signal_756, new_AGEMA_signal_755, new_AGEMA_signal_754, SB_29_n10}), .b ({new_AGEMA_signal_759, new_AGEMA_signal_758, new_AGEMA_signal_757, SB_29_T0}), .c ({new_AGEMA_signal_1674, new_AGEMA_signal_1673, new_AGEMA_signal_1672, SB_29_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U1 ( .a ({SubC_in_s3[125], SubC_in_s2[125], SubC_in_s1[125], SubC_in_s0[125]}), .b ({new_AGEMA_signal_768, new_AGEMA_signal_767, new_AGEMA_signal_766, SB_29_T3}), .c ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, new_AGEMA_signal_1675, SB_29_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_29_t0_AND_U1 ( .a ({SubC_in_s3[125], SubC_in_s2[125], SubC_in_s1[125], SubC_in_s0[125]}), .b ({SubC_in_s3[93], SubC_in_s2[93], SubC_in_s1[93], SubC_in_s0[93]}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_759, new_AGEMA_signal_758, new_AGEMA_signal_757, SB_29_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_29_t1_AND_U1 ( .a ({SubC_in_s3[125], SubC_in_s2[125], SubC_in_s1[125], SubC_in_s0[125]}), .b ({SubC_in_s3[61], SubC_in_s2[61], SubC_in_s1[61], SubC_in_s0[61]}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_762, new_AGEMA_signal_761, new_AGEMA_signal_760, SB_29_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_29_t2_AND_U1 ( .a ({SubC_in_s3[125], SubC_in_s2[125], SubC_in_s1[125], SubC_in_s0[125]}), .b ({SubC_in_s3[29], SubC_in_s2[29], SubC_in_s1[29], SubC_in_s0[29]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_765, new_AGEMA_signal_764, new_AGEMA_signal_763, SB_29_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_29_t3_AND_U1 ( .a ({SubC_in_s3[93], SubC_in_s2[93], SubC_in_s1[93], SubC_in_s0[93]}), .b ({SubC_in_s3[29], SubC_in_s2[29], SubC_in_s1[29], SubC_in_s0[29]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_768, new_AGEMA_signal_767, new_AGEMA_signal_766, SB_29_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U11 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, SB_28_n15}), .b ({new_AGEMA_signal_777, new_AGEMA_signal_776, new_AGEMA_signal_775, SB_28_n14}), .c ({SubC_out_s3[124], SubC_out_s2[124], SubC_out_s1[124], SubC_out_s0[124]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U9 ( .a ({new_AGEMA_signal_777, new_AGEMA_signal_776, new_AGEMA_signal_775, SB_28_n14}), .b ({new_AGEMA_signal_795, new_AGEMA_signal_794, new_AGEMA_signal_793, SB_28_T2}), .c ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, new_AGEMA_signal_1684, SB_28_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U6 ( .a ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, new_AGEMA_signal_2161, SB_28_n11}), .b ({new_AGEMA_signal_792, new_AGEMA_signal_791, new_AGEMA_signal_790, SB_28_T1}), .c ({SubC_out_s3[92], SubC_out_s2[92], SubC_out_s1[92], SubC_out_s0[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U5 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, SB_28_n15}), .b ({SubC_in_s3[60], SubC_in_s2[60], SubC_in_s1[60], SubC_in_s0[60]}), .c ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, new_AGEMA_signal_2161, SB_28_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U4 ( .a ({new_AGEMA_signal_786, new_AGEMA_signal_785, new_AGEMA_signal_784, SB_28_n10}), .b ({new_AGEMA_signal_789, new_AGEMA_signal_788, new_AGEMA_signal_787, SB_28_T0}), .c ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, SB_28_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U1 ( .a ({SubC_in_s3[124], SubC_in_s2[124], SubC_in_s1[124], SubC_in_s0[124]}), .b ({new_AGEMA_signal_798, new_AGEMA_signal_797, new_AGEMA_signal_796, SB_28_T3}), .c ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, new_AGEMA_signal_1690, SB_28_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_28_t0_AND_U1 ( .a ({SubC_in_s3[124], SubC_in_s2[124], SubC_in_s1[124], SubC_in_s0[124]}), .b ({SubC_in_s3[92], SubC_in_s2[92], SubC_in_s1[92], SubC_in_s0[92]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_789, new_AGEMA_signal_788, new_AGEMA_signal_787, SB_28_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_28_t1_AND_U1 ( .a ({SubC_in_s3[124], SubC_in_s2[124], SubC_in_s1[124], SubC_in_s0[124]}), .b ({SubC_in_s3[60], SubC_in_s2[60], SubC_in_s1[60], SubC_in_s0[60]}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_792, new_AGEMA_signal_791, new_AGEMA_signal_790, SB_28_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_28_t2_AND_U1 ( .a ({SubC_in_s3[124], SubC_in_s2[124], SubC_in_s1[124], SubC_in_s0[124]}), .b ({SubC_in_s3[28], SubC_in_s2[28], SubC_in_s1[28], SubC_in_s0[28]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_795, new_AGEMA_signal_794, new_AGEMA_signal_793, SB_28_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_28_t3_AND_U1 ( .a ({SubC_in_s3[92], SubC_in_s2[92], SubC_in_s1[92], SubC_in_s0[92]}), .b ({SubC_in_s3[28], SubC_in_s2[28], SubC_in_s1[28], SubC_in_s0[28]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_798, new_AGEMA_signal_797, new_AGEMA_signal_796, SB_28_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U11 ( .a ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, new_AGEMA_signal_1702, SB_27_n15}), .b ({new_AGEMA_signal_807, new_AGEMA_signal_806, new_AGEMA_signal_805, SB_27_n14}), .c ({SubC_out_s3[123], SubC_out_s2[123], SubC_out_s1[123], SubC_out_s0[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U9 ( .a ({new_AGEMA_signal_807, new_AGEMA_signal_806, new_AGEMA_signal_805, SB_27_n14}), .b ({new_AGEMA_signal_825, new_AGEMA_signal_824, new_AGEMA_signal_823, SB_27_T2}), .c ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, new_AGEMA_signal_1699, SB_27_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U6 ( .a ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, new_AGEMA_signal_2173, SB_27_n11}), .b ({new_AGEMA_signal_822, new_AGEMA_signal_821, new_AGEMA_signal_820, SB_27_T1}), .c ({SubC_out_s3[91], SubC_out_s2[91], SubC_out_s1[91], SubC_out_s0[91]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U5 ( .a ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, new_AGEMA_signal_1702, SB_27_n15}), .b ({SubC_in_s3[59], SubC_in_s2[59], SubC_in_s1[59], SubC_in_s0[59]}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, new_AGEMA_signal_2173, SB_27_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U4 ( .a ({new_AGEMA_signal_816, new_AGEMA_signal_815, new_AGEMA_signal_814, SB_27_n10}), .b ({new_AGEMA_signal_819, new_AGEMA_signal_818, new_AGEMA_signal_817, SB_27_T0}), .c ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, new_AGEMA_signal_1702, SB_27_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U1 ( .a ({SubC_in_s3[123], SubC_in_s2[123], SubC_in_s1[123], SubC_in_s0[123]}), .b ({new_AGEMA_signal_828, new_AGEMA_signal_827, new_AGEMA_signal_826, SB_27_T3}), .c ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, new_AGEMA_signal_1705, SB_27_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_27_t0_AND_U1 ( .a ({SubC_in_s3[123], SubC_in_s2[123], SubC_in_s1[123], SubC_in_s0[123]}), .b ({SubC_in_s3[91], SubC_in_s2[91], SubC_in_s1[91], SubC_in_s0[91]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_819, new_AGEMA_signal_818, new_AGEMA_signal_817, SB_27_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_27_t1_AND_U1 ( .a ({SubC_in_s3[123], SubC_in_s2[123], SubC_in_s1[123], SubC_in_s0[123]}), .b ({SubC_in_s3[59], SubC_in_s2[59], SubC_in_s1[59], SubC_in_s0[59]}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_822, new_AGEMA_signal_821, new_AGEMA_signal_820, SB_27_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_27_t2_AND_U1 ( .a ({SubC_in_s3[123], SubC_in_s2[123], SubC_in_s1[123], SubC_in_s0[123]}), .b ({SubC_in_s3[27], SubC_in_s2[27], SubC_in_s1[27], SubC_in_s0[27]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_825, new_AGEMA_signal_824, new_AGEMA_signal_823, SB_27_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_27_t3_AND_U1 ( .a ({SubC_in_s3[91], SubC_in_s2[91], SubC_in_s1[91], SubC_in_s0[91]}), .b ({SubC_in_s3[27], SubC_in_s2[27], SubC_in_s1[27], SubC_in_s0[27]}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_828, new_AGEMA_signal_827, new_AGEMA_signal_826, SB_27_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U11 ( .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, new_AGEMA_signal_1717, SB_26_n15}), .b ({new_AGEMA_signal_837, new_AGEMA_signal_836, new_AGEMA_signal_835, SB_26_n14}), .c ({SubC_out_s3[122], SubC_out_s2[122], SubC_out_s1[122], SubC_out_s0[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U9 ( .a ({new_AGEMA_signal_837, new_AGEMA_signal_836, new_AGEMA_signal_835, SB_26_n14}), .b ({new_AGEMA_signal_855, new_AGEMA_signal_854, new_AGEMA_signal_853, SB_26_T2}), .c ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, SB_26_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U6 ( .a ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, new_AGEMA_signal_2185, SB_26_n11}), .b ({new_AGEMA_signal_852, new_AGEMA_signal_851, new_AGEMA_signal_850, SB_26_T1}), .c ({SubC_out_s3[90], SubC_out_s2[90], SubC_out_s1[90], SubC_out_s0[90]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U5 ( .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, new_AGEMA_signal_1717, SB_26_n15}), .b ({SubC_in_s3[58], SubC_in_s2[58], SubC_in_s1[58], SubC_in_s0[58]}), .c ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, new_AGEMA_signal_2185, SB_26_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U4 ( .a ({new_AGEMA_signal_846, new_AGEMA_signal_845, new_AGEMA_signal_844, SB_26_n10}), .b ({new_AGEMA_signal_849, new_AGEMA_signal_848, new_AGEMA_signal_847, SB_26_T0}), .c ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, new_AGEMA_signal_1717, SB_26_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U1 ( .a ({SubC_in_s3[122], SubC_in_s2[122], SubC_in_s1[122], SubC_in_s0[122]}), .b ({new_AGEMA_signal_858, new_AGEMA_signal_857, new_AGEMA_signal_856, SB_26_T3}), .c ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, new_AGEMA_signal_1720, SB_26_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_26_t0_AND_U1 ( .a ({SubC_in_s3[122], SubC_in_s2[122], SubC_in_s1[122], SubC_in_s0[122]}), .b ({SubC_in_s3[90], SubC_in_s2[90], SubC_in_s1[90], SubC_in_s0[90]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_849, new_AGEMA_signal_848, new_AGEMA_signal_847, SB_26_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_26_t1_AND_U1 ( .a ({SubC_in_s3[122], SubC_in_s2[122], SubC_in_s1[122], SubC_in_s0[122]}), .b ({SubC_in_s3[58], SubC_in_s2[58], SubC_in_s1[58], SubC_in_s0[58]}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_852, new_AGEMA_signal_851, new_AGEMA_signal_850, SB_26_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_26_t2_AND_U1 ( .a ({SubC_in_s3[122], SubC_in_s2[122], SubC_in_s1[122], SubC_in_s0[122]}), .b ({SubC_in_s3[26], SubC_in_s2[26], SubC_in_s1[26], SubC_in_s0[26]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_855, new_AGEMA_signal_854, new_AGEMA_signal_853, SB_26_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_26_t3_AND_U1 ( .a ({SubC_in_s3[90], SubC_in_s2[90], SubC_in_s1[90], SubC_in_s0[90]}), .b ({SubC_in_s3[26], SubC_in_s2[26], SubC_in_s1[26], SubC_in_s0[26]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_858, new_AGEMA_signal_857, new_AGEMA_signal_856, SB_26_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U11 ( .a ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, new_AGEMA_signal_1732, SB_25_n15}), .b ({new_AGEMA_signal_867, new_AGEMA_signal_866, new_AGEMA_signal_865, SB_25_n14}), .c ({SubC_out_s3[121], SubC_out_s2[121], SubC_out_s1[121], SubC_out_s0[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U9 ( .a ({new_AGEMA_signal_867, new_AGEMA_signal_866, new_AGEMA_signal_865, SB_25_n14}), .b ({new_AGEMA_signal_885, new_AGEMA_signal_884, new_AGEMA_signal_883, SB_25_T2}), .c ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, new_AGEMA_signal_1729, SB_25_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U6 ( .a ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, new_AGEMA_signal_2197, SB_25_n11}), .b ({new_AGEMA_signal_882, new_AGEMA_signal_881, new_AGEMA_signal_880, SB_25_T1}), .c ({SubC_out_s3[89], SubC_out_s2[89], SubC_out_s1[89], SubC_out_s0[89]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U5 ( .a ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, new_AGEMA_signal_1732, SB_25_n15}), .b ({SubC_in_s3[57], SubC_in_s2[57], SubC_in_s1[57], SubC_in_s0[57]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, new_AGEMA_signal_2197, SB_25_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U4 ( .a ({new_AGEMA_signal_876, new_AGEMA_signal_875, new_AGEMA_signal_874, SB_25_n10}), .b ({new_AGEMA_signal_879, new_AGEMA_signal_878, new_AGEMA_signal_877, SB_25_T0}), .c ({new_AGEMA_signal_1734, new_AGEMA_signal_1733, new_AGEMA_signal_1732, SB_25_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U1 ( .a ({SubC_in_s3[121], SubC_in_s2[121], SubC_in_s1[121], SubC_in_s0[121]}), .b ({new_AGEMA_signal_888, new_AGEMA_signal_887, new_AGEMA_signal_886, SB_25_T3}), .c ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, new_AGEMA_signal_1735, SB_25_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_25_t0_AND_U1 ( .a ({SubC_in_s3[121], SubC_in_s2[121], SubC_in_s1[121], SubC_in_s0[121]}), .b ({SubC_in_s3[89], SubC_in_s2[89], SubC_in_s1[89], SubC_in_s0[89]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_879, new_AGEMA_signal_878, new_AGEMA_signal_877, SB_25_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_25_t1_AND_U1 ( .a ({SubC_in_s3[121], SubC_in_s2[121], SubC_in_s1[121], SubC_in_s0[121]}), .b ({SubC_in_s3[57], SubC_in_s2[57], SubC_in_s1[57], SubC_in_s0[57]}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_882, new_AGEMA_signal_881, new_AGEMA_signal_880, SB_25_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_25_t2_AND_U1 ( .a ({SubC_in_s3[121], SubC_in_s2[121], SubC_in_s1[121], SubC_in_s0[121]}), .b ({SubC_in_s3[25], SubC_in_s2[25], SubC_in_s1[25], SubC_in_s0[25]}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_885, new_AGEMA_signal_884, new_AGEMA_signal_883, SB_25_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_25_t3_AND_U1 ( .a ({SubC_in_s3[89], SubC_in_s2[89], SubC_in_s1[89], SubC_in_s0[89]}), .b ({SubC_in_s3[25], SubC_in_s2[25], SubC_in_s1[25], SubC_in_s0[25]}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_888, new_AGEMA_signal_887, new_AGEMA_signal_886, SB_25_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U11 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, SB_24_n15}), .b ({new_AGEMA_signal_897, new_AGEMA_signal_896, new_AGEMA_signal_895, SB_24_n14}), .c ({SubC_out_s3[120], SubC_out_s2[120], SubC_out_s1[120], SubC_out_s0[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U9 ( .a ({new_AGEMA_signal_897, new_AGEMA_signal_896, new_AGEMA_signal_895, SB_24_n14}), .b ({new_AGEMA_signal_915, new_AGEMA_signal_914, new_AGEMA_signal_913, SB_24_T2}), .c ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, new_AGEMA_signal_1744, SB_24_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U6 ( .a ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, new_AGEMA_signal_2209, SB_24_n11}), .b ({new_AGEMA_signal_912, new_AGEMA_signal_911, new_AGEMA_signal_910, SB_24_T1}), .c ({SubC_out_s3[88], SubC_out_s2[88], SubC_out_s1[88], SubC_out_s0[88]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U5 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, SB_24_n15}), .b ({SubC_in_s3[56], SubC_in_s2[56], SubC_in_s1[56], SubC_in_s0[56]}), .c ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, new_AGEMA_signal_2209, SB_24_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U4 ( .a ({new_AGEMA_signal_906, new_AGEMA_signal_905, new_AGEMA_signal_904, SB_24_n10}), .b ({new_AGEMA_signal_909, new_AGEMA_signal_908, new_AGEMA_signal_907, SB_24_T0}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, SB_24_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U1 ( .a ({SubC_in_s3[120], SubC_in_s2[120], SubC_in_s1[120], SubC_in_s0[120]}), .b ({new_AGEMA_signal_918, new_AGEMA_signal_917, new_AGEMA_signal_916, SB_24_T3}), .c ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, SB_24_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_24_t0_AND_U1 ( .a ({SubC_in_s3[120], SubC_in_s2[120], SubC_in_s1[120], SubC_in_s0[120]}), .b ({SubC_in_s3[88], SubC_in_s2[88], SubC_in_s1[88], SubC_in_s0[88]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_909, new_AGEMA_signal_908, new_AGEMA_signal_907, SB_24_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_24_t1_AND_U1 ( .a ({SubC_in_s3[120], SubC_in_s2[120], SubC_in_s1[120], SubC_in_s0[120]}), .b ({SubC_in_s3[56], SubC_in_s2[56], SubC_in_s1[56], SubC_in_s0[56]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_912, new_AGEMA_signal_911, new_AGEMA_signal_910, SB_24_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_24_t2_AND_U1 ( .a ({SubC_in_s3[120], SubC_in_s2[120], SubC_in_s1[120], SubC_in_s0[120]}), .b ({SubC_in_s3[24], SubC_in_s2[24], SubC_in_s1[24], SubC_in_s0[24]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_915, new_AGEMA_signal_914, new_AGEMA_signal_913, SB_24_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_24_t3_AND_U1 ( .a ({SubC_in_s3[88], SubC_in_s2[88], SubC_in_s1[88], SubC_in_s0[88]}), .b ({SubC_in_s3[24], SubC_in_s2[24], SubC_in_s1[24], SubC_in_s0[24]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_918, new_AGEMA_signal_917, new_AGEMA_signal_916, SB_24_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U11 ( .a ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, new_AGEMA_signal_1762, SB_23_n15}), .b ({new_AGEMA_signal_927, new_AGEMA_signal_926, new_AGEMA_signal_925, SB_23_n14}), .c ({SubC_out_s3[119], SubC_out_s2[119], SubC_out_s1[119], SubC_out_s0[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U9 ( .a ({new_AGEMA_signal_927, new_AGEMA_signal_926, new_AGEMA_signal_925, SB_23_n14}), .b ({new_AGEMA_signal_945, new_AGEMA_signal_944, new_AGEMA_signal_943, SB_23_T2}), .c ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, SB_23_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U6 ( .a ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, new_AGEMA_signal_2221, SB_23_n11}), .b ({new_AGEMA_signal_942, new_AGEMA_signal_941, new_AGEMA_signal_940, SB_23_T1}), .c ({SubC_out_s3[87], SubC_out_s2[87], SubC_out_s1[87], SubC_out_s0[87]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U5 ( .a ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, new_AGEMA_signal_1762, SB_23_n15}), .b ({SubC_in_s3[55], SubC_in_s2[55], SubC_in_s1[55], SubC_in_s0[55]}), .c ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, new_AGEMA_signal_2221, SB_23_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U4 ( .a ({new_AGEMA_signal_936, new_AGEMA_signal_935, new_AGEMA_signal_934, SB_23_n10}), .b ({new_AGEMA_signal_939, new_AGEMA_signal_938, new_AGEMA_signal_937, SB_23_T0}), .c ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, new_AGEMA_signal_1762, SB_23_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U1 ( .a ({SubC_in_s3[119], SubC_in_s2[119], SubC_in_s1[119], SubC_in_s0[119]}), .b ({new_AGEMA_signal_948, new_AGEMA_signal_947, new_AGEMA_signal_946, SB_23_T3}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, new_AGEMA_signal_1765, SB_23_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_23_t0_AND_U1 ( .a ({SubC_in_s3[119], SubC_in_s2[119], SubC_in_s1[119], SubC_in_s0[119]}), .b ({SubC_in_s3[87], SubC_in_s2[87], SubC_in_s1[87], SubC_in_s0[87]}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_939, new_AGEMA_signal_938, new_AGEMA_signal_937, SB_23_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_23_t1_AND_U1 ( .a ({SubC_in_s3[119], SubC_in_s2[119], SubC_in_s1[119], SubC_in_s0[119]}), .b ({SubC_in_s3[55], SubC_in_s2[55], SubC_in_s1[55], SubC_in_s0[55]}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_942, new_AGEMA_signal_941, new_AGEMA_signal_940, SB_23_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_23_t2_AND_U1 ( .a ({SubC_in_s3[119], SubC_in_s2[119], SubC_in_s1[119], SubC_in_s0[119]}), .b ({SubC_in_s3[23], SubC_in_s2[23], SubC_in_s1[23], SubC_in_s0[23]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_945, new_AGEMA_signal_944, new_AGEMA_signal_943, SB_23_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_23_t3_AND_U1 ( .a ({SubC_in_s3[87], SubC_in_s2[87], SubC_in_s1[87], SubC_in_s0[87]}), .b ({SubC_in_s3[23], SubC_in_s2[23], SubC_in_s1[23], SubC_in_s0[23]}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_948, new_AGEMA_signal_947, new_AGEMA_signal_946, SB_23_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U11 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, SB_22_n15}), .b ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, SB_22_n14}), .c ({SubC_out_s3[118], SubC_out_s2[118], SubC_out_s1[118], SubC_out_s0[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U9 ( .a ({new_AGEMA_signal_957, new_AGEMA_signal_956, new_AGEMA_signal_955, SB_22_n14}), .b ({new_AGEMA_signal_975, new_AGEMA_signal_974, new_AGEMA_signal_973, SB_22_T2}), .c ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, new_AGEMA_signal_1774, SB_22_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U6 ( .a ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, SB_22_n11}), .b ({new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, SB_22_T1}), .c ({SubC_out_s3[86], SubC_out_s2[86], SubC_out_s1[86], SubC_out_s0[86]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U5 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, SB_22_n15}), .b ({SubC_in_s3[54], SubC_in_s2[54], SubC_in_s1[54], SubC_in_s0[54]}), .c ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, SB_22_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U4 ( .a ({new_AGEMA_signal_966, new_AGEMA_signal_965, new_AGEMA_signal_964, SB_22_n10}), .b ({new_AGEMA_signal_969, new_AGEMA_signal_968, new_AGEMA_signal_967, SB_22_T0}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, SB_22_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U1 ( .a ({SubC_in_s3[118], SubC_in_s2[118], SubC_in_s1[118], SubC_in_s0[118]}), .b ({new_AGEMA_signal_978, new_AGEMA_signal_977, new_AGEMA_signal_976, SB_22_T3}), .c ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, new_AGEMA_signal_1780, SB_22_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_22_t0_AND_U1 ( .a ({SubC_in_s3[118], SubC_in_s2[118], SubC_in_s1[118], SubC_in_s0[118]}), .b ({SubC_in_s3[86], SubC_in_s2[86], SubC_in_s1[86], SubC_in_s0[86]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_969, new_AGEMA_signal_968, new_AGEMA_signal_967, SB_22_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_22_t1_AND_U1 ( .a ({SubC_in_s3[118], SubC_in_s2[118], SubC_in_s1[118], SubC_in_s0[118]}), .b ({SubC_in_s3[54], SubC_in_s2[54], SubC_in_s1[54], SubC_in_s0[54]}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_972, new_AGEMA_signal_971, new_AGEMA_signal_970, SB_22_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_22_t2_AND_U1 ( .a ({SubC_in_s3[118], SubC_in_s2[118], SubC_in_s1[118], SubC_in_s0[118]}), .b ({SubC_in_s3[22], SubC_in_s2[22], SubC_in_s1[22], SubC_in_s0[22]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_975, new_AGEMA_signal_974, new_AGEMA_signal_973, SB_22_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_22_t3_AND_U1 ( .a ({SubC_in_s3[86], SubC_in_s2[86], SubC_in_s1[86], SubC_in_s0[86]}), .b ({SubC_in_s3[22], SubC_in_s2[22], SubC_in_s1[22], SubC_in_s0[22]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_978, new_AGEMA_signal_977, new_AGEMA_signal_976, SB_22_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U11 ( .a ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, new_AGEMA_signal_1792, SB_21_n15}), .b ({new_AGEMA_signal_987, new_AGEMA_signal_986, new_AGEMA_signal_985, SB_21_n14}), .c ({SubC_out_s3[117], SubC_out_s2[117], SubC_out_s1[117], SubC_out_s0[117]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U9 ( .a ({new_AGEMA_signal_987, new_AGEMA_signal_986, new_AGEMA_signal_985, SB_21_n14}), .b ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, SB_21_T2}), .c ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, new_AGEMA_signal_1789, SB_21_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U6 ( .a ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, new_AGEMA_signal_2245, SB_21_n11}), .b ({new_AGEMA_signal_1002, new_AGEMA_signal_1001, new_AGEMA_signal_1000, SB_21_T1}), .c ({SubC_out_s3[85], SubC_out_s2[85], SubC_out_s1[85], SubC_out_s0[85]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U5 ( .a ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, new_AGEMA_signal_1792, SB_21_n15}), .b ({SubC_in_s3[53], SubC_in_s2[53], SubC_in_s1[53], SubC_in_s0[53]}), .c ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, new_AGEMA_signal_2245, SB_21_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U4 ( .a ({new_AGEMA_signal_996, new_AGEMA_signal_995, new_AGEMA_signal_994, SB_21_n10}), .b ({new_AGEMA_signal_999, new_AGEMA_signal_998, new_AGEMA_signal_997, SB_21_T0}), .c ({new_AGEMA_signal_1794, new_AGEMA_signal_1793, new_AGEMA_signal_1792, SB_21_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U1 ( .a ({SubC_in_s3[117], SubC_in_s2[117], SubC_in_s1[117], SubC_in_s0[117]}), .b ({new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, SB_21_T3}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, SB_21_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_21_t0_AND_U1 ( .a ({SubC_in_s3[117], SubC_in_s2[117], SubC_in_s1[117], SubC_in_s0[117]}), .b ({SubC_in_s3[85], SubC_in_s2[85], SubC_in_s1[85], SubC_in_s0[85]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_999, new_AGEMA_signal_998, new_AGEMA_signal_997, SB_21_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_21_t1_AND_U1 ( .a ({SubC_in_s3[117], SubC_in_s2[117], SubC_in_s1[117], SubC_in_s0[117]}), .b ({SubC_in_s3[53], SubC_in_s2[53], SubC_in_s1[53], SubC_in_s0[53]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1002, new_AGEMA_signal_1001, new_AGEMA_signal_1000, SB_21_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_21_t2_AND_U1 ( .a ({SubC_in_s3[117], SubC_in_s2[117], SubC_in_s1[117], SubC_in_s0[117]}), .b ({SubC_in_s3[21], SubC_in_s2[21], SubC_in_s1[21], SubC_in_s0[21]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, SB_21_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_21_t3_AND_U1 ( .a ({SubC_in_s3[85], SubC_in_s2[85], SubC_in_s1[85], SubC_in_s0[85]}), .b ({SubC_in_s3[21], SubC_in_s2[21], SubC_in_s1[21], SubC_in_s0[21]}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, SB_21_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U11 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, new_AGEMA_signal_1807, SB_20_n15}), .b ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, SB_20_n14}), .c ({SubC_out_s3[116], SubC_out_s2[116], SubC_out_s1[116], SubC_out_s0[116]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U9 ( .a ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, new_AGEMA_signal_1015, SB_20_n14}), .b ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, new_AGEMA_signal_1033, SB_20_T2}), .c ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, new_AGEMA_signal_1804, SB_20_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U6 ( .a ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, new_AGEMA_signal_2257, SB_20_n11}), .b ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, SB_20_T1}), .c ({SubC_out_s3[84], SubC_out_s2[84], SubC_out_s1[84], SubC_out_s0[84]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U5 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, new_AGEMA_signal_1807, SB_20_n15}), .b ({SubC_in_s3[52], SubC_in_s2[52], SubC_in_s1[52], SubC_in_s0[52]}), .c ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, new_AGEMA_signal_2257, SB_20_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U4 ( .a ({new_AGEMA_signal_1026, new_AGEMA_signal_1025, new_AGEMA_signal_1024, SB_20_n10}), .b ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, new_AGEMA_signal_1027, SB_20_T0}), .c ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, new_AGEMA_signal_1807, SB_20_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U1 ( .a ({SubC_in_s3[116], SubC_in_s2[116], SubC_in_s1[116], SubC_in_s0[116]}), .b ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, new_AGEMA_signal_1036, SB_20_T3}), .c ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, new_AGEMA_signal_1810, SB_20_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_20_t0_AND_U1 ( .a ({SubC_in_s3[116], SubC_in_s2[116], SubC_in_s1[116], SubC_in_s0[116]}), .b ({SubC_in_s3[84], SubC_in_s2[84], SubC_in_s1[84], SubC_in_s0[84]}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, new_AGEMA_signal_1027, SB_20_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_20_t1_AND_U1 ( .a ({SubC_in_s3[116], SubC_in_s2[116], SubC_in_s1[116], SubC_in_s0[116]}), .b ({SubC_in_s3[52], SubC_in_s2[52], SubC_in_s1[52], SubC_in_s0[52]}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1032, new_AGEMA_signal_1031, new_AGEMA_signal_1030, SB_20_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_20_t2_AND_U1 ( .a ({SubC_in_s3[116], SubC_in_s2[116], SubC_in_s1[116], SubC_in_s0[116]}), .b ({SubC_in_s3[20], SubC_in_s2[20], SubC_in_s1[20], SubC_in_s0[20]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, new_AGEMA_signal_1033, SB_20_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_20_t3_AND_U1 ( .a ({SubC_in_s3[84], SubC_in_s2[84], SubC_in_s1[84], SubC_in_s0[84]}), .b ({SubC_in_s3[20], SubC_in_s2[20], SubC_in_s1[20], SubC_in_s0[20]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, new_AGEMA_signal_1036, SB_20_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U11 ( .a ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, new_AGEMA_signal_1822, SB_19_n15}), .b ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, new_AGEMA_signal_1045, SB_19_n14}), .c ({SubC_out_s3[115], SubC_out_s2[115], SubC_out_s1[115], SubC_out_s0[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U9 ( .a ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, new_AGEMA_signal_1045, SB_19_n14}), .b ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, new_AGEMA_signal_1063, SB_19_T2}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, new_AGEMA_signal_1819, SB_19_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U6 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, new_AGEMA_signal_2269, SB_19_n11}), .b ({new_AGEMA_signal_1062, new_AGEMA_signal_1061, new_AGEMA_signal_1060, SB_19_T1}), .c ({SubC_out_s3[83], SubC_out_s2[83], SubC_out_s1[83], SubC_out_s0[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U5 ( .a ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, new_AGEMA_signal_1822, SB_19_n15}), .b ({SubC_in_s3[51], SubC_in_s2[51], SubC_in_s1[51], SubC_in_s0[51]}), .c ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, new_AGEMA_signal_2269, SB_19_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U4 ( .a ({new_AGEMA_signal_1056, new_AGEMA_signal_1055, new_AGEMA_signal_1054, SB_19_n10}), .b ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, new_AGEMA_signal_1057, SB_19_T0}), .c ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, new_AGEMA_signal_1822, SB_19_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U1 ( .a ({SubC_in_s3[115], SubC_in_s2[115], SubC_in_s1[115], SubC_in_s0[115]}), .b ({new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, SB_19_T3}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, new_AGEMA_signal_1825, SB_19_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_19_t0_AND_U1 ( .a ({SubC_in_s3[115], SubC_in_s2[115], SubC_in_s1[115], SubC_in_s0[115]}), .b ({SubC_in_s3[83], SubC_in_s2[83], SubC_in_s1[83], SubC_in_s0[83]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, new_AGEMA_signal_1057, SB_19_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_19_t1_AND_U1 ( .a ({SubC_in_s3[115], SubC_in_s2[115], SubC_in_s1[115], SubC_in_s0[115]}), .b ({SubC_in_s3[51], SubC_in_s2[51], SubC_in_s1[51], SubC_in_s0[51]}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1062, new_AGEMA_signal_1061, new_AGEMA_signal_1060, SB_19_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_19_t2_AND_U1 ( .a ({SubC_in_s3[115], SubC_in_s2[115], SubC_in_s1[115], SubC_in_s0[115]}), .b ({SubC_in_s3[19], SubC_in_s2[19], SubC_in_s1[19], SubC_in_s0[19]}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, new_AGEMA_signal_1063, SB_19_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_19_t3_AND_U1 ( .a ({SubC_in_s3[83], SubC_in_s2[83], SubC_in_s1[83], SubC_in_s0[83]}), .b ({SubC_in_s3[19], SubC_in_s2[19], SubC_in_s1[19], SubC_in_s0[19]}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, SB_19_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U11 ( .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, new_AGEMA_signal_1837, SB_18_n15}), .b ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, SB_18_n14}), .c ({SubC_out_s3[114], SubC_out_s2[114], SubC_out_s1[114], SubC_out_s0[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U9 ( .a ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, new_AGEMA_signal_1075, SB_18_n14}), .b ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, new_AGEMA_signal_1093, SB_18_T2}), .c ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, new_AGEMA_signal_1834, SB_18_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U6 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, SB_18_n11}), .b ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, SB_18_T1}), .c ({SubC_out_s3[82], SubC_out_s2[82], SubC_out_s1[82], SubC_out_s0[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U5 ( .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, new_AGEMA_signal_1837, SB_18_n15}), .b ({SubC_in_s3[50], SubC_in_s2[50], SubC_in_s1[50], SubC_in_s0[50]}), .c ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, SB_18_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U4 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, SB_18_n10}), .b ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, new_AGEMA_signal_1087, SB_18_T0}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, new_AGEMA_signal_1837, SB_18_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U1 ( .a ({SubC_in_s3[114], SubC_in_s2[114], SubC_in_s1[114], SubC_in_s0[114]}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, SB_18_T3}), .c ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, SB_18_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_18_t0_AND_U1 ( .a ({SubC_in_s3[114], SubC_in_s2[114], SubC_in_s1[114], SubC_in_s0[114]}), .b ({SubC_in_s3[82], SubC_in_s2[82], SubC_in_s1[82], SubC_in_s0[82]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, new_AGEMA_signal_1087, SB_18_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_18_t1_AND_U1 ( .a ({SubC_in_s3[114], SubC_in_s2[114], SubC_in_s1[114], SubC_in_s0[114]}), .b ({SubC_in_s3[50], SubC_in_s2[50], SubC_in_s1[50], SubC_in_s0[50]}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, SB_18_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_18_t2_AND_U1 ( .a ({SubC_in_s3[114], SubC_in_s2[114], SubC_in_s1[114], SubC_in_s0[114]}), .b ({SubC_in_s3[18], SubC_in_s2[18], SubC_in_s1[18], SubC_in_s0[18]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, new_AGEMA_signal_1093, SB_18_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_18_t3_AND_U1 ( .a ({SubC_in_s3[82], SubC_in_s2[82], SubC_in_s1[82], SubC_in_s0[82]}), .b ({SubC_in_s3[18], SubC_in_s2[18], SubC_in_s1[18], SubC_in_s0[18]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, SB_18_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U11 ( .a ({new_AGEMA_signal_1854, new_AGEMA_signal_1853, new_AGEMA_signal_1852, SB_17_n15}), .b ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, new_AGEMA_signal_1105, SB_17_n14}), .c ({SubC_out_s3[113], SubC_out_s2[113], SubC_out_s1[113], SubC_out_s0[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U9 ( .a ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, new_AGEMA_signal_1105, SB_17_n14}), .b ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, new_AGEMA_signal_1123, SB_17_T2}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, new_AGEMA_signal_1849, SB_17_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U6 ( .a ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, new_AGEMA_signal_2293, SB_17_n11}), .b ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, new_AGEMA_signal_1120, SB_17_T1}), .c ({SubC_out_s3[81], SubC_out_s2[81], SubC_out_s1[81], SubC_out_s0[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U5 ( .a ({new_AGEMA_signal_1854, new_AGEMA_signal_1853, new_AGEMA_signal_1852, SB_17_n15}), .b ({SubC_in_s3[49], SubC_in_s2[49], SubC_in_s1[49], SubC_in_s0[49]}), .c ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, new_AGEMA_signal_2293, SB_17_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U4 ( .a ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, new_AGEMA_signal_1114, SB_17_n10}), .b ({new_AGEMA_signal_1119, new_AGEMA_signal_1118, new_AGEMA_signal_1117, SB_17_T0}), .c ({new_AGEMA_signal_1854, new_AGEMA_signal_1853, new_AGEMA_signal_1852, SB_17_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U1 ( .a ({SubC_in_s3[113], SubC_in_s2[113], SubC_in_s1[113], SubC_in_s0[113]}), .b ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, SB_17_T3}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, new_AGEMA_signal_1855, SB_17_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_17_t0_AND_U1 ( .a ({SubC_in_s3[113], SubC_in_s2[113], SubC_in_s1[113], SubC_in_s0[113]}), .b ({SubC_in_s3[81], SubC_in_s2[81], SubC_in_s1[81], SubC_in_s0[81]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1119, new_AGEMA_signal_1118, new_AGEMA_signal_1117, SB_17_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_17_t1_AND_U1 ( .a ({SubC_in_s3[113], SubC_in_s2[113], SubC_in_s1[113], SubC_in_s0[113]}), .b ({SubC_in_s3[49], SubC_in_s2[49], SubC_in_s1[49], SubC_in_s0[49]}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, new_AGEMA_signal_1120, SB_17_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_17_t2_AND_U1 ( .a ({SubC_in_s3[113], SubC_in_s2[113], SubC_in_s1[113], SubC_in_s0[113]}), .b ({SubC_in_s3[17], SubC_in_s2[17], SubC_in_s1[17], SubC_in_s0[17]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, new_AGEMA_signal_1123, SB_17_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_17_t3_AND_U1 ( .a ({SubC_in_s3[81], SubC_in_s2[81], SubC_in_s1[81], SubC_in_s0[81]}), .b ({SubC_in_s3[17], SubC_in_s2[17], SubC_in_s1[17], SubC_in_s0[17]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, SB_17_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U11 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, SB_16_n15}), .b ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, new_AGEMA_signal_1135, SB_16_n14}), .c ({SubC_out_s3[112], SubC_out_s2[112], SubC_out_s1[112], SubC_out_s0[112]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U9 ( .a ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, new_AGEMA_signal_1135, SB_16_n14}), .b ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, new_AGEMA_signal_1153, SB_16_T2}), .c ({new_AGEMA_signal_1866, new_AGEMA_signal_1865, new_AGEMA_signal_1864, SB_16_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U6 ( .a ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, new_AGEMA_signal_2305, SB_16_n11}), .b ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, SB_16_T1}), .c ({SubC_out_s3[80], SubC_out_s2[80], SubC_out_s1[80], SubC_out_s0[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U5 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, SB_16_n15}), .b ({SubC_in_s3[48], SubC_in_s2[48], SubC_in_s1[48], SubC_in_s0[48]}), .c ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, new_AGEMA_signal_2305, SB_16_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U4 ( .a ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, new_AGEMA_signal_1144, SB_16_n10}), .b ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, new_AGEMA_signal_1147, SB_16_T0}), .c ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, SB_16_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U1 ( .a ({SubC_in_s3[112], SubC_in_s2[112], SubC_in_s1[112], SubC_in_s0[112]}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, SB_16_T3}), .c ({new_AGEMA_signal_1872, new_AGEMA_signal_1871, new_AGEMA_signal_1870, SB_16_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_16_t0_AND_U1 ( .a ({SubC_in_s3[112], SubC_in_s2[112], SubC_in_s1[112], SubC_in_s0[112]}), .b ({SubC_in_s3[80], SubC_in_s2[80], SubC_in_s1[80], SubC_in_s0[80]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, new_AGEMA_signal_1147, SB_16_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_16_t1_AND_U1 ( .a ({SubC_in_s3[112], SubC_in_s2[112], SubC_in_s1[112], SubC_in_s0[112]}), .b ({SubC_in_s3[48], SubC_in_s2[48], SubC_in_s1[48], SubC_in_s0[48]}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, SB_16_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_16_t2_AND_U1 ( .a ({SubC_in_s3[112], SubC_in_s2[112], SubC_in_s1[112], SubC_in_s0[112]}), .b ({SubC_in_s3[16], SubC_in_s2[16], SubC_in_s1[16], SubC_in_s0[16]}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, new_AGEMA_signal_1153, SB_16_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_16_t3_AND_U1 ( .a ({SubC_in_s3[80], SubC_in_s2[80], SubC_in_s1[80], SubC_in_s0[80]}), .b ({SubC_in_s3[16], SubC_in_s2[16], SubC_in_s1[16], SubC_in_s0[16]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, SB_16_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U11 ( .a ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, new_AGEMA_signal_1882, SB_15_n15}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, new_AGEMA_signal_1165, SB_15_n14}), .c ({SubC_out_s3[111], SubC_out_s2[111], SubC_out_s1[111], SubC_out_s0[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U9 ( .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, new_AGEMA_signal_1165, SB_15_n14}), .b ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, SB_15_T2}), .c ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, new_AGEMA_signal_1879, SB_15_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U6 ( .a ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, new_AGEMA_signal_2317, SB_15_n11}), .b ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, new_AGEMA_signal_1180, SB_15_T1}), .c ({SubC_out_s3[79], SubC_out_s2[79], SubC_out_s1[79], SubC_out_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U5 ( .a ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, new_AGEMA_signal_1882, SB_15_n15}), .b ({SubC_in_s3[47], SubC_in_s2[47], SubC_in_s1[47], SubC_in_s0[47]}), .c ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, new_AGEMA_signal_2317, SB_15_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U4 ( .a ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, new_AGEMA_signal_1174, SB_15_n10}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, new_AGEMA_signal_1177, SB_15_T0}), .c ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, new_AGEMA_signal_1882, SB_15_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U1 ( .a ({SubC_in_s3[111], SubC_in_s2[111], SubC_in_s1[111], SubC_in_s0[111]}), .b ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, new_AGEMA_signal_1186, SB_15_T3}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, new_AGEMA_signal_1885, SB_15_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_15_t0_AND_U1 ( .a ({SubC_in_s3[111], SubC_in_s2[111], SubC_in_s1[111], SubC_in_s0[111]}), .b ({SubC_in_s3[79], SubC_in_s2[79], SubC_in_s1[79], SubC_in_s0[79]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, new_AGEMA_signal_1177, SB_15_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_15_t1_AND_U1 ( .a ({SubC_in_s3[111], SubC_in_s2[111], SubC_in_s1[111], SubC_in_s0[111]}), .b ({SubC_in_s3[47], SubC_in_s2[47], SubC_in_s1[47], SubC_in_s0[47]}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, new_AGEMA_signal_1180, SB_15_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_15_t2_AND_U1 ( .a ({SubC_in_s3[111], SubC_in_s2[111], SubC_in_s1[111], SubC_in_s0[111]}), .b ({SubC_in_s3[15], SubC_in_s2[15], SubC_in_s1[15], SubC_in_s0[15]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, SB_15_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_15_t3_AND_U1 ( .a ({SubC_in_s3[79], SubC_in_s2[79], SubC_in_s1[79], SubC_in_s0[79]}), .b ({SubC_in_s3[15], SubC_in_s2[15], SubC_in_s1[15], SubC_in_s0[15]}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, new_AGEMA_signal_1186, SB_15_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U11 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, new_AGEMA_signal_1897, SB_14_n15}), .b ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, SB_14_n14}), .c ({SubC_out_s3[110], SubC_out_s2[110], SubC_out_s1[110], SubC_out_s0[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U9 ( .a ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, SB_14_n14}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, new_AGEMA_signal_1213, SB_14_T2}), .c ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, SB_14_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U6 ( .a ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, SB_14_n11}), .b ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, new_AGEMA_signal_1210, SB_14_T1}), .c ({SubC_out_s3[78], SubC_out_s2[78], SubC_out_s1[78], SubC_out_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U5 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, new_AGEMA_signal_1897, SB_14_n15}), .b ({SubC_in_s3[46], SubC_in_s2[46], SubC_in_s1[46], SubC_in_s0[46]}), .c ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, SB_14_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U4 ( .a ({new_AGEMA_signal_1206, new_AGEMA_signal_1205, new_AGEMA_signal_1204, SB_14_n10}), .b ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, SB_14_T0}), .c ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, new_AGEMA_signal_1897, SB_14_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U1 ( .a ({SubC_in_s3[110], SubC_in_s2[110], SubC_in_s1[110], SubC_in_s0[110]}), .b ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, new_AGEMA_signal_1216, SB_14_T3}), .c ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, new_AGEMA_signal_1900, SB_14_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_14_t0_AND_U1 ( .a ({SubC_in_s3[110], SubC_in_s2[110], SubC_in_s1[110], SubC_in_s0[110]}), .b ({SubC_in_s3[78], SubC_in_s2[78], SubC_in_s1[78], SubC_in_s0[78]}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, SB_14_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_14_t1_AND_U1 ( .a ({SubC_in_s3[110], SubC_in_s2[110], SubC_in_s1[110], SubC_in_s0[110]}), .b ({SubC_in_s3[46], SubC_in_s2[46], SubC_in_s1[46], SubC_in_s0[46]}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, new_AGEMA_signal_1210, SB_14_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_14_t2_AND_U1 ( .a ({SubC_in_s3[110], SubC_in_s2[110], SubC_in_s1[110], SubC_in_s0[110]}), .b ({SubC_in_s3[14], SubC_in_s2[14], SubC_in_s1[14], SubC_in_s0[14]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, new_AGEMA_signal_1213, SB_14_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_14_t3_AND_U1 ( .a ({SubC_in_s3[78], SubC_in_s2[78], SubC_in_s1[78], SubC_in_s0[78]}), .b ({SubC_in_s3[14], SubC_in_s2[14], SubC_in_s1[14], SubC_in_s0[14]}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, new_AGEMA_signal_1216, SB_14_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U11 ( .a ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, new_AGEMA_signal_1912, SB_13_n15}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, new_AGEMA_signal_1225, SB_13_n14}), .c ({SubC_out_s3[109], SubC_out_s2[109], SubC_out_s1[109], SubC_out_s0[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U9 ( .a ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, new_AGEMA_signal_1225, SB_13_n14}), .b ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, SB_13_T2}), .c ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, new_AGEMA_signal_1909, SB_13_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U6 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, SB_13_n11}), .b ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, new_AGEMA_signal_1240, SB_13_T1}), .c ({SubC_out_s3[77], SubC_out_s2[77], SubC_out_s1[77], SubC_out_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U5 ( .a ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, new_AGEMA_signal_1912, SB_13_n15}), .b ({SubC_in_s3[45], SubC_in_s2[45], SubC_in_s1[45], SubC_in_s0[45]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, SB_13_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U4 ( .a ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, new_AGEMA_signal_1234, SB_13_n10}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, new_AGEMA_signal_1237, SB_13_T0}), .c ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, new_AGEMA_signal_1912, SB_13_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U1 ( .a ({SubC_in_s3[109], SubC_in_s2[109], SubC_in_s1[109], SubC_in_s0[109]}), .b ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, new_AGEMA_signal_1246, SB_13_T3}), .c ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, new_AGEMA_signal_1915, SB_13_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_13_t0_AND_U1 ( .a ({SubC_in_s3[109], SubC_in_s2[109], SubC_in_s1[109], SubC_in_s0[109]}), .b ({SubC_in_s3[77], SubC_in_s2[77], SubC_in_s1[77], SubC_in_s0[77]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, new_AGEMA_signal_1237, SB_13_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_13_t1_AND_U1 ( .a ({SubC_in_s3[109], SubC_in_s2[109], SubC_in_s1[109], SubC_in_s0[109]}), .b ({SubC_in_s3[45], SubC_in_s2[45], SubC_in_s1[45], SubC_in_s0[45]}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, new_AGEMA_signal_1240, SB_13_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_13_t2_AND_U1 ( .a ({SubC_in_s3[109], SubC_in_s2[109], SubC_in_s1[109], SubC_in_s0[109]}), .b ({SubC_in_s3[13], SubC_in_s2[13], SubC_in_s1[13], SubC_in_s0[13]}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, SB_13_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_13_t3_AND_U1 ( .a ({SubC_in_s3[77], SubC_in_s2[77], SubC_in_s1[77], SubC_in_s0[77]}), .b ({SubC_in_s3[13], SubC_in_s2[13], SubC_in_s1[13], SubC_in_s0[13]}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, new_AGEMA_signal_1246, SB_13_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U11 ( .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, SB_12_n15}), .b ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, new_AGEMA_signal_1255, SB_12_n14}), .c ({SubC_out_s3[108], SubC_out_s2[108], SubC_out_s1[108], SubC_out_s0[108]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U9 ( .a ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, new_AGEMA_signal_1255, SB_12_n14}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, new_AGEMA_signal_1273, SB_12_T2}), .c ({new_AGEMA_signal_1926, new_AGEMA_signal_1925, new_AGEMA_signal_1924, SB_12_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U6 ( .a ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, SB_12_n11}), .b ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, SB_12_T1}), .c ({SubC_out_s3[76], SubC_out_s2[76], SubC_out_s1[76], SubC_out_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U5 ( .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, SB_12_n15}), .b ({SubC_in_s3[44], SubC_in_s2[44], SubC_in_s1[44], SubC_in_s0[44]}), .c ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, SB_12_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U4 ( .a ({new_AGEMA_signal_1266, new_AGEMA_signal_1265, new_AGEMA_signal_1264, SB_12_n10}), .b ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, SB_12_T0}), .c ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, SB_12_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U1 ( .a ({SubC_in_s3[108], SubC_in_s2[108], SubC_in_s1[108], SubC_in_s0[108]}), .b ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, new_AGEMA_signal_1276, SB_12_T3}), .c ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, SB_12_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_12_t0_AND_U1 ( .a ({SubC_in_s3[108], SubC_in_s2[108], SubC_in_s1[108], SubC_in_s0[108]}), .b ({SubC_in_s3[76], SubC_in_s2[76], SubC_in_s1[76], SubC_in_s0[76]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, SB_12_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_12_t1_AND_U1 ( .a ({SubC_in_s3[108], SubC_in_s2[108], SubC_in_s1[108], SubC_in_s0[108]}), .b ({SubC_in_s3[44], SubC_in_s2[44], SubC_in_s1[44], SubC_in_s0[44]}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, SB_12_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_12_t2_AND_U1 ( .a ({SubC_in_s3[108], SubC_in_s2[108], SubC_in_s1[108], SubC_in_s0[108]}), .b ({SubC_in_s3[12], SubC_in_s2[12], SubC_in_s1[12], SubC_in_s0[12]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, new_AGEMA_signal_1273, SB_12_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_12_t3_AND_U1 ( .a ({SubC_in_s3[76], SubC_in_s2[76], SubC_in_s1[76], SubC_in_s0[76]}), .b ({SubC_in_s3[12], SubC_in_s2[12], SubC_in_s1[12], SubC_in_s0[12]}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, new_AGEMA_signal_1276, SB_12_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U11 ( .a ({new_AGEMA_signal_1944, new_AGEMA_signal_1943, new_AGEMA_signal_1942, SB_11_n15}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, new_AGEMA_signal_1285, SB_11_n14}), .c ({SubC_out_s3[107], SubC_out_s2[107], SubC_out_s1[107], SubC_out_s0[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U9 ( .a ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, new_AGEMA_signal_1285, SB_11_n14}), .b ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, new_AGEMA_signal_1303, SB_11_T2}), .c ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, new_AGEMA_signal_1939, SB_11_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U6 ( .a ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, new_AGEMA_signal_2365, SB_11_n11}), .b ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, new_AGEMA_signal_1300, SB_11_T1}), .c ({SubC_out_s3[75], SubC_out_s2[75], SubC_out_s1[75], SubC_out_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U5 ( .a ({new_AGEMA_signal_1944, new_AGEMA_signal_1943, new_AGEMA_signal_1942, SB_11_n15}), .b ({SubC_in_s3[43], SubC_in_s2[43], SubC_in_s1[43], SubC_in_s0[43]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, new_AGEMA_signal_2365, SB_11_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U4 ( .a ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, new_AGEMA_signal_1294, SB_11_n10}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, new_AGEMA_signal_1297, SB_11_T0}), .c ({new_AGEMA_signal_1944, new_AGEMA_signal_1943, new_AGEMA_signal_1942, SB_11_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U1 ( .a ({SubC_in_s3[107], SubC_in_s2[107], SubC_in_s1[107], SubC_in_s0[107]}), .b ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, SB_11_T3}), .c ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, new_AGEMA_signal_1945, SB_11_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_11_t0_AND_U1 ( .a ({SubC_in_s3[107], SubC_in_s2[107], SubC_in_s1[107], SubC_in_s0[107]}), .b ({SubC_in_s3[75], SubC_in_s2[75], SubC_in_s1[75], SubC_in_s0[75]}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, new_AGEMA_signal_1297, SB_11_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_11_t1_AND_U1 ( .a ({SubC_in_s3[107], SubC_in_s2[107], SubC_in_s1[107], SubC_in_s0[107]}), .b ({SubC_in_s3[43], SubC_in_s2[43], SubC_in_s1[43], SubC_in_s0[43]}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, new_AGEMA_signal_1300, SB_11_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_11_t2_AND_U1 ( .a ({SubC_in_s3[107], SubC_in_s2[107], SubC_in_s1[107], SubC_in_s0[107]}), .b ({SubC_in_s3[11], SubC_in_s2[11], SubC_in_s1[11], SubC_in_s0[11]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, new_AGEMA_signal_1303, SB_11_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_11_t3_AND_U1 ( .a ({SubC_in_s3[75], SubC_in_s2[75], SubC_in_s1[75], SubC_in_s0[75]}), .b ({SubC_in_s3[11], SubC_in_s2[11], SubC_in_s1[11], SubC_in_s0[11]}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, SB_11_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U11 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, SB_10_n15}), .b ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, SB_10_n14}), .c ({SubC_out_s3[106], SubC_out_s2[106], SubC_out_s1[106], SubC_out_s0[106]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U9 ( .a ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, SB_10_n14}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, new_AGEMA_signal_1333, SB_10_T2}), .c ({new_AGEMA_signal_1956, new_AGEMA_signal_1955, new_AGEMA_signal_1954, SB_10_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U6 ( .a ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, SB_10_n11}), .b ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, SB_10_T1}), .c ({SubC_out_s3[74], SubC_out_s2[74], SubC_out_s1[74], SubC_out_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U5 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, SB_10_n15}), .b ({SubC_in_s3[42], SubC_in_s2[42], SubC_in_s1[42], SubC_in_s0[42]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, SB_10_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U4 ( .a ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, new_AGEMA_signal_1324, SB_10_n10}), .b ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, SB_10_T0}), .c ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, SB_10_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U1 ( .a ({SubC_in_s3[106], SubC_in_s2[106], SubC_in_s1[106], SubC_in_s0[106]}), .b ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, new_AGEMA_signal_1336, SB_10_T3}), .c ({new_AGEMA_signal_1962, new_AGEMA_signal_1961, new_AGEMA_signal_1960, SB_10_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_10_t0_AND_U1 ( .a ({SubC_in_s3[106], SubC_in_s2[106], SubC_in_s1[106], SubC_in_s0[106]}), .b ({SubC_in_s3[74], SubC_in_s2[74], SubC_in_s1[74], SubC_in_s0[74]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, SB_10_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_10_t1_AND_U1 ( .a ({SubC_in_s3[106], SubC_in_s2[106], SubC_in_s1[106], SubC_in_s0[106]}), .b ({SubC_in_s3[42], SubC_in_s2[42], SubC_in_s1[42], SubC_in_s0[42]}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, SB_10_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_10_t2_AND_U1 ( .a ({SubC_in_s3[106], SubC_in_s2[106], SubC_in_s1[106], SubC_in_s0[106]}), .b ({SubC_in_s3[10], SubC_in_s2[10], SubC_in_s1[10], SubC_in_s0[10]}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, new_AGEMA_signal_1333, SB_10_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_10_t3_AND_U1 ( .a ({SubC_in_s3[74], SubC_in_s2[74], SubC_in_s1[74], SubC_in_s0[74]}), .b ({SubC_in_s3[10], SubC_in_s2[10], SubC_in_s1[10], SubC_in_s0[10]}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, new_AGEMA_signal_1336, SB_10_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U11 ( .a ({new_AGEMA_signal_1974, new_AGEMA_signal_1973, new_AGEMA_signal_1972, SB_9_n15}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, new_AGEMA_signal_1345, SB_9_n14}), .c ({SubC_out_s3[105], SubC_out_s2[105], SubC_out_s1[105], SubC_out_s0[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U9 ( .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, new_AGEMA_signal_1345, SB_9_n14}), .b ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, new_AGEMA_signal_1363, SB_9_T2}), .c ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, new_AGEMA_signal_1969, SB_9_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U6 ( .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, SB_9_n11}), .b ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, new_AGEMA_signal_1360, SB_9_T1}), .c ({SubC_out_s3[73], SubC_out_s2[73], SubC_out_s1[73], SubC_out_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U5 ( .a ({new_AGEMA_signal_1974, new_AGEMA_signal_1973, new_AGEMA_signal_1972, SB_9_n15}), .b ({SubC_in_s3[41], SubC_in_s2[41], SubC_in_s1[41], SubC_in_s0[41]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, SB_9_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U4 ( .a ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, new_AGEMA_signal_1354, SB_9_n10}), .b ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, new_AGEMA_signal_1357, SB_9_T0}), .c ({new_AGEMA_signal_1974, new_AGEMA_signal_1973, new_AGEMA_signal_1972, SB_9_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U1 ( .a ({SubC_in_s3[105], SubC_in_s2[105], SubC_in_s1[105], SubC_in_s0[105]}), .b ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, SB_9_T3}), .c ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, SB_9_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_9_t0_AND_U1 ( .a ({SubC_in_s3[105], SubC_in_s2[105], SubC_in_s1[105], SubC_in_s0[105]}), .b ({SubC_in_s3[73], SubC_in_s2[73], SubC_in_s1[73], SubC_in_s0[73]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, new_AGEMA_signal_1357, SB_9_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_9_t1_AND_U1 ( .a ({SubC_in_s3[105], SubC_in_s2[105], SubC_in_s1[105], SubC_in_s0[105]}), .b ({SubC_in_s3[41], SubC_in_s2[41], SubC_in_s1[41], SubC_in_s0[41]}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, new_AGEMA_signal_1360, SB_9_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_9_t2_AND_U1 ( .a ({SubC_in_s3[105], SubC_in_s2[105], SubC_in_s1[105], SubC_in_s0[105]}), .b ({SubC_in_s3[9], SubC_in_s2[9], SubC_in_s1[9], SubC_in_s0[9]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, new_AGEMA_signal_1363, SB_9_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_9_t3_AND_U1 ( .a ({SubC_in_s3[73], SubC_in_s2[73], SubC_in_s1[73], SubC_in_s0[73]}), .b ({SubC_in_s3[9], SubC_in_s2[9], SubC_in_s1[9], SubC_in_s0[9]}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, SB_9_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U11 ( .a ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, new_AGEMA_signal_1987, SB_8_n15}), .b ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, SB_8_n14}), .c ({SubC_out_s3[104], SubC_out_s2[104], SubC_out_s1[104], SubC_out_s0[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U9 ( .a ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, SB_8_n14}), .b ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, new_AGEMA_signal_1393, SB_8_T2}), .c ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, new_AGEMA_signal_1984, SB_8_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U6 ( .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, SB_8_n11}), .b ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, new_AGEMA_signal_1390, SB_8_T1}), .c ({SubC_out_s3[72], SubC_out_s2[72], SubC_out_s1[72], SubC_out_s0[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U5 ( .a ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, new_AGEMA_signal_1987, SB_8_n15}), .b ({SubC_in_s3[40], SubC_in_s2[40], SubC_in_s1[40], SubC_in_s0[40]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, SB_8_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U4 ( .a ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, new_AGEMA_signal_1384, SB_8_n10}), .b ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, SB_8_T0}), .c ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, new_AGEMA_signal_1987, SB_8_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U1 ( .a ({SubC_in_s3[104], SubC_in_s2[104], SubC_in_s1[104], SubC_in_s0[104]}), .b ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, new_AGEMA_signal_1396, SB_8_T3}), .c ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, new_AGEMA_signal_1990, SB_8_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_8_t0_AND_U1 ( .a ({SubC_in_s3[104], SubC_in_s2[104], SubC_in_s1[104], SubC_in_s0[104]}), .b ({SubC_in_s3[72], SubC_in_s2[72], SubC_in_s1[72], SubC_in_s0[72]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, SB_8_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_8_t1_AND_U1 ( .a ({SubC_in_s3[104], SubC_in_s2[104], SubC_in_s1[104], SubC_in_s0[104]}), .b ({SubC_in_s3[40], SubC_in_s2[40], SubC_in_s1[40], SubC_in_s0[40]}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, new_AGEMA_signal_1390, SB_8_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_8_t2_AND_U1 ( .a ({SubC_in_s3[104], SubC_in_s2[104], SubC_in_s1[104], SubC_in_s0[104]}), .b ({SubC_in_s3[8], SubC_in_s2[8], SubC_in_s1[8], SubC_in_s0[8]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, new_AGEMA_signal_1393, SB_8_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_8_t3_AND_U1 ( .a ({SubC_in_s3[72], SubC_in_s2[72], SubC_in_s1[72], SubC_in_s0[72]}), .b ({SubC_in_s3[8], SubC_in_s2[8], SubC_in_s1[8], SubC_in_s0[8]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, new_AGEMA_signal_1396, SB_8_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U11 ( .a ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, SB_7_n15}), .b ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, new_AGEMA_signal_1405, SB_7_n14}), .c ({SubC_out_s3[103], SubC_out_s2[103], SubC_out_s1[103], SubC_out_s0[103]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U9 ( .a ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, new_AGEMA_signal_1405, SB_7_n14}), .b ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, SB_7_T2}), .c ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, new_AGEMA_signal_1999, SB_7_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U6 ( .a ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2413, SB_7_n11}), .b ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, new_AGEMA_signal_1420, SB_7_T1}), .c ({SubC_out_s3[71], SubC_out_s2[71], SubC_out_s1[71], SubC_out_s0[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U5 ( .a ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, SB_7_n15}), .b ({SubC_in_s3[39], SubC_in_s2[39], SubC_in_s1[39], SubC_in_s0[39]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2413, SB_7_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U4 ( .a ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, new_AGEMA_signal_1414, SB_7_n10}), .b ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, new_AGEMA_signal_1417, SB_7_T0}), .c ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, new_AGEMA_signal_2002, SB_7_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U1 ( .a ({SubC_in_s3[103], SubC_in_s2[103], SubC_in_s1[103], SubC_in_s0[103]}), .b ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, SB_7_T3}), .c ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, new_AGEMA_signal_2005, SB_7_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_7_t0_AND_U1 ( .a ({SubC_in_s3[103], SubC_in_s2[103], SubC_in_s1[103], SubC_in_s0[103]}), .b ({SubC_in_s3[71], SubC_in_s2[71], SubC_in_s1[71], SubC_in_s0[71]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, new_AGEMA_signal_1417, SB_7_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_7_t1_AND_U1 ( .a ({SubC_in_s3[103], SubC_in_s2[103], SubC_in_s1[103], SubC_in_s0[103]}), .b ({SubC_in_s3[39], SubC_in_s2[39], SubC_in_s1[39], SubC_in_s0[39]}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, new_AGEMA_signal_1420, SB_7_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_7_t2_AND_U1 ( .a ({SubC_in_s3[103], SubC_in_s2[103], SubC_in_s1[103], SubC_in_s0[103]}), .b ({SubC_in_s3[7], SubC_in_s2[7], SubC_in_s1[7], SubC_in_s0[7]}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, SB_7_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_7_t3_AND_U1 ( .a ({SubC_in_s3[71], SubC_in_s2[71], SubC_in_s1[71], SubC_in_s0[71]}), .b ({SubC_in_s3[7], SubC_in_s2[7], SubC_in_s1[7], SubC_in_s0[7]}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, SB_7_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U11 ( .a ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, new_AGEMA_signal_2017, SB_6_n15}), .b ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, new_AGEMA_signal_1435, SB_6_n14}), .c ({SubC_out_s3[102], SubC_out_s2[102], SubC_out_s1[102], SubC_out_s0[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U9 ( .a ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, new_AGEMA_signal_1435, SB_6_n14}), .b ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, new_AGEMA_signal_1453, SB_6_T2}), .c ({new_AGEMA_signal_2016, new_AGEMA_signal_2015, new_AGEMA_signal_2014, SB_6_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U6 ( .a ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, SB_6_n11}), .b ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, new_AGEMA_signal_1450, SB_6_T1}), .c ({SubC_out_s3[70], SubC_out_s2[70], SubC_out_s1[70], SubC_out_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U5 ( .a ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, new_AGEMA_signal_2017, SB_6_n15}), .b ({SubC_in_s3[38], SubC_in_s2[38], SubC_in_s1[38], SubC_in_s0[38]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, SB_6_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U4 ( .a ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, new_AGEMA_signal_1444, SB_6_n10}), .b ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, SB_6_T0}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, new_AGEMA_signal_2017, SB_6_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U1 ( .a ({SubC_in_s3[102], SubC_in_s2[102], SubC_in_s1[102], SubC_in_s0[102]}), .b ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, new_AGEMA_signal_1456, SB_6_T3}), .c ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, SB_6_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_6_t0_AND_U1 ( .a ({SubC_in_s3[102], SubC_in_s2[102], SubC_in_s1[102], SubC_in_s0[102]}), .b ({SubC_in_s3[70], SubC_in_s2[70], SubC_in_s1[70], SubC_in_s0[70]}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, SB_6_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_6_t1_AND_U1 ( .a ({SubC_in_s3[102], SubC_in_s2[102], SubC_in_s1[102], SubC_in_s0[102]}), .b ({SubC_in_s3[38], SubC_in_s2[38], SubC_in_s1[38], SubC_in_s0[38]}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, new_AGEMA_signal_1450, SB_6_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_6_t2_AND_U1 ( .a ({SubC_in_s3[102], SubC_in_s2[102], SubC_in_s1[102], SubC_in_s0[102]}), .b ({SubC_in_s3[6], SubC_in_s2[6], SubC_in_s1[6], SubC_in_s0[6]}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, new_AGEMA_signal_1453, SB_6_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_6_t3_AND_U1 ( .a ({SubC_in_s3[70], SubC_in_s2[70], SubC_in_s1[70], SubC_in_s0[70]}), .b ({SubC_in_s3[6], SubC_in_s2[6], SubC_in_s1[6], SubC_in_s0[6]}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, new_AGEMA_signal_1456, SB_6_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U11 ( .a ({new_AGEMA_signal_2034, new_AGEMA_signal_2033, new_AGEMA_signal_2032, SB_5_n15}), .b ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, new_AGEMA_signal_1465, SB_5_n14}), .c ({SubC_out_s3[101], SubC_out_s2[101], SubC_out_s1[101], SubC_out_s0[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U9 ( .a ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, new_AGEMA_signal_1465, SB_5_n14}), .b ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, SB_5_T2}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, new_AGEMA_signal_2029, SB_5_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U6 ( .a ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, new_AGEMA_signal_2437, SB_5_n11}), .b ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, SB_5_T1}), .c ({SubC_out_s3[69], SubC_out_s2[69], SubC_out_s1[69], SubC_out_s0[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U5 ( .a ({new_AGEMA_signal_2034, new_AGEMA_signal_2033, new_AGEMA_signal_2032, SB_5_n15}), .b ({SubC_in_s3[37], SubC_in_s2[37], SubC_in_s1[37], SubC_in_s0[37]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, new_AGEMA_signal_2437, SB_5_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U4 ( .a ({new_AGEMA_signal_1476, new_AGEMA_signal_1475, new_AGEMA_signal_1474, SB_5_n10}), .b ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, new_AGEMA_signal_1477, SB_5_T0}), .c ({new_AGEMA_signal_2034, new_AGEMA_signal_2033, new_AGEMA_signal_2032, SB_5_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U1 ( .a ({SubC_in_s3[101], SubC_in_s2[101], SubC_in_s1[101], SubC_in_s0[101]}), .b ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, new_AGEMA_signal_1486, SB_5_T3}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, new_AGEMA_signal_2035, SB_5_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_5_t0_AND_U1 ( .a ({SubC_in_s3[101], SubC_in_s2[101], SubC_in_s1[101], SubC_in_s0[101]}), .b ({SubC_in_s3[69], SubC_in_s2[69], SubC_in_s1[69], SubC_in_s0[69]}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, new_AGEMA_signal_1477, SB_5_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_5_t1_AND_U1 ( .a ({SubC_in_s3[101], SubC_in_s2[101], SubC_in_s1[101], SubC_in_s0[101]}), .b ({SubC_in_s3[37], SubC_in_s2[37], SubC_in_s1[37], SubC_in_s0[37]}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, SB_5_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_5_t2_AND_U1 ( .a ({SubC_in_s3[101], SubC_in_s2[101], SubC_in_s1[101], SubC_in_s0[101]}), .b ({SubC_in_s3[5], SubC_in_s2[5], SubC_in_s1[5], SubC_in_s0[5]}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, SB_5_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_5_t3_AND_U1 ( .a ({SubC_in_s3[69], SubC_in_s2[69], SubC_in_s1[69], SubC_in_s0[69]}), .b ({SubC_in_s3[5], SubC_in_s2[5], SubC_in_s1[5], SubC_in_s0[5]}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, new_AGEMA_signal_1486, SB_5_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U11 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, SB_4_n15}), .b ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, new_AGEMA_signal_1495, SB_4_n14}), .c ({SubC_out_s3[100], SubC_out_s2[100], SubC_out_s1[100], SubC_out_s0[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U9 ( .a ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, new_AGEMA_signal_1495, SB_4_n14}), .b ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, new_AGEMA_signal_1513, SB_4_T2}), .c ({new_AGEMA_signal_2046, new_AGEMA_signal_2045, new_AGEMA_signal_2044, SB_4_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U6 ( .a ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, SB_4_n11}), .b ({new_AGEMA_signal_1512, new_AGEMA_signal_1511, new_AGEMA_signal_1510, SB_4_T1}), .c ({SubC_out_s3[68], SubC_out_s2[68], SubC_out_s1[68], SubC_out_s0[68]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U5 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, SB_4_n15}), .b ({SubC_in_s3[36], SubC_in_s2[36], SubC_in_s1[36], SubC_in_s0[36]}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, SB_4_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U4 ( .a ({new_AGEMA_signal_1506, new_AGEMA_signal_1505, new_AGEMA_signal_1504, SB_4_n10}), .b ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, SB_4_T0}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, SB_4_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U1 ( .a ({SubC_in_s3[100], SubC_in_s2[100], SubC_in_s1[100], SubC_in_s0[100]}), .b ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, SB_4_T3}), .c ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, new_AGEMA_signal_2050, SB_4_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_4_t0_AND_U1 ( .a ({SubC_in_s3[100], SubC_in_s2[100], SubC_in_s1[100], SubC_in_s0[100]}), .b ({SubC_in_s3[68], SubC_in_s2[68], SubC_in_s1[68], SubC_in_s0[68]}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, SB_4_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_4_t1_AND_U1 ( .a ({SubC_in_s3[100], SubC_in_s2[100], SubC_in_s1[100], SubC_in_s0[100]}), .b ({SubC_in_s3[36], SubC_in_s2[36], SubC_in_s1[36], SubC_in_s0[36]}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_1512, new_AGEMA_signal_1511, new_AGEMA_signal_1510, SB_4_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_4_t2_AND_U1 ( .a ({SubC_in_s3[100], SubC_in_s2[100], SubC_in_s1[100], SubC_in_s0[100]}), .b ({SubC_in_s3[4], SubC_in_s2[4], SubC_in_s1[4], SubC_in_s0[4]}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, new_AGEMA_signal_1513, SB_4_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_4_t3_AND_U1 ( .a ({SubC_in_s3[68], SubC_in_s2[68], SubC_in_s1[68], SubC_in_s0[68]}), .b ({SubC_in_s3[4], SubC_in_s2[4], SubC_in_s1[4], SubC_in_s0[4]}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, SB_4_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U11 ( .a ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, new_AGEMA_signal_2062, SB_3_n15}), .b ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, SB_3_n14}), .c ({SubC_out_s3[99], SubC_out_s2[99], SubC_out_s1[99], SubC_out_s0[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U9 ( .a ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, SB_3_n14}), .b ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, SB_3_T2}), .c ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, new_AGEMA_signal_2059, SB_3_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U6 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, new_AGEMA_signal_2461, SB_3_n11}), .b ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, new_AGEMA_signal_1540, SB_3_T1}), .c ({SubC_out_s3[67], SubC_out_s2[67], SubC_out_s1[67], SubC_out_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U5 ( .a ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, new_AGEMA_signal_2062, SB_3_n15}), .b ({SubC_in_s3[35], SubC_in_s2[35], SubC_in_s1[35], SubC_in_s0[35]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, new_AGEMA_signal_2461, SB_3_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U4 ( .a ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, new_AGEMA_signal_1534, SB_3_n10}), .b ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, new_AGEMA_signal_1537, SB_3_T0}), .c ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, new_AGEMA_signal_2062, SB_3_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U1 ( .a ({SubC_in_s3[99], SubC_in_s2[99], SubC_in_s1[99], SubC_in_s0[99]}), .b ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, new_AGEMA_signal_1546, SB_3_T3}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, new_AGEMA_signal_2065, SB_3_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_3_t0_AND_U1 ( .a ({SubC_in_s3[99], SubC_in_s2[99], SubC_in_s1[99], SubC_in_s0[99]}), .b ({SubC_in_s3[67], SubC_in_s2[67], SubC_in_s1[67], SubC_in_s0[67]}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, new_AGEMA_signal_1537, SB_3_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_3_t1_AND_U1 ( .a ({SubC_in_s3[99], SubC_in_s2[99], SubC_in_s1[99], SubC_in_s0[99]}), .b ({SubC_in_s3[35], SubC_in_s2[35], SubC_in_s1[35], SubC_in_s0[35]}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, new_AGEMA_signal_1540, SB_3_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_3_t2_AND_U1 ( .a ({SubC_in_s3[99], SubC_in_s2[99], SubC_in_s1[99], SubC_in_s0[99]}), .b ({SubC_in_s3[3], SubC_in_s2[3], SubC_in_s1[3], SubC_in_s0[3]}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, SB_3_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_3_t3_AND_U1 ( .a ({SubC_in_s3[67], SubC_in_s2[67], SubC_in_s1[67], SubC_in_s0[67]}), .b ({SubC_in_s3[3], SubC_in_s2[3], SubC_in_s1[3], SubC_in_s0[3]}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, new_AGEMA_signal_1546, SB_3_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U11 ( .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, new_AGEMA_signal_2077, SB_2_n15}), .b ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, new_AGEMA_signal_1555, SB_2_n14}), .c ({SubC_out_s3[98], SubC_out_s2[98], SubC_out_s1[98], SubC_out_s0[98]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U9 ( .a ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, new_AGEMA_signal_1555, SB_2_n14}), .b ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, new_AGEMA_signal_1573, SB_2_T2}), .c ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, SB_2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U6 ( .a ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, new_AGEMA_signal_2473, SB_2_n11}), .b ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, SB_2_T1}), .c ({SubC_out_s3[66], SubC_out_s2[66], SubC_out_s1[66], SubC_out_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U5 ( .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, new_AGEMA_signal_2077, SB_2_n15}), .b ({SubC_in_s3[34], SubC_in_s2[34], SubC_in_s1[34], SubC_in_s0[34]}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, new_AGEMA_signal_2473, SB_2_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U4 ( .a ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, new_AGEMA_signal_1564, SB_2_n10}), .b ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, new_AGEMA_signal_1567, SB_2_T0}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, new_AGEMA_signal_2077, SB_2_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U1 ( .a ({SubC_in_s3[98], SubC_in_s2[98], SubC_in_s1[98], SubC_in_s0[98]}), .b ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, new_AGEMA_signal_1576, SB_2_T3}), .c ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, SB_2_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_2_t0_AND_U1 ( .a ({SubC_in_s3[98], SubC_in_s2[98], SubC_in_s1[98], SubC_in_s0[98]}), .b ({SubC_in_s3[66], SubC_in_s2[66], SubC_in_s1[66], SubC_in_s0[66]}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, new_AGEMA_signal_1567, SB_2_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_2_t1_AND_U1 ( .a ({SubC_in_s3[98], SubC_in_s2[98], SubC_in_s1[98], SubC_in_s0[98]}), .b ({SubC_in_s3[34], SubC_in_s2[34], SubC_in_s1[34], SubC_in_s0[34]}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, SB_2_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_2_t2_AND_U1 ( .a ({SubC_in_s3[98], SubC_in_s2[98], SubC_in_s1[98], SubC_in_s0[98]}), .b ({SubC_in_s3[2], SubC_in_s2[2], SubC_in_s1[2], SubC_in_s0[2]}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, new_AGEMA_signal_1573, SB_2_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_2_t3_AND_U1 ( .a ({SubC_in_s3[66], SubC_in_s2[66], SubC_in_s1[66], SubC_in_s0[66]}), .b ({SubC_in_s3[2], SubC_in_s2[2], SubC_in_s1[2], SubC_in_s0[2]}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, new_AGEMA_signal_1576, SB_2_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U11 ( .a ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, new_AGEMA_signal_2092, SB_1_n15}), .b ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, new_AGEMA_signal_1585, SB_1_n14}), .c ({SubC_out_s3[97], SubC_out_s2[97], SubC_out_s1[97], SubC_out_s0[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U9 ( .a ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, new_AGEMA_signal_1585, SB_1_n14}), .b ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, new_AGEMA_signal_1603, SB_1_T2}), .c ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, new_AGEMA_signal_2089, SB_1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U6 ( .a ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, new_AGEMA_signal_2485, SB_1_n11}), .b ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, new_AGEMA_signal_1600, SB_1_T1}), .c ({SubC_out_s3[65], SubC_out_s2[65], SubC_out_s1[65], SubC_out_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U5 ( .a ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, new_AGEMA_signal_2092, SB_1_n15}), .b ({SubC_in_s3[33], SubC_in_s2[33], SubC_in_s1[33], SubC_in_s0[33]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, new_AGEMA_signal_2485, SB_1_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U4 ( .a ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, new_AGEMA_signal_1594, SB_1_n10}), .b ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, SB_1_T0}), .c ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, new_AGEMA_signal_2092, SB_1_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U1 ( .a ({SubC_in_s3[97], SubC_in_s2[97], SubC_in_s1[97], SubC_in_s0[97]}), .b ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, SB_1_T3}), .c ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, SB_1_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_1_t0_AND_U1 ( .a ({SubC_in_s3[97], SubC_in_s2[97], SubC_in_s1[97], SubC_in_s0[97]}), .b ({SubC_in_s3[65], SubC_in_s2[65], SubC_in_s1[65], SubC_in_s0[65]}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, SB_1_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_1_t1_AND_U1 ( .a ({SubC_in_s3[97], SubC_in_s2[97], SubC_in_s1[97], SubC_in_s0[97]}), .b ({SubC_in_s3[33], SubC_in_s2[33], SubC_in_s1[33], SubC_in_s0[33]}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, new_AGEMA_signal_1600, SB_1_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_1_t2_AND_U1 ( .a ({SubC_in_s3[97], SubC_in_s2[97], SubC_in_s1[97], SubC_in_s0[97]}), .b ({SubC_in_s3[1], SubC_in_s2[1], SubC_in_s1[1], SubC_in_s0[1]}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, new_AGEMA_signal_1603, SB_1_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_1_t3_AND_U1 ( .a ({SubC_in_s3[65], SubC_in_s2[65], SubC_in_s1[65], SubC_in_s0[65]}), .b ({SubC_in_s3[1], SubC_in_s2[1], SubC_in_s1[1], SubC_in_s0[1]}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, SB_1_T3}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U11 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, SB_0_n15}), .b ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, SB_0_n14}), .c ({SubC_out_s3[96], SubC_out_s2[96], SubC_out_s1[96], SubC_out_s0[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U9 ( .a ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, SB_0_n14}), .b ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, SB_0_T2}), .c ({new_AGEMA_signal_2106, new_AGEMA_signal_2105, new_AGEMA_signal_2104, SB_0_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U6 ( .a ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, new_AGEMA_signal_2497, SB_0_n11}), .b ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, new_AGEMA_signal_1630, SB_0_T1}), .c ({SubC_out_s3[64], SubC_out_s2[64], SubC_out_s1[64], SubC_out_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U5 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, SB_0_n15}), .b ({SubC_in_s3[32], SubC_in_s2[32], SubC_in_s1[32], SubC_in_s0[32]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, new_AGEMA_signal_2497, SB_0_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U4 ( .a ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, new_AGEMA_signal_1624, SB_0_n10}), .b ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, new_AGEMA_signal_1627, SB_0_T0}), .c ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, SB_0_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U1 ( .a ({SubC_in_s3[96], SubC_in_s2[96], SubC_in_s1[96], SubC_in_s0[96]}), .b ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, new_AGEMA_signal_1636, SB_0_T3}), .c ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, SB_0_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_0_t0_AND_U1 ( .a ({SubC_in_s3[96], SubC_in_s2[96], SubC_in_s1[96], SubC_in_s0[96]}), .b ({SubC_in_s3[64], SubC_in_s2[64], SubC_in_s1[64], SubC_in_s0[64]}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, new_AGEMA_signal_1627, SB_0_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_0_t1_AND_U1 ( .a ({SubC_in_s3[96], SubC_in_s2[96], SubC_in_s1[96], SubC_in_s0[96]}), .b ({SubC_in_s3[32], SubC_in_s2[32], SubC_in_s1[32], SubC_in_s0[32]}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, new_AGEMA_signal_1630, SB_0_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_0_t2_AND_U1 ( .a ({SubC_in_s3[96], SubC_in_s2[96], SubC_in_s1[96], SubC_in_s0[96]}), .b ({SubC_in_s3[0], SubC_in_s2[0], SubC_in_s1[0], SubC_in_s0[0]}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, SB_0_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_0_t3_AND_U1 ( .a ({SubC_in_s3[64], SubC_in_s2[64], SubC_in_s1[64], SubC_in_s0[64]}), .b ({SubC_in_s3[0], SubC_in_s2[0], SubC_in_s1[0], SubC_in_s0[0]}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, new_AGEMA_signal_1636, SB_0_T3}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U10 ( .a ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, new_AGEMA_signal_2122, SB_31_n13}), .b ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, new_AGEMA_signal_1639, SB_31_n12}), .c ({SubC_out_s3[63], SubC_out_s2[63], SubC_out_s1[63], SubC_out_s0[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U7 ( .a ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, new_AGEMA_signal_1648, SB_31_T4}), .b ({new_AGEMA_signal_708, new_AGEMA_signal_707, new_AGEMA_signal_706, SB_31_T3}), .c ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, new_AGEMA_signal_2122, SB_31_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_31_U2 ( .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, new_AGEMA_signal_1645, SB_31_n9}), .b ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, new_AGEMA_signal_1651, SB_31_T5}), .c ({SubC_out_s3[31], SubC_out_s2[31], SubC_out_s1[31], SubC_out_s0[31]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_31_t4_AND_U1 ( .a ({SubC_in_s3[63], SubC_in_s2[63], SubC_in_s1[63], SubC_in_s0[63]}), .b ({new_AGEMA_signal_708, new_AGEMA_signal_707, new_AGEMA_signal_706, SB_31_T3}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, new_AGEMA_signal_1648, SB_31_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_31_t5_AND_U1 ( .a ({SubC_in_s3[63], SubC_in_s2[63], SubC_in_s1[63], SubC_in_s0[63]}), .b ({new_AGEMA_signal_705, new_AGEMA_signal_704, new_AGEMA_signal_703, SB_31_T2}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, new_AGEMA_signal_1651, SB_31_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U10 ( .a ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, new_AGEMA_signal_2134, SB_30_n13}), .b ({new_AGEMA_signal_1656, new_AGEMA_signal_1655, new_AGEMA_signal_1654, SB_30_n12}), .c ({SubC_out_s3[62], SubC_out_s2[62], SubC_out_s1[62], SubC_out_s0[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U7 ( .a ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, new_AGEMA_signal_1663, SB_30_T4}), .b ({new_AGEMA_signal_738, new_AGEMA_signal_737, new_AGEMA_signal_736, SB_30_T3}), .c ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, new_AGEMA_signal_2134, SB_30_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_30_U2 ( .a ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, SB_30_n9}), .b ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, new_AGEMA_signal_1666, SB_30_T5}), .c ({SubC_out_s3[30], SubC_out_s2[30], SubC_out_s1[30], SubC_out_s0[30]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_30_t4_AND_U1 ( .a ({SubC_in_s3[62], SubC_in_s2[62], SubC_in_s1[62], SubC_in_s0[62]}), .b ({new_AGEMA_signal_738, new_AGEMA_signal_737, new_AGEMA_signal_736, SB_30_T3}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, new_AGEMA_signal_1663, SB_30_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_30_t5_AND_U1 ( .a ({SubC_in_s3[62], SubC_in_s2[62], SubC_in_s1[62], SubC_in_s0[62]}), .b ({new_AGEMA_signal_735, new_AGEMA_signal_734, new_AGEMA_signal_733, SB_30_T2}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, new_AGEMA_signal_1666, SB_30_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U10 ( .a ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, SB_29_n13}), .b ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, new_AGEMA_signal_1669, SB_29_n12}), .c ({SubC_out_s3[61], SubC_out_s2[61], SubC_out_s1[61], SubC_out_s0[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U7 ( .a ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, SB_29_T4}), .b ({new_AGEMA_signal_768, new_AGEMA_signal_767, new_AGEMA_signal_766, SB_29_T3}), .c ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, SB_29_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_29_U2 ( .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, new_AGEMA_signal_1675, SB_29_n9}), .b ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, new_AGEMA_signal_1681, SB_29_T5}), .c ({SubC_out_s3[29], SubC_out_s2[29], SubC_out_s1[29], SubC_out_s0[29]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_29_t4_AND_U1 ( .a ({SubC_in_s3[61], SubC_in_s2[61], SubC_in_s1[61], SubC_in_s0[61]}), .b ({new_AGEMA_signal_768, new_AGEMA_signal_767, new_AGEMA_signal_766, SB_29_T3}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, SB_29_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_29_t5_AND_U1 ( .a ({SubC_in_s3[61], SubC_in_s2[61], SubC_in_s1[61], SubC_in_s0[61]}), .b ({new_AGEMA_signal_765, new_AGEMA_signal_764, new_AGEMA_signal_763, SB_29_T2}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, new_AGEMA_signal_1681, SB_29_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U10 ( .a ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, SB_28_n13}), .b ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, new_AGEMA_signal_1684, SB_28_n12}), .c ({SubC_out_s3[60], SubC_out_s2[60], SubC_out_s1[60], SubC_out_s0[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U7 ( .a ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, new_AGEMA_signal_1693, SB_28_T4}), .b ({new_AGEMA_signal_798, new_AGEMA_signal_797, new_AGEMA_signal_796, SB_28_T3}), .c ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, SB_28_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_28_U2 ( .a ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, new_AGEMA_signal_1690, SB_28_n9}), .b ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, new_AGEMA_signal_1696, SB_28_T5}), .c ({SubC_out_s3[28], SubC_out_s2[28], SubC_out_s1[28], SubC_out_s0[28]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_28_t4_AND_U1 ( .a ({SubC_in_s3[60], SubC_in_s2[60], SubC_in_s1[60], SubC_in_s0[60]}), .b ({new_AGEMA_signal_798, new_AGEMA_signal_797, new_AGEMA_signal_796, SB_28_T3}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, new_AGEMA_signal_1693, SB_28_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_28_t5_AND_U1 ( .a ({SubC_in_s3[60], SubC_in_s2[60], SubC_in_s1[60], SubC_in_s0[60]}), .b ({new_AGEMA_signal_795, new_AGEMA_signal_794, new_AGEMA_signal_793, SB_28_T2}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, new_AGEMA_signal_1696, SB_28_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U10 ( .a ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, SB_27_n13}), .b ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, new_AGEMA_signal_1699, SB_27_n12}), .c ({SubC_out_s3[59], SubC_out_s2[59], SubC_out_s1[59], SubC_out_s0[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U7 ( .a ({new_AGEMA_signal_1710, new_AGEMA_signal_1709, new_AGEMA_signal_1708, SB_27_T4}), .b ({new_AGEMA_signal_828, new_AGEMA_signal_827, new_AGEMA_signal_826, SB_27_T3}), .c ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, SB_27_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_27_U2 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, new_AGEMA_signal_1705, SB_27_n9}), .b ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, new_AGEMA_signal_1711, SB_27_T5}), .c ({SubC_out_s3[27], SubC_out_s2[27], SubC_out_s1[27], SubC_out_s0[27]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_27_t4_AND_U1 ( .a ({SubC_in_s3[59], SubC_in_s2[59], SubC_in_s1[59], SubC_in_s0[59]}), .b ({new_AGEMA_signal_828, new_AGEMA_signal_827, new_AGEMA_signal_826, SB_27_T3}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_1710, new_AGEMA_signal_1709, new_AGEMA_signal_1708, SB_27_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_27_t5_AND_U1 ( .a ({SubC_in_s3[59], SubC_in_s2[59], SubC_in_s1[59], SubC_in_s0[59]}), .b ({new_AGEMA_signal_825, new_AGEMA_signal_824, new_AGEMA_signal_823, SB_27_T2}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, new_AGEMA_signal_1711, SB_27_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U10 ( .a ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, new_AGEMA_signal_2182, SB_26_n13}), .b ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, new_AGEMA_signal_1714, SB_26_n12}), .c ({SubC_out_s3[58], SubC_out_s2[58], SubC_out_s1[58], SubC_out_s0[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U7 ( .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, SB_26_T4}), .b ({new_AGEMA_signal_858, new_AGEMA_signal_857, new_AGEMA_signal_856, SB_26_T3}), .c ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, new_AGEMA_signal_2182, SB_26_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_26_U2 ( .a ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, new_AGEMA_signal_1720, SB_26_n9}), .b ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, new_AGEMA_signal_1726, SB_26_T5}), .c ({SubC_out_s3[26], SubC_out_s2[26], SubC_out_s1[26], SubC_out_s0[26]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_26_t4_AND_U1 ( .a ({SubC_in_s3[58], SubC_in_s2[58], SubC_in_s1[58], SubC_in_s0[58]}), .b ({new_AGEMA_signal_858, new_AGEMA_signal_857, new_AGEMA_signal_856, SB_26_T3}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, SB_26_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_26_t5_AND_U1 ( .a ({SubC_in_s3[58], SubC_in_s2[58], SubC_in_s1[58], SubC_in_s0[58]}), .b ({new_AGEMA_signal_855, new_AGEMA_signal_854, new_AGEMA_signal_853, SB_26_T2}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, new_AGEMA_signal_1726, SB_26_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U10 ( .a ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, SB_25_n13}), .b ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, new_AGEMA_signal_1729, SB_25_n12}), .c ({SubC_out_s3[57], SubC_out_s2[57], SubC_out_s1[57], SubC_out_s0[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U7 ( .a ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, new_AGEMA_signal_1738, SB_25_T4}), .b ({new_AGEMA_signal_888, new_AGEMA_signal_887, new_AGEMA_signal_886, SB_25_T3}), .c ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, new_AGEMA_signal_2194, SB_25_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_25_U2 ( .a ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, new_AGEMA_signal_1735, SB_25_n9}), .b ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, new_AGEMA_signal_1741, SB_25_T5}), .c ({SubC_out_s3[25], SubC_out_s2[25], SubC_out_s1[25], SubC_out_s0[25]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_25_t4_AND_U1 ( .a ({SubC_in_s3[57], SubC_in_s2[57], SubC_in_s1[57], SubC_in_s0[57]}), .b ({new_AGEMA_signal_888, new_AGEMA_signal_887, new_AGEMA_signal_886, SB_25_T3}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, new_AGEMA_signal_1738, SB_25_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_25_t5_AND_U1 ( .a ({SubC_in_s3[57], SubC_in_s2[57], SubC_in_s1[57], SubC_in_s0[57]}), .b ({new_AGEMA_signal_885, new_AGEMA_signal_884, new_AGEMA_signal_883, SB_25_T2}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, new_AGEMA_signal_1741, SB_25_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U10 ( .a ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, SB_24_n13}), .b ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, new_AGEMA_signal_1744, SB_24_n12}), .c ({SubC_out_s3[56], SubC_out_s2[56], SubC_out_s1[56], SubC_out_s0[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U7 ( .a ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, new_AGEMA_signal_1753, SB_24_T4}), .b ({new_AGEMA_signal_918, new_AGEMA_signal_917, new_AGEMA_signal_916, SB_24_T3}), .c ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, SB_24_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_24_U2 ( .a ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, SB_24_n9}), .b ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, new_AGEMA_signal_1756, SB_24_T5}), .c ({SubC_out_s3[24], SubC_out_s2[24], SubC_out_s1[24], SubC_out_s0[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_24_t4_AND_U1 ( .a ({SubC_in_s3[56], SubC_in_s2[56], SubC_in_s1[56], SubC_in_s0[56]}), .b ({new_AGEMA_signal_918, new_AGEMA_signal_917, new_AGEMA_signal_916, SB_24_T3}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, new_AGEMA_signal_1753, SB_24_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_24_t5_AND_U1 ( .a ({SubC_in_s3[56], SubC_in_s2[56], SubC_in_s1[56], SubC_in_s0[56]}), .b ({new_AGEMA_signal_915, new_AGEMA_signal_914, new_AGEMA_signal_913, SB_24_T2}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, new_AGEMA_signal_1756, SB_24_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U10 ( .a ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, SB_23_n13}), .b ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, new_AGEMA_signal_1759, SB_23_n12}), .c ({SubC_out_s3[55], SubC_out_s2[55], SubC_out_s1[55], SubC_out_s0[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U7 ( .a ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, new_AGEMA_signal_1768, SB_23_T4}), .b ({new_AGEMA_signal_948, new_AGEMA_signal_947, new_AGEMA_signal_946, SB_23_T3}), .c ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, SB_23_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_23_U2 ( .a ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, new_AGEMA_signal_1765, SB_23_n9}), .b ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, new_AGEMA_signal_1771, SB_23_T5}), .c ({SubC_out_s3[23], SubC_out_s2[23], SubC_out_s1[23], SubC_out_s0[23]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_23_t4_AND_U1 ( .a ({SubC_in_s3[55], SubC_in_s2[55], SubC_in_s1[55], SubC_in_s0[55]}), .b ({new_AGEMA_signal_948, new_AGEMA_signal_947, new_AGEMA_signal_946, SB_23_T3}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, new_AGEMA_signal_1768, SB_23_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_23_t5_AND_U1 ( .a ({SubC_in_s3[55], SubC_in_s2[55], SubC_in_s1[55], SubC_in_s0[55]}), .b ({new_AGEMA_signal_945, new_AGEMA_signal_944, new_AGEMA_signal_943, SB_23_T2}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, new_AGEMA_signal_1771, SB_23_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U10 ( .a ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, SB_22_n13}), .b ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, new_AGEMA_signal_1774, SB_22_n12}), .c ({SubC_out_s3[54], SubC_out_s2[54], SubC_out_s1[54], SubC_out_s0[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U7 ( .a ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, new_AGEMA_signal_1783, SB_22_T4}), .b ({new_AGEMA_signal_978, new_AGEMA_signal_977, new_AGEMA_signal_976, SB_22_T3}), .c ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, SB_22_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_22_U2 ( .a ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, new_AGEMA_signal_1780, SB_22_n9}), .b ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, SB_22_T5}), .c ({SubC_out_s3[22], SubC_out_s2[22], SubC_out_s1[22], SubC_out_s0[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_22_t4_AND_U1 ( .a ({SubC_in_s3[54], SubC_in_s2[54], SubC_in_s1[54], SubC_in_s0[54]}), .b ({new_AGEMA_signal_978, new_AGEMA_signal_977, new_AGEMA_signal_976, SB_22_T3}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, new_AGEMA_signal_1783, SB_22_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_22_t5_AND_U1 ( .a ({SubC_in_s3[54], SubC_in_s2[54], SubC_in_s1[54], SubC_in_s0[54]}), .b ({new_AGEMA_signal_975, new_AGEMA_signal_974, new_AGEMA_signal_973, SB_22_T2}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, SB_22_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U10 ( .a ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, SB_21_n13}), .b ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, new_AGEMA_signal_1789, SB_21_n12}), .c ({SubC_out_s3[53], SubC_out_s2[53], SubC_out_s1[53], SubC_out_s0[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U7 ( .a ({new_AGEMA_signal_1800, new_AGEMA_signal_1799, new_AGEMA_signal_1798, SB_21_T4}), .b ({new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, SB_21_T3}), .c ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, SB_21_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_21_U2 ( .a ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, SB_21_n9}), .b ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, new_AGEMA_signal_1801, SB_21_T5}), .c ({SubC_out_s3[21], SubC_out_s2[21], SubC_out_s1[21], SubC_out_s0[21]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_21_t4_AND_U1 ( .a ({SubC_in_s3[53], SubC_in_s2[53], SubC_in_s1[53], SubC_in_s0[53]}), .b ({new_AGEMA_signal_1008, new_AGEMA_signal_1007, new_AGEMA_signal_1006, SB_21_T3}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_1800, new_AGEMA_signal_1799, new_AGEMA_signal_1798, SB_21_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_21_t5_AND_U1 ( .a ({SubC_in_s3[53], SubC_in_s2[53], SubC_in_s1[53], SubC_in_s0[53]}), .b ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, new_AGEMA_signal_1003, SB_21_T2}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, new_AGEMA_signal_1801, SB_21_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U10 ( .a ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, SB_20_n13}), .b ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, new_AGEMA_signal_1804, SB_20_n12}), .c ({SubC_out_s3[52], SubC_out_s2[52], SubC_out_s1[52], SubC_out_s0[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U7 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, SB_20_T4}), .b ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, new_AGEMA_signal_1036, SB_20_T3}), .c ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, SB_20_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_20_U2 ( .a ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, new_AGEMA_signal_1810, SB_20_n9}), .b ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, new_AGEMA_signal_1816, SB_20_T5}), .c ({SubC_out_s3[20], SubC_out_s2[20], SubC_out_s1[20], SubC_out_s0[20]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_20_t4_AND_U1 ( .a ({SubC_in_s3[52], SubC_in_s2[52], SubC_in_s1[52], SubC_in_s0[52]}), .b ({new_AGEMA_signal_1038, new_AGEMA_signal_1037, new_AGEMA_signal_1036, SB_20_T3}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, SB_20_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_20_t5_AND_U1 ( .a ({SubC_in_s3[52], SubC_in_s2[52], SubC_in_s1[52], SubC_in_s0[52]}), .b ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, new_AGEMA_signal_1033, SB_20_T2}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, new_AGEMA_signal_1816, SB_20_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U10 ( .a ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, SB_19_n13}), .b ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, new_AGEMA_signal_1819, SB_19_n12}), .c ({SubC_out_s3[51], SubC_out_s2[51], SubC_out_s1[51], SubC_out_s0[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U7 ( .a ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, new_AGEMA_signal_1828, SB_19_T4}), .b ({new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, SB_19_T3}), .c ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, SB_19_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_19_U2 ( .a ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, new_AGEMA_signal_1825, SB_19_n9}), .b ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, new_AGEMA_signal_1831, SB_19_T5}), .c ({SubC_out_s3[19], SubC_out_s2[19], SubC_out_s1[19], SubC_out_s0[19]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_19_t4_AND_U1 ( .a ({SubC_in_s3[51], SubC_in_s2[51], SubC_in_s1[51], SubC_in_s0[51]}), .b ({new_AGEMA_signal_1068, new_AGEMA_signal_1067, new_AGEMA_signal_1066, SB_19_T3}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, new_AGEMA_signal_1828, SB_19_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_19_t5_AND_U1 ( .a ({SubC_in_s3[51], SubC_in_s2[51], SubC_in_s1[51], SubC_in_s0[51]}), .b ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, new_AGEMA_signal_1063, SB_19_T2}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, new_AGEMA_signal_1831, SB_19_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U10 ( .a ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, new_AGEMA_signal_2278, SB_18_n13}), .b ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, new_AGEMA_signal_1834, SB_18_n12}), .c ({SubC_out_s3[50], SubC_out_s2[50], SubC_out_s1[50], SubC_out_s0[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U7 ( .a ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, new_AGEMA_signal_1843, SB_18_T4}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, SB_18_T3}), .c ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, new_AGEMA_signal_2278, SB_18_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_18_U2 ( .a ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, SB_18_n9}), .b ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, new_AGEMA_signal_1846, SB_18_T5}), .c ({SubC_out_s3[18], SubC_out_s2[18], SubC_out_s1[18], SubC_out_s0[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_18_t4_AND_U1 ( .a ({SubC_in_s3[50], SubC_in_s2[50], SubC_in_s1[50], SubC_in_s0[50]}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, SB_18_T3}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, new_AGEMA_signal_1843, SB_18_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_18_t5_AND_U1 ( .a ({SubC_in_s3[50], SubC_in_s2[50], SubC_in_s1[50], SubC_in_s0[50]}), .b ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, new_AGEMA_signal_1093, SB_18_T2}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, new_AGEMA_signal_1846, SB_18_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U10 ( .a ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, SB_17_n13}), .b ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, new_AGEMA_signal_1849, SB_17_n12}), .c ({SubC_out_s3[49], SubC_out_s2[49], SubC_out_s1[49], SubC_out_s0[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U7 ( .a ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, SB_17_T4}), .b ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, SB_17_T3}), .c ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, SB_17_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_17_U2 ( .a ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, new_AGEMA_signal_1855, SB_17_n9}), .b ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, new_AGEMA_signal_1861, SB_17_T5}), .c ({SubC_out_s3[17], SubC_out_s2[17], SubC_out_s1[17], SubC_out_s0[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_17_t4_AND_U1 ( .a ({SubC_in_s3[49], SubC_in_s2[49], SubC_in_s1[49], SubC_in_s0[49]}), .b ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, SB_17_T3}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, SB_17_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_17_t5_AND_U1 ( .a ({SubC_in_s3[49], SubC_in_s2[49], SubC_in_s1[49], SubC_in_s0[49]}), .b ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, new_AGEMA_signal_1123, SB_17_T2}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, new_AGEMA_signal_1861, SB_17_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U10 ( .a ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, SB_16_n13}), .b ({new_AGEMA_signal_1866, new_AGEMA_signal_1865, new_AGEMA_signal_1864, SB_16_n12}), .c ({SubC_out_s3[48], SubC_out_s2[48], SubC_out_s1[48], SubC_out_s0[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U7 ( .a ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, new_AGEMA_signal_1873, SB_16_T4}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, SB_16_T3}), .c ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, SB_16_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_16_U2 ( .a ({new_AGEMA_signal_1872, new_AGEMA_signal_1871, new_AGEMA_signal_1870, SB_16_n9}), .b ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, new_AGEMA_signal_1876, SB_16_T5}), .c ({SubC_out_s3[16], SubC_out_s2[16], SubC_out_s1[16], SubC_out_s0[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_16_t4_AND_U1 ( .a ({SubC_in_s3[48], SubC_in_s2[48], SubC_in_s1[48], SubC_in_s0[48]}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, SB_16_T3}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, new_AGEMA_signal_1873, SB_16_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_16_t5_AND_U1 ( .a ({SubC_in_s3[48], SubC_in_s2[48], SubC_in_s1[48], SubC_in_s0[48]}), .b ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, new_AGEMA_signal_1153, SB_16_T2}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, new_AGEMA_signal_1876, SB_16_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U10 ( .a ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, SB_15_n13}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, new_AGEMA_signal_1879, SB_15_n12}), .c ({SubC_out_s3[47], SubC_out_s2[47], SubC_out_s1[47], SubC_out_s0[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U7 ( .a ({new_AGEMA_signal_1890, new_AGEMA_signal_1889, new_AGEMA_signal_1888, SB_15_T4}), .b ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, new_AGEMA_signal_1186, SB_15_T3}), .c ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, SB_15_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_15_U2 ( .a ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, new_AGEMA_signal_1885, SB_15_n9}), .b ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, new_AGEMA_signal_1891, SB_15_T5}), .c ({SubC_out_s3[15], SubC_out_s2[15], SubC_out_s1[15], SubC_out_s0[15]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_15_t4_AND_U1 ( .a ({SubC_in_s3[47], SubC_in_s2[47], SubC_in_s1[47], SubC_in_s0[47]}), .b ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, new_AGEMA_signal_1186, SB_15_T3}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_1890, new_AGEMA_signal_1889, new_AGEMA_signal_1888, SB_15_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_15_t5_AND_U1 ( .a ({SubC_in_s3[47], SubC_in_s2[47], SubC_in_s1[47], SubC_in_s0[47]}), .b ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, SB_15_T2}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, new_AGEMA_signal_1891, SB_15_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U10 ( .a ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, SB_14_n13}), .b ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, new_AGEMA_signal_1894, SB_14_n12}), .c ({SubC_out_s3[46], SubC_out_s2[46], SubC_out_s1[46], SubC_out_s0[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U7 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, SB_14_T4}), .b ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, new_AGEMA_signal_1216, SB_14_T3}), .c ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, SB_14_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_14_U2 ( .a ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, new_AGEMA_signal_1900, SB_14_n9}), .b ({new_AGEMA_signal_1908, new_AGEMA_signal_1907, new_AGEMA_signal_1906, SB_14_T5}), .c ({SubC_out_s3[14], SubC_out_s2[14], SubC_out_s1[14], SubC_out_s0[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_14_t4_AND_U1 ( .a ({SubC_in_s3[46], SubC_in_s2[46], SubC_in_s1[46], SubC_in_s0[46]}), .b ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, new_AGEMA_signal_1216, SB_14_T3}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, SB_14_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_14_t5_AND_U1 ( .a ({SubC_in_s3[46], SubC_in_s2[46], SubC_in_s1[46], SubC_in_s0[46]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, new_AGEMA_signal_1213, SB_14_T2}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_1908, new_AGEMA_signal_1907, new_AGEMA_signal_1906, SB_14_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U10 ( .a ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, SB_13_n13}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, new_AGEMA_signal_1909, SB_13_n12}), .c ({SubC_out_s3[45], SubC_out_s2[45], SubC_out_s1[45], SubC_out_s0[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U7 ( .a ({new_AGEMA_signal_1920, new_AGEMA_signal_1919, new_AGEMA_signal_1918, SB_13_T4}), .b ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, new_AGEMA_signal_1246, SB_13_T3}), .c ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, SB_13_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_13_U2 ( .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, new_AGEMA_signal_1915, SB_13_n9}), .b ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, new_AGEMA_signal_1921, SB_13_T5}), .c ({SubC_out_s3[13], SubC_out_s2[13], SubC_out_s1[13], SubC_out_s0[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_13_t4_AND_U1 ( .a ({SubC_in_s3[45], SubC_in_s2[45], SubC_in_s1[45], SubC_in_s0[45]}), .b ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, new_AGEMA_signal_1246, SB_13_T3}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_1920, new_AGEMA_signal_1919, new_AGEMA_signal_1918, SB_13_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_13_t5_AND_U1 ( .a ({SubC_in_s3[45], SubC_in_s2[45], SubC_in_s1[45], SubC_in_s0[45]}), .b ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, SB_13_T2}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, new_AGEMA_signal_1921, SB_13_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U10 ( .a ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, SB_12_n13}), .b ({new_AGEMA_signal_1926, new_AGEMA_signal_1925, new_AGEMA_signal_1924, SB_12_n12}), .c ({SubC_out_s3[44], SubC_out_s2[44], SubC_out_s1[44], SubC_out_s0[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U7 ( .a ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, new_AGEMA_signal_1933, SB_12_T4}), .b ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, new_AGEMA_signal_1276, SB_12_T3}), .c ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, SB_12_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_12_U2 ( .a ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, SB_12_n9}), .b ({new_AGEMA_signal_1938, new_AGEMA_signal_1937, new_AGEMA_signal_1936, SB_12_T5}), .c ({SubC_out_s3[12], SubC_out_s2[12], SubC_out_s1[12], SubC_out_s0[12]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_12_t4_AND_U1 ( .a ({SubC_in_s3[44], SubC_in_s2[44], SubC_in_s1[44], SubC_in_s0[44]}), .b ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, new_AGEMA_signal_1276, SB_12_T3}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, new_AGEMA_signal_1933, SB_12_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_12_t5_AND_U1 ( .a ({SubC_in_s3[44], SubC_in_s2[44], SubC_in_s1[44], SubC_in_s0[44]}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, new_AGEMA_signal_1273, SB_12_T2}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_1938, new_AGEMA_signal_1937, new_AGEMA_signal_1936, SB_12_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U10 ( .a ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, SB_11_n13}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, new_AGEMA_signal_1939, SB_11_n12}), .c ({SubC_out_s3[43], SubC_out_s2[43], SubC_out_s1[43], SubC_out_s0[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U7 ( .a ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, new_AGEMA_signal_1948, SB_11_T4}), .b ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, SB_11_T3}), .c ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, SB_11_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_11_U2 ( .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, new_AGEMA_signal_1945, SB_11_n9}), .b ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, new_AGEMA_signal_1951, SB_11_T5}), .c ({SubC_out_s3[11], SubC_out_s2[11], SubC_out_s1[11], SubC_out_s0[11]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_11_t4_AND_U1 ( .a ({SubC_in_s3[43], SubC_in_s2[43], SubC_in_s1[43], SubC_in_s0[43]}), .b ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, SB_11_T3}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, new_AGEMA_signal_1948, SB_11_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_11_t5_AND_U1 ( .a ({SubC_in_s3[43], SubC_in_s2[43], SubC_in_s1[43], SubC_in_s0[43]}), .b ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, new_AGEMA_signal_1303, SB_11_T2}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, new_AGEMA_signal_1951, SB_11_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U10 ( .a ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, SB_10_n13}), .b ({new_AGEMA_signal_1956, new_AGEMA_signal_1955, new_AGEMA_signal_1954, SB_10_n12}), .c ({SubC_out_s3[42], SubC_out_s2[42], SubC_out_s1[42], SubC_out_s0[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U7 ( .a ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, new_AGEMA_signal_1963, SB_10_T4}), .b ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, new_AGEMA_signal_1336, SB_10_T3}), .c ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, SB_10_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_10_U2 ( .a ({new_AGEMA_signal_1962, new_AGEMA_signal_1961, new_AGEMA_signal_1960, SB_10_n9}), .b ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, SB_10_T5}), .c ({SubC_out_s3[10], SubC_out_s2[10], SubC_out_s1[10], SubC_out_s0[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_10_t4_AND_U1 ( .a ({SubC_in_s3[42], SubC_in_s2[42], SubC_in_s1[42], SubC_in_s0[42]}), .b ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, new_AGEMA_signal_1336, SB_10_T3}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, new_AGEMA_signal_1963, SB_10_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_10_t5_AND_U1 ( .a ({SubC_in_s3[42], SubC_in_s2[42], SubC_in_s1[42], SubC_in_s0[42]}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, new_AGEMA_signal_1333, SB_10_T2}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, SB_10_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U10 ( .a ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, SB_9_n13}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, new_AGEMA_signal_1969, SB_9_n12}), .c ({SubC_out_s3[41], SubC_out_s2[41], SubC_out_s1[41], SubC_out_s0[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U7 ( .a ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, new_AGEMA_signal_1978, SB_9_T4}), .b ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, SB_9_T3}), .c ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, SB_9_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_9_U2 ( .a ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, SB_9_n9}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, new_AGEMA_signal_1981, SB_9_T5}), .c ({SubC_out_s3[9], SubC_out_s2[9], SubC_out_s1[9], SubC_out_s0[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_9_t4_AND_U1 ( .a ({SubC_in_s3[41], SubC_in_s2[41], SubC_in_s1[41], SubC_in_s0[41]}), .b ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, SB_9_T3}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, new_AGEMA_signal_1978, SB_9_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_9_t5_AND_U1 ( .a ({SubC_in_s3[41], SubC_in_s2[41], SubC_in_s1[41], SubC_in_s0[41]}), .b ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, new_AGEMA_signal_1363, SB_9_T2}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, new_AGEMA_signal_1981, SB_9_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U10 ( .a ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, SB_8_n13}), .b ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, new_AGEMA_signal_1984, SB_8_n12}), .c ({SubC_out_s3[40], SubC_out_s2[40], SubC_out_s1[40], SubC_out_s0[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U7 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, SB_8_T4}), .b ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, new_AGEMA_signal_1396, SB_8_T3}), .c ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, SB_8_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_8_U2 ( .a ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, new_AGEMA_signal_1990, SB_8_n9}), .b ({new_AGEMA_signal_1998, new_AGEMA_signal_1997, new_AGEMA_signal_1996, SB_8_T5}), .c ({SubC_out_s3[8], SubC_out_s2[8], SubC_out_s1[8], SubC_out_s0[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_8_t4_AND_U1 ( .a ({SubC_in_s3[40], SubC_in_s2[40], SubC_in_s1[40], SubC_in_s0[40]}), .b ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, new_AGEMA_signal_1396, SB_8_T3}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, SB_8_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_8_t5_AND_U1 ( .a ({SubC_in_s3[40], SubC_in_s2[40], SubC_in_s1[40], SubC_in_s0[40]}), .b ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, new_AGEMA_signal_1393, SB_8_T2}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_1998, new_AGEMA_signal_1997, new_AGEMA_signal_1996, SB_8_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U10 ( .a ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, SB_7_n13}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, new_AGEMA_signal_1999, SB_7_n12}), .c ({SubC_out_s3[39], SubC_out_s2[39], SubC_out_s1[39], SubC_out_s0[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U7 ( .a ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, new_AGEMA_signal_2008, SB_7_T4}), .b ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, SB_7_T3}), .c ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, SB_7_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_7_U2 ( .a ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, new_AGEMA_signal_2005, SB_7_n9}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, new_AGEMA_signal_2011, SB_7_T5}), .c ({SubC_out_s3[7], SubC_out_s2[7], SubC_out_s1[7], SubC_out_s0[7]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_7_t4_AND_U1 ( .a ({SubC_in_s3[39], SubC_in_s2[39], SubC_in_s1[39], SubC_in_s0[39]}), .b ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, SB_7_T3}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, new_AGEMA_signal_2008, SB_7_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_7_t5_AND_U1 ( .a ({SubC_in_s3[39], SubC_in_s2[39], SubC_in_s1[39], SubC_in_s0[39]}), .b ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, SB_7_T2}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, new_AGEMA_signal_2011, SB_7_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U10 ( .a ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, SB_6_n13}), .b ({new_AGEMA_signal_2016, new_AGEMA_signal_2015, new_AGEMA_signal_2014, SB_6_n12}), .c ({SubC_out_s3[38], SubC_out_s2[38], SubC_out_s1[38], SubC_out_s0[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U7 ( .a ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, new_AGEMA_signal_2023, SB_6_T4}), .b ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, new_AGEMA_signal_1456, SB_6_T3}), .c ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, SB_6_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_6_U2 ( .a ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, SB_6_n9}), .b ({new_AGEMA_signal_2028, new_AGEMA_signal_2027, new_AGEMA_signal_2026, SB_6_T5}), .c ({SubC_out_s3[6], SubC_out_s2[6], SubC_out_s1[6], SubC_out_s0[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_6_t4_AND_U1 ( .a ({SubC_in_s3[38], SubC_in_s2[38], SubC_in_s1[38], SubC_in_s0[38]}), .b ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, new_AGEMA_signal_1456, SB_6_T3}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, new_AGEMA_signal_2023, SB_6_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_6_t5_AND_U1 ( .a ({SubC_in_s3[38], SubC_in_s2[38], SubC_in_s1[38], SubC_in_s0[38]}), .b ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, new_AGEMA_signal_1453, SB_6_T2}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_2028, new_AGEMA_signal_2027, new_AGEMA_signal_2026, SB_6_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U10 ( .a ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, SB_5_n13}), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, new_AGEMA_signal_2029, SB_5_n12}), .c ({SubC_out_s3[37], SubC_out_s2[37], SubC_out_s1[37], SubC_out_s0[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U7 ( .a ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, SB_5_T4}), .b ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, new_AGEMA_signal_1486, SB_5_T3}), .c ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, SB_5_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_5_U2 ( .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, new_AGEMA_signal_2035, SB_5_n9}), .b ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, new_AGEMA_signal_2041, SB_5_T5}), .c ({SubC_out_s3[5], SubC_out_s2[5], SubC_out_s1[5], SubC_out_s0[5]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_5_t4_AND_U1 ( .a ({SubC_in_s3[37], SubC_in_s2[37], SubC_in_s1[37], SubC_in_s0[37]}), .b ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, new_AGEMA_signal_1486, SB_5_T3}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, SB_5_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_5_t5_AND_U1 ( .a ({SubC_in_s3[37], SubC_in_s2[37], SubC_in_s1[37], SubC_in_s0[37]}), .b ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, SB_5_T2}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, new_AGEMA_signal_2041, SB_5_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U10 ( .a ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, SB_4_n13}), .b ({new_AGEMA_signal_2046, new_AGEMA_signal_2045, new_AGEMA_signal_2044, SB_4_n12}), .c ({SubC_out_s3[36], SubC_out_s2[36], SubC_out_s1[36], SubC_out_s0[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U7 ( .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, new_AGEMA_signal_2053, SB_4_T4}), .b ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, SB_4_T3}), .c ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, SB_4_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_4_U2 ( .a ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, new_AGEMA_signal_2050, SB_4_n9}), .b ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, new_AGEMA_signal_2056, SB_4_T5}), .c ({SubC_out_s3[4], SubC_out_s2[4], SubC_out_s1[4], SubC_out_s0[4]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_4_t4_AND_U1 ( .a ({SubC_in_s3[36], SubC_in_s2[36], SubC_in_s1[36], SubC_in_s0[36]}), .b ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, SB_4_T3}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, new_AGEMA_signal_2053, SB_4_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_4_t5_AND_U1 ( .a ({SubC_in_s3[36], SubC_in_s2[36], SubC_in_s1[36], SubC_in_s0[36]}), .b ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, new_AGEMA_signal_1513, SB_4_T2}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, new_AGEMA_signal_2056, SB_4_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U10 ( .a ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, SB_3_n13}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, new_AGEMA_signal_2059, SB_3_n12}), .c ({SubC_out_s3[35], SubC_out_s2[35], SubC_out_s1[35], SubC_out_s0[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U7 ( .a ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, new_AGEMA_signal_2068, SB_3_T4}), .b ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, new_AGEMA_signal_1546, SB_3_T3}), .c ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, SB_3_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_3_U2 ( .a ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, new_AGEMA_signal_2065, SB_3_n9}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, new_AGEMA_signal_2071, SB_3_T5}), .c ({SubC_out_s3[3], SubC_out_s2[3], SubC_out_s1[3], SubC_out_s0[3]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_3_t4_AND_U1 ( .a ({SubC_in_s3[35], SubC_in_s2[35], SubC_in_s1[35], SubC_in_s0[35]}), .b ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, new_AGEMA_signal_1546, SB_3_T3}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, new_AGEMA_signal_2068, SB_3_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_3_t5_AND_U1 ( .a ({SubC_in_s3[35], SubC_in_s2[35], SubC_in_s1[35], SubC_in_s0[35]}), .b ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, SB_3_T2}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, new_AGEMA_signal_2071, SB_3_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U10 ( .a ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, SB_2_n13}), .b ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, new_AGEMA_signal_2074, SB_2_n12}), .c ({SubC_out_s3[34], SubC_out_s2[34], SubC_out_s1[34], SubC_out_s0[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U7 ( .a ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, SB_2_T4}), .b ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, new_AGEMA_signal_1576, SB_2_T3}), .c ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, SB_2_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_2_U2 ( .a ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, SB_2_n9}), .b ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, SB_2_T5}), .c ({SubC_out_s3[2], SubC_out_s2[2], SubC_out_s1[2], SubC_out_s0[2]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_2_t4_AND_U1 ( .a ({SubC_in_s3[34], SubC_in_s2[34], SubC_in_s1[34], SubC_in_s0[34]}), .b ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, new_AGEMA_signal_1576, SB_2_T3}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, SB_2_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_2_t5_AND_U1 ( .a ({SubC_in_s3[34], SubC_in_s2[34], SubC_in_s1[34], SubC_in_s0[34]}), .b ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, new_AGEMA_signal_1573, SB_2_T2}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, SB_2_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U10 ( .a ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, SB_1_n13}), .b ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, new_AGEMA_signal_2089, SB_1_n12}), .c ({SubC_out_s3[33], SubC_out_s2[33], SubC_out_s1[33], SubC_out_s0[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U7 ( .a ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, SB_1_T4}), .b ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, SB_1_T3}), .c ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, SB_1_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_1_U2 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, SB_1_n9}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, new_AGEMA_signal_2101, SB_1_T5}), .c ({SubC_out_s3[1], SubC_out_s2[1], SubC_out_s1[1], SubC_out_s0[1]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_1_t4_AND_U1 ( .a ({SubC_in_s3[33], SubC_in_s2[33], SubC_in_s1[33], SubC_in_s0[33]}), .b ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, SB_1_T3}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, SB_1_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_1_t5_AND_U1 ( .a ({SubC_in_s3[33], SubC_in_s2[33], SubC_in_s1[33], SubC_in_s0[33]}), .b ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, new_AGEMA_signal_1603, SB_1_T2}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, new_AGEMA_signal_2101, SB_1_T5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U10 ( .a ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, SB_0_n13}), .b ({new_AGEMA_signal_2106, new_AGEMA_signal_2105, new_AGEMA_signal_2104, SB_0_n12}), .c ({SubC_out_s3[32], SubC_out_s2[32], SubC_out_s1[32], SubC_out_s0[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U7 ( .a ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, SB_0_T4}), .b ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, new_AGEMA_signal_1636, SB_0_T3}), .c ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, SB_0_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SB_0_U2 ( .a ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, SB_0_n9}), .b ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, new_AGEMA_signal_2116, SB_0_T5}), .c ({SubC_out_s3[0], SubC_out_s2[0], SubC_out_s1[0], SubC_out_s0[0]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_0_t4_AND_U1 ( .a ({SubC_in_s3[32], SubC_in_s2[32], SubC_in_s1[32], SubC_in_s0[32]}), .b ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, new_AGEMA_signal_1636, SB_0_T3}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, SB_0_T4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SB_0_t5_AND_U1 ( .a ({SubC_in_s3[32], SubC_in_s2[32], SubC_in_s1[32], SubC_in_s0[32]}), .b ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, SB_0_T2}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, new_AGEMA_signal_2116, SB_0_T5}) ) ;

endmodule
