/* modified netlist. Source: module arx_round in file ./test/arx_round.v */
/* clock gating is added to the circuit, the latency increased 10 time(s)  */

module arx_round_HPC2_ClockGating_d2 (round_constant, round, x_round_in_s0, y_round_in_s0, clk, y_round_in_s1, y_round_in_s2, x_round_in_s1, x_round_in_s2, Fresh, /*rst,*/ x_round_out_s0, y_round_out_s0, x_round_out_s1, x_round_out_s2, y_round_out_s1, y_round_out_s2/*, Synch*/);
    input [31:0] round_constant ;
    input [1:0] round ;
    input [31:0] x_round_in_s0 ;
    input [31:0] y_round_in_s0 ;
    input clk ;
    input [31:0] y_round_in_s1 ;
    input [31:0] y_round_in_s2 ;
    input [31:0] x_round_in_s1 ;
    input [31:0] x_round_in_s2 ;
    //input rst ;
    input [767:0] Fresh ;
    output [31:0] x_round_out_s0 ;
    output [31:0] y_round_out_s0 ;
    output [31:0] x_round_out_s1 ;
    output [31:0] x_round_out_s2 ;
    output [31:0] y_round_out_s1 ;
    output [31:0] y_round_out_s2 ;
    //output Synch ;
    wire AdderIns_s2_gc_0_a1_t ;
    wire AdderIns_s2_bc_0_a1_t ;
    wire AdderIns_s2_bc_1_a1_t ;
    wire AdderIns_s2_bc_2_a1_t ;
    wire AdderIns_s2_bc_3_a1_t ;
    wire AdderIns_s2_bc_4_a1_t ;
    wire AdderIns_s2_bc_5_a1_t ;
    wire AdderIns_s2_bc_6_a1_t ;
    wire AdderIns_s2_bc_7_a1_t ;
    wire AdderIns_s2_bc_8_a1_t ;
    wire AdderIns_s2_bc_9_a1_t ;
    wire AdderIns_s2_bc_10_a1_t ;
    wire AdderIns_s2_bc_11_a1_t ;
    wire AdderIns_s2_bc_12_a1_t ;
    wire AdderIns_s2_bc_13_a1_t ;
    wire AdderIns_s2_bc_14_a1_t ;
    wire AdderIns_s2_bc_15_a1_t ;
    wire AdderIns_s2_bc_16_a1_t ;
    wire AdderIns_s2_bc_17_a1_t ;
    wire AdderIns_s2_bc_18_a1_t ;
    wire AdderIns_s2_bc_19_a1_t ;
    wire AdderIns_s2_bc_20_a1_t ;
    wire AdderIns_s2_bc_21_a1_t ;
    wire AdderIns_s2_bc_22_a1_t ;
    wire AdderIns_s2_bc_23_a1_t ;
    wire AdderIns_s2_bc_24_a1_t ;
    wire AdderIns_s2_bc_25_a1_t ;
    wire AdderIns_s2_bc_26_a1_t ;
    wire AdderIns_s2_bc_27_a1_t ;
    wire AdderIns_s2_bc_28_a1_t ;
    wire AdderIns_s2_bc_29_a1_t ;
    wire AdderIns_s3_gc_0_a1_t ;
    wire AdderIns_s3_gc_1_a1_t ;
    wire AdderIns_s3_bc_0_a1_t ;
    wire AdderIns_s3_bc_1_a1_t ;
    wire AdderIns_s3_bc_2_a1_t ;
    wire AdderIns_s3_bc_3_a1_t ;
    wire AdderIns_s3_bc_4_a1_t ;
    wire AdderIns_s3_bc_5_a1_t ;
    wire AdderIns_s3_bc_6_a1_t ;
    wire AdderIns_s3_bc_7_a1_t ;
    wire AdderIns_s3_bc_8_a1_t ;
    wire AdderIns_s3_bc_9_a1_t ;
    wire AdderIns_s3_bc_10_a1_t ;
    wire AdderIns_s3_bc_11_a1_t ;
    wire AdderIns_s3_bc_12_a1_t ;
    wire AdderIns_s3_bc_13_a1_t ;
    wire AdderIns_s3_bc_14_a1_t ;
    wire AdderIns_s3_bc_15_a1_t ;
    wire AdderIns_s3_bc_16_a1_t ;
    wire AdderIns_s3_bc_17_a1_t ;
    wire AdderIns_s3_bc_18_a1_t ;
    wire AdderIns_s3_bc_19_a1_t ;
    wire AdderIns_s3_bc_20_a1_t ;
    wire AdderIns_s3_bc_21_a1_t ;
    wire AdderIns_s3_bc_22_a1_t ;
    wire AdderIns_s3_bc_23_a1_t ;
    wire AdderIns_s3_bc_24_a1_t ;
    wire AdderIns_s3_bc_25_a1_t ;
    wire AdderIns_s3_bc_26_a1_t ;
    wire AdderIns_s3_bc_27_a1_t ;
    wire AdderIns_s4_gc_0_a1_t ;
    wire AdderIns_s4_gc_1_a1_t ;
    wire AdderIns_s4_gc_2_a1_t ;
    wire AdderIns_s4_gc_3_a1_t ;
    wire AdderIns_s4_bc_0_a1_t ;
    wire AdderIns_s4_bc_1_a1_t ;
    wire AdderIns_s4_bc_2_a1_t ;
    wire AdderIns_s4_bc_3_a1_t ;
    wire AdderIns_s4_bc_4_a1_t ;
    wire AdderIns_s4_bc_5_a1_t ;
    wire AdderIns_s4_bc_6_a1_t ;
    wire AdderIns_s4_bc_7_a1_t ;
    wire AdderIns_s4_bc_8_a1_t ;
    wire AdderIns_s4_bc_9_a1_t ;
    wire AdderIns_s4_bc_10_a1_t ;
    wire AdderIns_s4_bc_11_a1_t ;
    wire AdderIns_s4_bc_12_a1_t ;
    wire AdderIns_s4_bc_13_a1_t ;
    wire AdderIns_s4_bc_14_a1_t ;
    wire AdderIns_s4_bc_15_a1_t ;
    wire AdderIns_s4_bc_16_a1_t ;
    wire AdderIns_s4_bc_17_a1_t ;
    wire AdderIns_s4_bc_18_a1_t ;
    wire AdderIns_s4_bc_19_a1_t ;
    wire AdderIns_s4_bc_20_a1_t ;
    wire AdderIns_s4_bc_21_a1_t ;
    wire AdderIns_s4_bc_22_a1_t ;
    wire AdderIns_s4_bc_23_a1_t ;
    wire AdderIns_s5_gc_0_a1_t ;
    wire AdderIns_s5_gc_1_a1_t ;
    wire AdderIns_s5_gc_2_a1_t ;
    wire AdderIns_s5_gc_3_a1_t ;
    wire AdderIns_s5_gc_4_a1_t ;
    wire AdderIns_s5_gc_5_a1_t ;
    wire AdderIns_s5_gc_6_a1_t ;
    wire AdderIns_s5_gc_7_a1_t ;
    wire AdderIns_s5_bc_0_a1_t ;
    wire AdderIns_s5_bc_1_a1_t ;
    wire AdderIns_s5_bc_2_a1_t ;
    wire AdderIns_s5_bc_3_a1_t ;
    wire AdderIns_s5_bc_4_a1_t ;
    wire AdderIns_s5_bc_5_a1_t ;
    wire AdderIns_s5_bc_6_a1_t ;
    wire AdderIns_s5_bc_7_a1_t ;
    wire AdderIns_s5_bc_8_a1_t ;
    wire AdderIns_s5_bc_9_a1_t ;
    wire AdderIns_s5_bc_10_a1_t ;
    wire AdderIns_s5_bc_11_a1_t ;
    wire AdderIns_s5_bc_12_a1_t ;
    wire AdderIns_s5_bc_13_a1_t ;
    wire AdderIns_s5_bc_14_a1_t ;
    wire AdderIns_s5_bc_15_a1_t ;
    wire AdderIns_s6_gc_1_a1_t ;
    wire AdderIns_s6_gc_2_a1_t ;
    wire AdderIns_s6_gc_3_a1_t ;
    wire AdderIns_s6_gc_4_a1_t ;
    wire AdderIns_s6_gc_5_a1_t ;
    wire AdderIns_s6_gc_6_a1_t ;
    wire AdderIns_s6_gc_7_a1_t ;
    wire AdderIns_s6_gc_8_a1_t ;
    wire AdderIns_s6_gc_9_a1_t ;
    wire AdderIns_s6_gc_10_a1_t ;
    wire AdderIns_s6_gc_11_a1_t ;
    wire AdderIns_s6_gc_12_a1_t ;
    wire AdderIns_s6_gc_13_a1_t ;
    wire AdderIns_s6_gc_14_a1_t ;
    wire AdderIns_s6_gc_15_a1_t ;
    wire [31:0] y_rotated01 ;
    wire [31:0] y_rotated23 ;
    wire [31:0] y_rotated ;
    wire [31:0] sum ;
    wire [31:0] sum_rotated01 ;
    wire [31:0] sum_rotated23 ;
    wire [31:0] sum_rotated ;
    wire [30:0] AdderIns_g6 ;
    wire [31:1] AdderIns_p6 ;
    wire [30:16] AdderIns_g5 ;
    wire [15:1] AdderIns_p5 ;
    wire [30:7] AdderIns_g4 ;
    wire [23:0] AdderIns_p4 ;
    wire [30:3] AdderIns_g3 ;
    wire [27:0] AdderIns_p3 ;
    wire [30:1] AdderIns_g2 ;
    wire [29:0] AdderIns_p2 ;
    wire [30:0] AdderIns_g1 ;
    wire new_AGEMA_signal_828 ;
    wire new_AGEMA_signal_829 ;
    wire new_AGEMA_signal_834 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_840 ;
    wire new_AGEMA_signal_841 ;
    wire new_AGEMA_signal_846 ;
    wire new_AGEMA_signal_847 ;
    wire new_AGEMA_signal_852 ;
    wire new_AGEMA_signal_853 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_859 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_870 ;
    wire new_AGEMA_signal_871 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_900 ;
    wire new_AGEMA_signal_901 ;
    wire new_AGEMA_signal_906 ;
    wire new_AGEMA_signal_907 ;
    wire new_AGEMA_signal_910 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_915 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_919 ;
    wire new_AGEMA_signal_922 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_924 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_928 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_930 ;
    wire new_AGEMA_signal_931 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_934 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_939 ;
    wire new_AGEMA_signal_940 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_942 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) U129 ( .a ({1'b0, 1'b0, round_constant[0]}), .b ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, sum[0]}), .c ({x_round_out_s2[0], x_round_out_s1[0], x_round_out_s0[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_0_U1 ( .s (round[0]), .b ({y_round_in_s2[31], y_round_in_s1[31], y_round_in_s0[31]}), .a ({y_round_in_s2[17], y_round_in_s1[17], y_round_in_s0[17]}), .c ({new_AGEMA_signal_829, new_AGEMA_signal_828, y_rotated01[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_1_U1 ( .s (round[0]), .b ({y_round_in_s2[0], y_round_in_s1[0], y_round_in_s0[0]}), .a ({y_round_in_s2[18], y_round_in_s1[18], y_round_in_s0[18]}), .c ({new_AGEMA_signal_835, new_AGEMA_signal_834, y_rotated01[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_2_U1 ( .s (round[0]), .b ({y_round_in_s2[1], y_round_in_s1[1], y_round_in_s0[1]}), .a ({y_round_in_s2[19], y_round_in_s1[19], y_round_in_s0[19]}), .c ({new_AGEMA_signal_841, new_AGEMA_signal_840, y_rotated01[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_3_U1 ( .s (round[0]), .b ({y_round_in_s2[2], y_round_in_s1[2], y_round_in_s0[2]}), .a ({y_round_in_s2[20], y_round_in_s1[20], y_round_in_s0[20]}), .c ({new_AGEMA_signal_847, new_AGEMA_signal_846, y_rotated01[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_4_U1 ( .s (round[0]), .b ({y_round_in_s2[3], y_round_in_s1[3], y_round_in_s0[3]}), .a ({y_round_in_s2[21], y_round_in_s1[21], y_round_in_s0[21]}), .c ({new_AGEMA_signal_853, new_AGEMA_signal_852, y_rotated01[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_5_U1 ( .s (round[0]), .b ({y_round_in_s2[4], y_round_in_s1[4], y_round_in_s0[4]}), .a ({y_round_in_s2[22], y_round_in_s1[22], y_round_in_s0[22]}), .c ({new_AGEMA_signal_859, new_AGEMA_signal_858, y_rotated01[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_6_U1 ( .s (round[0]), .b ({y_round_in_s2[5], y_round_in_s1[5], y_round_in_s0[5]}), .a ({y_round_in_s2[23], y_round_in_s1[23], y_round_in_s0[23]}), .c ({new_AGEMA_signal_865, new_AGEMA_signal_864, y_rotated01[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_7_U1 ( .s (round[0]), .b ({y_round_in_s2[6], y_round_in_s1[6], y_round_in_s0[6]}), .a ({y_round_in_s2[24], y_round_in_s1[24], y_round_in_s0[24]}), .c ({new_AGEMA_signal_871, new_AGEMA_signal_870, y_rotated01[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_8_U1 ( .s (round[0]), .b ({y_round_in_s2[7], y_round_in_s1[7], y_round_in_s0[7]}), .a ({y_round_in_s2[25], y_round_in_s1[25], y_round_in_s0[25]}), .c ({new_AGEMA_signal_877, new_AGEMA_signal_876, y_rotated01[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_9_U1 ( .s (round[0]), .b ({y_round_in_s2[8], y_round_in_s1[8], y_round_in_s0[8]}), .a ({y_round_in_s2[26], y_round_in_s1[26], y_round_in_s0[26]}), .c ({new_AGEMA_signal_883, new_AGEMA_signal_882, y_rotated01[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_10_U1 ( .s (round[0]), .b ({y_round_in_s2[9], y_round_in_s1[9], y_round_in_s0[9]}), .a ({y_round_in_s2[27], y_round_in_s1[27], y_round_in_s0[27]}), .c ({new_AGEMA_signal_889, new_AGEMA_signal_888, y_rotated01[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_11_U1 ( .s (round[0]), .b ({y_round_in_s2[10], y_round_in_s1[10], y_round_in_s0[10]}), .a ({y_round_in_s2[28], y_round_in_s1[28], y_round_in_s0[28]}), .c ({new_AGEMA_signal_895, new_AGEMA_signal_894, y_rotated01[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_12_U1 ( .s (round[0]), .b ({y_round_in_s2[11], y_round_in_s1[11], y_round_in_s0[11]}), .a ({y_round_in_s2[29], y_round_in_s1[29], y_round_in_s0[29]}), .c ({new_AGEMA_signal_901, new_AGEMA_signal_900, y_rotated01[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_13_U1 ( .s (round[0]), .b ({y_round_in_s2[12], y_round_in_s1[12], y_round_in_s0[12]}), .a ({y_round_in_s2[30], y_round_in_s1[30], y_round_in_s0[30]}), .c ({new_AGEMA_signal_907, new_AGEMA_signal_906, y_rotated01[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_14_U1 ( .s (round[0]), .b ({y_round_in_s2[13], y_round_in_s1[13], y_round_in_s0[13]}), .a ({y_round_in_s2[31], y_round_in_s1[31], y_round_in_s0[31]}), .c ({new_AGEMA_signal_911, new_AGEMA_signal_910, y_rotated01[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_15_U1 ( .s (round[0]), .b ({y_round_in_s2[14], y_round_in_s1[14], y_round_in_s0[14]}), .a ({y_round_in_s2[0], y_round_in_s1[0], y_round_in_s0[0]}), .c ({new_AGEMA_signal_915, new_AGEMA_signal_914, y_rotated01[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_16_U1 ( .s (round[0]), .b ({y_round_in_s2[15], y_round_in_s1[15], y_round_in_s0[15]}), .a ({y_round_in_s2[1], y_round_in_s1[1], y_round_in_s0[1]}), .c ({new_AGEMA_signal_919, new_AGEMA_signal_918, y_rotated01[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_17_U1 ( .s (round[0]), .b ({y_round_in_s2[16], y_round_in_s1[16], y_round_in_s0[16]}), .a ({y_round_in_s2[2], y_round_in_s1[2], y_round_in_s0[2]}), .c ({new_AGEMA_signal_923, new_AGEMA_signal_922, y_rotated01[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_18_U1 ( .s (round[0]), .b ({y_round_in_s2[17], y_round_in_s1[17], y_round_in_s0[17]}), .a ({y_round_in_s2[3], y_round_in_s1[3], y_round_in_s0[3]}), .c ({new_AGEMA_signal_925, new_AGEMA_signal_924, y_rotated01[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_19_U1 ( .s (round[0]), .b ({y_round_in_s2[18], y_round_in_s1[18], y_round_in_s0[18]}), .a ({y_round_in_s2[4], y_round_in_s1[4], y_round_in_s0[4]}), .c ({new_AGEMA_signal_927, new_AGEMA_signal_926, y_rotated01[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_20_U1 ( .s (round[0]), .b ({y_round_in_s2[19], y_round_in_s1[19], y_round_in_s0[19]}), .a ({y_round_in_s2[5], y_round_in_s1[5], y_round_in_s0[5]}), .c ({new_AGEMA_signal_929, new_AGEMA_signal_928, y_rotated01[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_21_U1 ( .s (round[0]), .b ({y_round_in_s2[20], y_round_in_s1[20], y_round_in_s0[20]}), .a ({y_round_in_s2[6], y_round_in_s1[6], y_round_in_s0[6]}), .c ({new_AGEMA_signal_931, new_AGEMA_signal_930, y_rotated01[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_22_U1 ( .s (round[0]), .b ({y_round_in_s2[21], y_round_in_s1[21], y_round_in_s0[21]}), .a ({y_round_in_s2[7], y_round_in_s1[7], y_round_in_s0[7]}), .c ({new_AGEMA_signal_933, new_AGEMA_signal_932, y_rotated01[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_23_U1 ( .s (round[0]), .b ({y_round_in_s2[22], y_round_in_s1[22], y_round_in_s0[22]}), .a ({y_round_in_s2[8], y_round_in_s1[8], y_round_in_s0[8]}), .c ({new_AGEMA_signal_935, new_AGEMA_signal_934, y_rotated01[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_24_U1 ( .s (round[0]), .b ({y_round_in_s2[23], y_round_in_s1[23], y_round_in_s0[23]}), .a ({y_round_in_s2[9], y_round_in_s1[9], y_round_in_s0[9]}), .c ({new_AGEMA_signal_937, new_AGEMA_signal_936, y_rotated01[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_25_U1 ( .s (round[0]), .b ({y_round_in_s2[24], y_round_in_s1[24], y_round_in_s0[24]}), .a ({y_round_in_s2[10], y_round_in_s1[10], y_round_in_s0[10]}), .c ({new_AGEMA_signal_939, new_AGEMA_signal_938, y_rotated01[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_26_U1 ( .s (round[0]), .b ({y_round_in_s2[25], y_round_in_s1[25], y_round_in_s0[25]}), .a ({y_round_in_s2[11], y_round_in_s1[11], y_round_in_s0[11]}), .c ({new_AGEMA_signal_941, new_AGEMA_signal_940, y_rotated01[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_27_U1 ( .s (round[0]), .b ({y_round_in_s2[26], y_round_in_s1[26], y_round_in_s0[26]}), .a ({y_round_in_s2[12], y_round_in_s1[12], y_round_in_s0[12]}), .c ({new_AGEMA_signal_943, new_AGEMA_signal_942, y_rotated01[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_28_U1 ( .s (round[0]), .b ({y_round_in_s2[27], y_round_in_s1[27], y_round_in_s0[27]}), .a ({y_round_in_s2[13], y_round_in_s1[13], y_round_in_s0[13]}), .c ({new_AGEMA_signal_945, new_AGEMA_signal_944, y_rotated01[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_29_U1 ( .s (round[0]), .b ({y_round_in_s2[28], y_round_in_s1[28], y_round_in_s0[28]}), .a ({y_round_in_s2[14], y_round_in_s1[14], y_round_in_s0[14]}), .c ({new_AGEMA_signal_947, new_AGEMA_signal_946, y_rotated01[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_30_U1 ( .s (round[0]), .b ({y_round_in_s2[29], y_round_in_s1[29], y_round_in_s0[29]}), .a ({y_round_in_s2[15], y_round_in_s1[15], y_round_in_s0[15]}), .c ({new_AGEMA_signal_949, new_AGEMA_signal_948, y_rotated01[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M0_mux_inst_31_U1 ( .s (round[0]), .b ({y_round_in_s2[30], y_round_in_s1[30], y_round_in_s0[30]}), .a ({y_round_in_s2[16], y_round_in_s1[16], y_round_in_s0[16]}), .c ({new_AGEMA_signal_951, new_AGEMA_signal_950, y_rotated01[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_0_U1 ( .s (round[0]), .b ({y_round_in_s2[0], y_round_in_s1[0], y_round_in_s0[0]}), .a ({y_round_in_s2[24], y_round_in_s1[24], y_round_in_s0[24]}), .c ({new_AGEMA_signal_953, new_AGEMA_signal_952, y_rotated23[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_1_U1 ( .s (round[0]), .b ({y_round_in_s2[1], y_round_in_s1[1], y_round_in_s0[1]}), .a ({y_round_in_s2[25], y_round_in_s1[25], y_round_in_s0[25]}), .c ({new_AGEMA_signal_955, new_AGEMA_signal_954, y_rotated23[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_2_U1 ( .s (round[0]), .b ({y_round_in_s2[2], y_round_in_s1[2], y_round_in_s0[2]}), .a ({y_round_in_s2[26], y_round_in_s1[26], y_round_in_s0[26]}), .c ({new_AGEMA_signal_957, new_AGEMA_signal_956, y_rotated23[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_3_U1 ( .s (round[0]), .b ({y_round_in_s2[3], y_round_in_s1[3], y_round_in_s0[3]}), .a ({y_round_in_s2[27], y_round_in_s1[27], y_round_in_s0[27]}), .c ({new_AGEMA_signal_959, new_AGEMA_signal_958, y_rotated23[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_4_U1 ( .s (round[0]), .b ({y_round_in_s2[4], y_round_in_s1[4], y_round_in_s0[4]}), .a ({y_round_in_s2[28], y_round_in_s1[28], y_round_in_s0[28]}), .c ({new_AGEMA_signal_961, new_AGEMA_signal_960, y_rotated23[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_5_U1 ( .s (round[0]), .b ({y_round_in_s2[5], y_round_in_s1[5], y_round_in_s0[5]}), .a ({y_round_in_s2[29], y_round_in_s1[29], y_round_in_s0[29]}), .c ({new_AGEMA_signal_963, new_AGEMA_signal_962, y_rotated23[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_6_U1 ( .s (round[0]), .b ({y_round_in_s2[6], y_round_in_s1[6], y_round_in_s0[6]}), .a ({y_round_in_s2[30], y_round_in_s1[30], y_round_in_s0[30]}), .c ({new_AGEMA_signal_965, new_AGEMA_signal_964, y_rotated23[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_7_U1 ( .s (round[0]), .b ({y_round_in_s2[7], y_round_in_s1[7], y_round_in_s0[7]}), .a ({y_round_in_s2[31], y_round_in_s1[31], y_round_in_s0[31]}), .c ({new_AGEMA_signal_967, new_AGEMA_signal_966, y_rotated23[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_8_U1 ( .s (round[0]), .b ({y_round_in_s2[8], y_round_in_s1[8], y_round_in_s0[8]}), .a ({y_round_in_s2[0], y_round_in_s1[0], y_round_in_s0[0]}), .c ({new_AGEMA_signal_969, new_AGEMA_signal_968, y_rotated23[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_9_U1 ( .s (round[0]), .b ({y_round_in_s2[9], y_round_in_s1[9], y_round_in_s0[9]}), .a ({y_round_in_s2[1], y_round_in_s1[1], y_round_in_s0[1]}), .c ({new_AGEMA_signal_971, new_AGEMA_signal_970, y_rotated23[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_10_U1 ( .s (round[0]), .b ({y_round_in_s2[10], y_round_in_s1[10], y_round_in_s0[10]}), .a ({y_round_in_s2[2], y_round_in_s1[2], y_round_in_s0[2]}), .c ({new_AGEMA_signal_973, new_AGEMA_signal_972, y_rotated23[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_11_U1 ( .s (round[0]), .b ({y_round_in_s2[11], y_round_in_s1[11], y_round_in_s0[11]}), .a ({y_round_in_s2[3], y_round_in_s1[3], y_round_in_s0[3]}), .c ({new_AGEMA_signal_975, new_AGEMA_signal_974, y_rotated23[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_12_U1 ( .s (round[0]), .b ({y_round_in_s2[12], y_round_in_s1[12], y_round_in_s0[12]}), .a ({y_round_in_s2[4], y_round_in_s1[4], y_round_in_s0[4]}), .c ({new_AGEMA_signal_977, new_AGEMA_signal_976, y_rotated23[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_13_U1 ( .s (round[0]), .b ({y_round_in_s2[13], y_round_in_s1[13], y_round_in_s0[13]}), .a ({y_round_in_s2[5], y_round_in_s1[5], y_round_in_s0[5]}), .c ({new_AGEMA_signal_979, new_AGEMA_signal_978, y_rotated23[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_14_U1 ( .s (round[0]), .b ({y_round_in_s2[14], y_round_in_s1[14], y_round_in_s0[14]}), .a ({y_round_in_s2[6], y_round_in_s1[6], y_round_in_s0[6]}), .c ({new_AGEMA_signal_981, new_AGEMA_signal_980, y_rotated23[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_15_U1 ( .s (round[0]), .b ({y_round_in_s2[15], y_round_in_s1[15], y_round_in_s0[15]}), .a ({y_round_in_s2[7], y_round_in_s1[7], y_round_in_s0[7]}), .c ({new_AGEMA_signal_983, new_AGEMA_signal_982, y_rotated23[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_16_U1 ( .s (round[0]), .b ({y_round_in_s2[16], y_round_in_s1[16], y_round_in_s0[16]}), .a ({y_round_in_s2[8], y_round_in_s1[8], y_round_in_s0[8]}), .c ({new_AGEMA_signal_985, new_AGEMA_signal_984, y_rotated23[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_17_U1 ( .s (round[0]), .b ({y_round_in_s2[17], y_round_in_s1[17], y_round_in_s0[17]}), .a ({y_round_in_s2[9], y_round_in_s1[9], y_round_in_s0[9]}), .c ({new_AGEMA_signal_987, new_AGEMA_signal_986, y_rotated23[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_18_U1 ( .s (round[0]), .b ({y_round_in_s2[18], y_round_in_s1[18], y_round_in_s0[18]}), .a ({y_round_in_s2[10], y_round_in_s1[10], y_round_in_s0[10]}), .c ({new_AGEMA_signal_989, new_AGEMA_signal_988, y_rotated23[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_19_U1 ( .s (round[0]), .b ({y_round_in_s2[19], y_round_in_s1[19], y_round_in_s0[19]}), .a ({y_round_in_s2[11], y_round_in_s1[11], y_round_in_s0[11]}), .c ({new_AGEMA_signal_991, new_AGEMA_signal_990, y_rotated23[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_20_U1 ( .s (round[0]), .b ({y_round_in_s2[20], y_round_in_s1[20], y_round_in_s0[20]}), .a ({y_round_in_s2[12], y_round_in_s1[12], y_round_in_s0[12]}), .c ({new_AGEMA_signal_993, new_AGEMA_signal_992, y_rotated23[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_21_U1 ( .s (round[0]), .b ({y_round_in_s2[21], y_round_in_s1[21], y_round_in_s0[21]}), .a ({y_round_in_s2[13], y_round_in_s1[13], y_round_in_s0[13]}), .c ({new_AGEMA_signal_995, new_AGEMA_signal_994, y_rotated23[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_22_U1 ( .s (round[0]), .b ({y_round_in_s2[22], y_round_in_s1[22], y_round_in_s0[22]}), .a ({y_round_in_s2[14], y_round_in_s1[14], y_round_in_s0[14]}), .c ({new_AGEMA_signal_997, new_AGEMA_signal_996, y_rotated23[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_23_U1 ( .s (round[0]), .b ({y_round_in_s2[23], y_round_in_s1[23], y_round_in_s0[23]}), .a ({y_round_in_s2[15], y_round_in_s1[15], y_round_in_s0[15]}), .c ({new_AGEMA_signal_999, new_AGEMA_signal_998, y_rotated23[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_24_U1 ( .s (round[0]), .b ({y_round_in_s2[24], y_round_in_s1[24], y_round_in_s0[24]}), .a ({y_round_in_s2[16], y_round_in_s1[16], y_round_in_s0[16]}), .c ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, y_rotated23[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_25_U1 ( .s (round[0]), .b ({y_round_in_s2[25], y_round_in_s1[25], y_round_in_s0[25]}), .a ({y_round_in_s2[17], y_round_in_s1[17], y_round_in_s0[17]}), .c ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, y_rotated23[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_26_U1 ( .s (round[0]), .b ({y_round_in_s2[26], y_round_in_s1[26], y_round_in_s0[26]}), .a ({y_round_in_s2[18], y_round_in_s1[18], y_round_in_s0[18]}), .c ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, y_rotated23[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_27_U1 ( .s (round[0]), .b ({y_round_in_s2[27], y_round_in_s1[27], y_round_in_s0[27]}), .a ({y_round_in_s2[19], y_round_in_s1[19], y_round_in_s0[19]}), .c ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, y_rotated23[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_28_U1 ( .s (round[0]), .b ({y_round_in_s2[28], y_round_in_s1[28], y_round_in_s0[28]}), .a ({y_round_in_s2[20], y_round_in_s1[20], y_round_in_s0[20]}), .c ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, y_rotated23[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_29_U1 ( .s (round[0]), .b ({y_round_in_s2[29], y_round_in_s1[29], y_round_in_s0[29]}), .a ({y_round_in_s2[21], y_round_in_s1[21], y_round_in_s0[21]}), .c ({new_AGEMA_signal_1011, new_AGEMA_signal_1010, y_rotated23[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_30_U1 ( .s (round[0]), .b ({y_round_in_s2[30], y_round_in_s1[30], y_round_in_s0[30]}), .a ({y_round_in_s2[22], y_round_in_s1[22], y_round_in_s0[22]}), .c ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, y_rotated23[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M1_mux_inst_31_U1 ( .s (round[0]), .b ({y_round_in_s2[31], y_round_in_s1[31], y_round_in_s0[31]}), .a ({y_round_in_s2[23], y_round_in_s1[23], y_round_in_s0[23]}), .c ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, y_rotated23[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_0_U1 ( .s (round[1]), .b ({new_AGEMA_signal_829, new_AGEMA_signal_828, y_rotated01[0]}), .a ({new_AGEMA_signal_953, new_AGEMA_signal_952, y_rotated23[0]}), .c ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, y_rotated[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_1_U1 ( .s (round[1]), .b ({new_AGEMA_signal_835, new_AGEMA_signal_834, y_rotated01[1]}), .a ({new_AGEMA_signal_955, new_AGEMA_signal_954, y_rotated23[1]}), .c ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, y_rotated[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_2_U1 ( .s (round[1]), .b ({new_AGEMA_signal_841, new_AGEMA_signal_840, y_rotated01[2]}), .a ({new_AGEMA_signal_957, new_AGEMA_signal_956, y_rotated23[2]}), .c ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, y_rotated[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_3_U1 ( .s (round[1]), .b ({new_AGEMA_signal_847, new_AGEMA_signal_846, y_rotated01[3]}), .a ({new_AGEMA_signal_959, new_AGEMA_signal_958, y_rotated23[3]}), .c ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, y_rotated[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_4_U1 ( .s (round[1]), .b ({new_AGEMA_signal_853, new_AGEMA_signal_852, y_rotated01[4]}), .a ({new_AGEMA_signal_961, new_AGEMA_signal_960, y_rotated23[4]}), .c ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, y_rotated[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_5_U1 ( .s (round[1]), .b ({new_AGEMA_signal_859, new_AGEMA_signal_858, y_rotated01[5]}), .a ({new_AGEMA_signal_963, new_AGEMA_signal_962, y_rotated23[5]}), .c ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, y_rotated[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_6_U1 ( .s (round[1]), .b ({new_AGEMA_signal_865, new_AGEMA_signal_864, y_rotated01[6]}), .a ({new_AGEMA_signal_965, new_AGEMA_signal_964, y_rotated23[6]}), .c ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, y_rotated[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_7_U1 ( .s (round[1]), .b ({new_AGEMA_signal_871, new_AGEMA_signal_870, y_rotated01[7]}), .a ({new_AGEMA_signal_967, new_AGEMA_signal_966, y_rotated23[7]}), .c ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, y_rotated[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_8_U1 ( .s (round[1]), .b ({new_AGEMA_signal_877, new_AGEMA_signal_876, y_rotated01[8]}), .a ({new_AGEMA_signal_969, new_AGEMA_signal_968, y_rotated23[8]}), .c ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, y_rotated[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_9_U1 ( .s (round[1]), .b ({new_AGEMA_signal_883, new_AGEMA_signal_882, y_rotated01[9]}), .a ({new_AGEMA_signal_971, new_AGEMA_signal_970, y_rotated23[9]}), .c ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, y_rotated[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_10_U1 ( .s (round[1]), .b ({new_AGEMA_signal_889, new_AGEMA_signal_888, y_rotated01[10]}), .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, y_rotated23[10]}), .c ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, y_rotated[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_11_U1 ( .s (round[1]), .b ({new_AGEMA_signal_895, new_AGEMA_signal_894, y_rotated01[11]}), .a ({new_AGEMA_signal_975, new_AGEMA_signal_974, y_rotated23[11]}), .c ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, y_rotated[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_12_U1 ( .s (round[1]), .b ({new_AGEMA_signal_901, new_AGEMA_signal_900, y_rotated01[12]}), .a ({new_AGEMA_signal_977, new_AGEMA_signal_976, y_rotated23[12]}), .c ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, y_rotated[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_13_U1 ( .s (round[1]), .b ({new_AGEMA_signal_907, new_AGEMA_signal_906, y_rotated01[13]}), .a ({new_AGEMA_signal_979, new_AGEMA_signal_978, y_rotated23[13]}), .c ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, y_rotated[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_14_U1 ( .s (round[1]), .b ({new_AGEMA_signal_911, new_AGEMA_signal_910, y_rotated01[14]}), .a ({new_AGEMA_signal_981, new_AGEMA_signal_980, y_rotated23[14]}), .c ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, y_rotated[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_15_U1 ( .s (round[1]), .b ({new_AGEMA_signal_915, new_AGEMA_signal_914, y_rotated01[15]}), .a ({new_AGEMA_signal_983, new_AGEMA_signal_982, y_rotated23[15]}), .c ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, y_rotated[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_16_U1 ( .s (round[1]), .b ({new_AGEMA_signal_919, new_AGEMA_signal_918, y_rotated01[16]}), .a ({new_AGEMA_signal_985, new_AGEMA_signal_984, y_rotated23[16]}), .c ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, y_rotated[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_17_U1 ( .s (round[1]), .b ({new_AGEMA_signal_923, new_AGEMA_signal_922, y_rotated01[17]}), .a ({new_AGEMA_signal_987, new_AGEMA_signal_986, y_rotated23[17]}), .c ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, y_rotated[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_18_U1 ( .s (round[1]), .b ({new_AGEMA_signal_925, new_AGEMA_signal_924, y_rotated01[18]}), .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, y_rotated23[18]}), .c ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, y_rotated[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_19_U1 ( .s (round[1]), .b ({new_AGEMA_signal_927, new_AGEMA_signal_926, y_rotated01[19]}), .a ({new_AGEMA_signal_991, new_AGEMA_signal_990, y_rotated23[19]}), .c ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, y_rotated[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_20_U1 ( .s (round[1]), .b ({new_AGEMA_signal_929, new_AGEMA_signal_928, y_rotated01[20]}), .a ({new_AGEMA_signal_993, new_AGEMA_signal_992, y_rotated23[20]}), .c ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, y_rotated[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_21_U1 ( .s (round[1]), .b ({new_AGEMA_signal_931, new_AGEMA_signal_930, y_rotated01[21]}), .a ({new_AGEMA_signal_995, new_AGEMA_signal_994, y_rotated23[21]}), .c ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, y_rotated[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_22_U1 ( .s (round[1]), .b ({new_AGEMA_signal_933, new_AGEMA_signal_932, y_rotated01[22]}), .a ({new_AGEMA_signal_997, new_AGEMA_signal_996, y_rotated23[22]}), .c ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, y_rotated[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_23_U1 ( .s (round[1]), .b ({new_AGEMA_signal_935, new_AGEMA_signal_934, y_rotated01[23]}), .a ({new_AGEMA_signal_999, new_AGEMA_signal_998, y_rotated23[23]}), .c ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, y_rotated[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_24_U1 ( .s (round[1]), .b ({new_AGEMA_signal_937, new_AGEMA_signal_936, y_rotated01[24]}), .a ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, y_rotated23[24]}), .c ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, y_rotated[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_25_U1 ( .s (round[1]), .b ({new_AGEMA_signal_939, new_AGEMA_signal_938, y_rotated01[25]}), .a ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, y_rotated23[25]}), .c ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, y_rotated[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_26_U1 ( .s (round[1]), .b ({new_AGEMA_signal_941, new_AGEMA_signal_940, y_rotated01[26]}), .a ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, y_rotated23[26]}), .c ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, y_rotated[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_27_U1 ( .s (round[1]), .b ({new_AGEMA_signal_943, new_AGEMA_signal_942, y_rotated01[27]}), .a ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, y_rotated23[27]}), .c ({new_AGEMA_signal_1071, new_AGEMA_signal_1070, y_rotated[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_28_U1 ( .s (round[1]), .b ({new_AGEMA_signal_945, new_AGEMA_signal_944, y_rotated01[28]}), .a ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, y_rotated23[28]}), .c ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, y_rotated[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_29_U1 ( .s (round[1]), .b ({new_AGEMA_signal_947, new_AGEMA_signal_946, y_rotated01[29]}), .a ({new_AGEMA_signal_1011, new_AGEMA_signal_1010, y_rotated23[29]}), .c ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, y_rotated[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_30_U1 ( .s (round[1]), .b ({new_AGEMA_signal_949, new_AGEMA_signal_948, y_rotated01[30]}), .a ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, y_rotated23[30]}), .c ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, y_rotated[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M3_mux_inst_31_U1 ( .s (round[1]), .b ({new_AGEMA_signal_951, new_AGEMA_signal_950, y_rotated01[31]}), .a ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, y_rotated23[31]}), .c ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, y_rotated[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_0_U1 ( .a ({x_round_in_s2[0], x_round_in_s1[0], x_round_in_s0[0]}), .b ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, y_rotated[0]}), .c ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, sum[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_1_U1 ( .a ({x_round_in_s2[1], x_round_in_s1[1], x_round_in_s0[1]}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, y_rotated[1]}), .c ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, AdderIns_p6[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_2_U1 ( .a ({x_round_in_s2[2], x_round_in_s1[2], x_round_in_s0[2]}), .b ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, y_rotated[2]}), .c ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, AdderIns_p6[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_3_U1 ( .a ({x_round_in_s2[3], x_round_in_s1[3], x_round_in_s0[3]}), .b ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, y_rotated[3]}), .c ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, AdderIns_p6[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_4_U1 ( .a ({x_round_in_s2[4], x_round_in_s1[4], x_round_in_s0[4]}), .b ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, y_rotated[4]}), .c ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, AdderIns_p6[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_5_U1 ( .a ({x_round_in_s2[5], x_round_in_s1[5], x_round_in_s0[5]}), .b ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, y_rotated[5]}), .c ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, AdderIns_p6[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_6_U1 ( .a ({x_round_in_s2[6], x_round_in_s1[6], x_round_in_s0[6]}), .b ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, y_rotated[6]}), .c ({new_AGEMA_signal_1119, new_AGEMA_signal_1118, AdderIns_p6[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_7_U1 ( .a ({x_round_in_s2[7], x_round_in_s1[7], x_round_in_s0[7]}), .b ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, y_rotated[7]}), .c ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, AdderIns_p6[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_8_U1 ( .a ({x_round_in_s2[8], x_round_in_s1[8], x_round_in_s0[8]}), .b ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, y_rotated[8]}), .c ({new_AGEMA_signal_1131, new_AGEMA_signal_1130, AdderIns_p6[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_9_U1 ( .a ({x_round_in_s2[9], x_round_in_s1[9], x_round_in_s0[9]}), .b ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, y_rotated[9]}), .c ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, AdderIns_p6[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_10_U1 ( .a ({x_round_in_s2[10], x_round_in_s1[10], x_round_in_s0[10]}), .b ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, y_rotated[10]}), .c ({new_AGEMA_signal_1143, new_AGEMA_signal_1142, AdderIns_p6[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_11_U1 ( .a ({x_round_in_s2[11], x_round_in_s1[11], x_round_in_s0[11]}), .b ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, y_rotated[11]}), .c ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, AdderIns_p6[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_12_U1 ( .a ({x_round_in_s2[12], x_round_in_s1[12], x_round_in_s0[12]}), .b ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, y_rotated[12]}), .c ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, AdderIns_p6[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_13_U1 ( .a ({x_round_in_s2[13], x_round_in_s1[13], x_round_in_s0[13]}), .b ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, y_rotated[13]}), .c ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, AdderIns_p6[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_14_U1 ( .a ({x_round_in_s2[14], x_round_in_s1[14], x_round_in_s0[14]}), .b ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, y_rotated[14]}), .c ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, AdderIns_p6[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_15_U1 ( .a ({x_round_in_s2[15], x_round_in_s1[15], x_round_in_s0[15]}), .b ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, y_rotated[15]}), .c ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, AdderIns_p6[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_16_U1 ( .a ({x_round_in_s2[16], x_round_in_s1[16], x_round_in_s0[16]}), .b ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, y_rotated[16]}), .c ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, AdderIns_p6[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_17_U1 ( .a ({x_round_in_s2[17], x_round_in_s1[17], x_round_in_s0[17]}), .b ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, y_rotated[17]}), .c ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, AdderIns_p6[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_18_U1 ( .a ({x_round_in_s2[18], x_round_in_s1[18], x_round_in_s0[18]}), .b ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, y_rotated[18]}), .c ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, AdderIns_p6[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_19_U1 ( .a ({x_round_in_s2[19], x_round_in_s1[19], x_round_in_s0[19]}), .b ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, y_rotated[19]}), .c ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, AdderIns_p6[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_20_U1 ( .a ({x_round_in_s2[20], x_round_in_s1[20], x_round_in_s0[20]}), .b ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, y_rotated[20]}), .c ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, AdderIns_p6[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_21_U1 ( .a ({x_round_in_s2[21], x_round_in_s1[21], x_round_in_s0[21]}), .b ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, y_rotated[21]}), .c ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, AdderIns_p6[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_22_U1 ( .a ({x_round_in_s2[22], x_round_in_s1[22], x_round_in_s0[22]}), .b ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, y_rotated[22]}), .c ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, AdderIns_p6[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_23_U1 ( .a ({x_round_in_s2[23], x_round_in_s1[23], x_round_in_s0[23]}), .b ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, y_rotated[23]}), .c ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, AdderIns_p6[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_24_U1 ( .a ({x_round_in_s2[24], x_round_in_s1[24], x_round_in_s0[24]}), .b ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, y_rotated[24]}), .c ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, AdderIns_p6[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_25_U1 ( .a ({x_round_in_s2[25], x_round_in_s1[25], x_round_in_s0[25]}), .b ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, y_rotated[25]}), .c ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, AdderIns_p6[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_26_U1 ( .a ({x_round_in_s2[26], x_round_in_s1[26], x_round_in_s0[26]}), .b ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, y_rotated[26]}), .c ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, AdderIns_p6[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_27_U1 ( .a ({x_round_in_s2[27], x_round_in_s1[27], x_round_in_s0[27]}), .b ({new_AGEMA_signal_1071, new_AGEMA_signal_1070, y_rotated[27]}), .c ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, AdderIns_p6[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_28_U1 ( .a ({x_round_in_s2[28], x_round_in_s1[28], x_round_in_s0[28]}), .b ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, y_rotated[28]}), .c ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, AdderIns_p6[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_29_U1 ( .a ({x_round_in_s2[29], x_round_in_s1[29], x_round_in_s0[29]}), .b ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, y_rotated[29]}), .c ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, AdderIns_p6[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_30_U1 ( .a ({x_round_in_s2[30], x_round_in_s1[30], x_round_in_s0[30]}), .b ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, y_rotated[30]}), .c ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, AdderIns_p6[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_31_U1 ( .a ({x_round_in_s2[31], x_round_in_s1[31], x_round_in_s0[31]}), .b ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, y_rotated[31]}), .c ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, AdderIns_p6[31]}) ) ;
    //ClockGatingController #(10) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) U140 ( .a ({1'b0, 1'b0, round_constant[1]}), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, sum[1]}), .c ({x_round_out_s2[1], x_round_out_s1[1], x_round_out_s0[1]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_0_a1_U1 ( .a ({x_round_in_s2[0], x_round_in_s1[0], x_round_in_s0[0]}), .b ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, y_rotated[0]}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, AdderIns_g1[0]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_1_a1_U1 ( .a ({x_round_in_s2[1], x_round_in_s1[1], x_round_in_s0[1]}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, y_rotated[1]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, AdderIns_g1[1]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_2_a1_U1 ( .a ({x_round_in_s2[2], x_round_in_s1[2], x_round_in_s0[2]}), .b ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, y_rotated[2]}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, AdderIns_g1[2]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_3_a1_U1 ( .a ({x_round_in_s2[3], x_round_in_s1[3], x_round_in_s0[3]}), .b ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, y_rotated[3]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, AdderIns_g1[3]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_4_a1_U1 ( .a ({x_round_in_s2[4], x_round_in_s1[4], x_round_in_s0[4]}), .b ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, y_rotated[4]}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, AdderIns_g1[4]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_5_a1_U1 ( .a ({x_round_in_s2[5], x_round_in_s1[5], x_round_in_s0[5]}), .b ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, y_rotated[5]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, AdderIns_g1[5]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_6_a1_U1 ( .a ({x_round_in_s2[6], x_round_in_s1[6], x_round_in_s0[6]}), .b ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, y_rotated[6]}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, AdderIns_g1[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_7_a1_U1 ( .a ({x_round_in_s2[7], x_round_in_s1[7], x_round_in_s0[7]}), .b ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, y_rotated[7]}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, AdderIns_g1[7]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_8_a1_U1 ( .a ({x_round_in_s2[8], x_round_in_s1[8], x_round_in_s0[8]}), .b ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, y_rotated[8]}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, AdderIns_g1[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_9_a1_U1 ( .a ({x_round_in_s2[9], x_round_in_s1[9], x_round_in_s0[9]}), .b ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, y_rotated[9]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, AdderIns_g1[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_10_a1_U1 ( .a ({x_round_in_s2[10], x_round_in_s1[10], x_round_in_s0[10]}), .b ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, y_rotated[10]}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, AdderIns_g1[10]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_11_a1_U1 ( .a ({x_round_in_s2[11], x_round_in_s1[11], x_round_in_s0[11]}), .b ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, y_rotated[11]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, AdderIns_g1[11]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_12_a1_U1 ( .a ({x_round_in_s2[12], x_round_in_s1[12], x_round_in_s0[12]}), .b ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, y_rotated[12]}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, AdderIns_g1[12]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_13_a1_U1 ( .a ({x_round_in_s2[13], x_round_in_s1[13], x_round_in_s0[13]}), .b ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, y_rotated[13]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, AdderIns_g1[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_14_a1_U1 ( .a ({x_round_in_s2[14], x_round_in_s1[14], x_round_in_s0[14]}), .b ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, y_rotated[14]}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, AdderIns_g1[14]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_15_a1_U1 ( .a ({x_round_in_s2[15], x_round_in_s1[15], x_round_in_s0[15]}), .b ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, y_rotated[15]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, AdderIns_g1[15]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_16_a1_U1 ( .a ({x_round_in_s2[16], x_round_in_s1[16], x_round_in_s0[16]}), .b ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, y_rotated[16]}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, AdderIns_g1[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_17_a1_U1 ( .a ({x_round_in_s2[17], x_round_in_s1[17], x_round_in_s0[17]}), .b ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, y_rotated[17]}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, AdderIns_g1[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_18_a1_U1 ( .a ({x_round_in_s2[18], x_round_in_s1[18], x_round_in_s0[18]}), .b ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, y_rotated[18]}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, AdderIns_g1[18]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_19_a1_U1 ( .a ({x_round_in_s2[19], x_round_in_s1[19], x_round_in_s0[19]}), .b ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, y_rotated[19]}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, AdderIns_g1[19]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_20_a1_U1 ( .a ({x_round_in_s2[20], x_round_in_s1[20], x_round_in_s0[20]}), .b ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, y_rotated[20]}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, AdderIns_g1[20]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_21_a1_U1 ( .a ({x_round_in_s2[21], x_round_in_s1[21], x_round_in_s0[21]}), .b ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, y_rotated[21]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, AdderIns_g1[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_22_a1_U1 ( .a ({x_round_in_s2[22], x_round_in_s1[22], x_round_in_s0[22]}), .b ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, y_rotated[22]}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, AdderIns_g1[22]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_23_a1_U1 ( .a ({x_round_in_s2[23], x_round_in_s1[23], x_round_in_s0[23]}), .b ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, y_rotated[23]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, AdderIns_g1[23]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_24_a1_U1 ( .a ({x_round_in_s2[24], x_round_in_s1[24], x_round_in_s0[24]}), .b ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, y_rotated[24]}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, AdderIns_g1[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_25_a1_U1 ( .a ({x_round_in_s2[25], x_round_in_s1[25], x_round_in_s0[25]}), .b ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, y_rotated[25]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, AdderIns_g1[25]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_26_a1_U1 ( .a ({x_round_in_s2[26], x_round_in_s1[26], x_round_in_s0[26]}), .b ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, y_rotated[26]}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, AdderIns_g1[26]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_27_a1_U1 ( .a ({x_round_in_s2[27], x_round_in_s1[27], x_round_in_s0[27]}), .b ({new_AGEMA_signal_1071, new_AGEMA_signal_1070, y_rotated[27]}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, AdderIns_g1[27]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_28_a1_U1 ( .a ({x_round_in_s2[28], x_round_in_s1[28], x_round_in_s0[28]}), .b ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, y_rotated[28]}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, AdderIns_g1[28]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_29_a1_U1 ( .a ({x_round_in_s2[29], x_round_in_s1[29], x_round_in_s0[29]}), .b ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, y_rotated[29]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, AdderIns_g1[29]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s1_pg_30_a1_U1 ( .a ({x_round_in_s2[30], x_round_in_s1[30], x_round_in_s0[30]}), .b ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, y_rotated[30]}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, AdderIns_g1[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_gc_0_a1_U1 ( .a ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, AdderIns_g1[0]}), .b ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, AdderIns_s2_gc_0_a1_t}), .c ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, AdderIns_g6[0]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, sum[0]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, AdderIns_s2_gc_0_a1_t}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_0_a2_U1 ( .a ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, sum[0]}), .b ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, AdderIns_p6[1]}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, AdderIns_p2[0]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, AdderIns_p6[1]}), .b ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, AdderIns_p6[2]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, AdderIns_p2[1]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, AdderIns_p6[2]}), .b ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, AdderIns_p6[3]}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, AdderIns_p2[2]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, AdderIns_p6[3]}), .b ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, AdderIns_p6[4]}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, AdderIns_p2[3]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, AdderIns_p6[4]}), .b ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, AdderIns_p6[5]}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, AdderIns_p2[4]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, AdderIns_p6[5]}), .b ({new_AGEMA_signal_1119, new_AGEMA_signal_1118, AdderIns_p6[6]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, AdderIns_p2[5]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1119, new_AGEMA_signal_1118, AdderIns_p6[6]}), .b ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, AdderIns_p6[7]}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, AdderIns_p2[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, AdderIns_p6[7]}), .b ({new_AGEMA_signal_1131, new_AGEMA_signal_1130, AdderIns_p6[8]}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, AdderIns_p2[7]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1131, new_AGEMA_signal_1130, AdderIns_p6[8]}), .b ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, AdderIns_p6[9]}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, AdderIns_p2[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, AdderIns_p6[9]}), .b ({new_AGEMA_signal_1143, new_AGEMA_signal_1142, AdderIns_p6[10]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, AdderIns_p2[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1143, new_AGEMA_signal_1142, AdderIns_p6[10]}), .b ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, AdderIns_p6[11]}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, AdderIns_p2[10]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, AdderIns_p6[11]}), .b ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, AdderIns_p6[12]}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, AdderIns_p2[11]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, AdderIns_p6[12]}), .b ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, AdderIns_p6[13]}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, AdderIns_p2[12]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, AdderIns_p6[13]}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, AdderIns_p6[14]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, AdderIns_p2[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, AdderIns_p6[14]}), .b ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, AdderIns_p6[15]}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, AdderIns_p2[14]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_15_a2_U1 ( .a ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, AdderIns_p6[15]}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, AdderIns_p6[16]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, AdderIns_p2[15]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_16_a2_U1 ( .a ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, AdderIns_p6[16]}), .b ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, AdderIns_p6[17]}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, AdderIns_p2[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_17_a2_U1 ( .a ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, AdderIns_p6[17]}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, AdderIns_p6[18]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, AdderIns_p2[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_18_a2_U1 ( .a ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, AdderIns_p6[18]}), .b ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, AdderIns_p6[19]}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, AdderIns_p2[18]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_19_a2_U1 ( .a ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, AdderIns_p6[19]}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, AdderIns_p6[20]}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, AdderIns_p2[19]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_20_a2_U1 ( .a ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, AdderIns_p6[20]}), .b ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, AdderIns_p6[21]}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, AdderIns_p2[20]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_21_a2_U1 ( .a ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, AdderIns_p6[21]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, AdderIns_p6[22]}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, AdderIns_p2[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_22_a2_U1 ( .a ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, AdderIns_p6[22]}), .b ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, AdderIns_p6[23]}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, AdderIns_p2[22]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_23_a2_U1 ( .a ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, AdderIns_p6[23]}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, AdderIns_p6[24]}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, AdderIns_p2[23]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_24_a2_U1 ( .a ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, AdderIns_p6[24]}), .b ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, AdderIns_p6[25]}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, AdderIns_p2[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_25_a2_U1 ( .a ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, AdderIns_p6[25]}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, AdderIns_p6[26]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, AdderIns_p2[25]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_26_a2_U1 ( .a ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, AdderIns_p6[26]}), .b ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, AdderIns_p6[27]}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, AdderIns_p2[26]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_27_a2_U1 ( .a ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, AdderIns_p6[27]}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, AdderIns_p6[28]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, AdderIns_p2[27]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_28_a2_U1 ( .a ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, AdderIns_p6[28]}), .b ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, AdderIns_p6[29]}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, AdderIns_p2[28]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_29_a2_U1 ( .a ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, AdderIns_p6[29]}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, AdderIns_p6[30]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, AdderIns_p2[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U11 ( .a ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, AdderIns_p6[1]}), .c ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, sum[1]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) U151 ( .a ({1'b0, 1'b0, round_constant[2]}), .b ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, sum[2]}), .c ({x_round_out_s2[2], x_round_out_s1[2], x_round_out_s0[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U154 ( .a ({1'b0, 1'b0, round_constant[3]}), .b ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, sum[3]}), .c ({x_round_out_s2[3], x_round_out_s1[3], x_round_out_s0[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_0_a1_U1 ( .a ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, AdderIns_g1[1]}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, AdderIns_s2_bc_0_a1_t}), .c ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, AdderIns_g2[1]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, AdderIns_g1[0]}), .b ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, AdderIns_p6[1]}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, AdderIns_s2_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_1_a1_U1 ( .a ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, AdderIns_g1[2]}), .b ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, AdderIns_s2_bc_1_a1_t}), .c ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, AdderIns_g2[2]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, AdderIns_g1[1]}), .b ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, AdderIns_p6[2]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, AdderIns_s2_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_2_a1_U1 ( .a ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, AdderIns_g1[3]}), .b ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, AdderIns_s2_bc_2_a1_t}), .c ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, AdderIns_g2[3]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, AdderIns_g1[2]}), .b ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, AdderIns_p6[3]}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, AdderIns_s2_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_3_a1_U1 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, AdderIns_g1[4]}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, AdderIns_s2_bc_3_a1_t}), .c ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, AdderIns_g2[4]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, AdderIns_g1[3]}), .b ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, AdderIns_p6[4]}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, AdderIns_s2_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_4_a1_U1 ( .a ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, AdderIns_g1[5]}), .b ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, AdderIns_s2_bc_4_a1_t}), .c ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, AdderIns_g2[5]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, AdderIns_g1[4]}), .b ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, AdderIns_p6[5]}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, AdderIns_s2_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_5_a1_U1 ( .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, AdderIns_g1[6]}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, AdderIns_s2_bc_5_a1_t}), .c ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, AdderIns_g2[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, AdderIns_g1[5]}), .b ({new_AGEMA_signal_1119, new_AGEMA_signal_1118, AdderIns_p6[6]}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, AdderIns_s2_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_6_a1_U1 ( .a ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, AdderIns_g1[7]}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, AdderIns_s2_bc_6_a1_t}), .c ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, AdderIns_g2[7]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, AdderIns_g1[6]}), .b ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, AdderIns_p6[7]}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, AdderIns_s2_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_7_a1_U1 ( .a ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, AdderIns_g1[8]}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, AdderIns_s2_bc_7_a1_t}), .c ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, AdderIns_g2[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, AdderIns_g1[7]}), .b ({new_AGEMA_signal_1131, new_AGEMA_signal_1130, AdderIns_p6[8]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, AdderIns_s2_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_8_a1_U1 ( .a ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, AdderIns_g1[9]}), .b ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, AdderIns_s2_bc_8_a1_t}), .c ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, AdderIns_g2[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, AdderIns_g1[8]}), .b ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, AdderIns_p6[9]}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, AdderIns_s2_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_9_a1_U1 ( .a ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, AdderIns_g1[10]}), .b ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, AdderIns_s2_bc_9_a1_t}), .c ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, AdderIns_g2[10]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, AdderIns_g1[9]}), .b ({new_AGEMA_signal_1143, new_AGEMA_signal_1142, AdderIns_p6[10]}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, AdderIns_s2_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_10_a1_U1 ( .a ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, AdderIns_g1[11]}), .b ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, AdderIns_s2_bc_10_a1_t}), .c ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, AdderIns_g2[11]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, AdderIns_g1[10]}), .b ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, AdderIns_p6[11]}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, AdderIns_s2_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_11_a1_U1 ( .a ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, AdderIns_g1[12]}), .b ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, AdderIns_s2_bc_11_a1_t}), .c ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, AdderIns_g2[12]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, AdderIns_g1[11]}), .b ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, AdderIns_p6[12]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, AdderIns_s2_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_12_a1_U1 ( .a ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, AdderIns_g1[13]}), .b ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, AdderIns_s2_bc_12_a1_t}), .c ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, AdderIns_g2[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, AdderIns_g1[12]}), .b ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, AdderIns_p6[13]}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, AdderIns_s2_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_13_a1_U1 ( .a ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, AdderIns_g1[14]}), .b ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, AdderIns_s2_bc_13_a1_t}), .c ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, AdderIns_g2[14]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, AdderIns_g1[13]}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, AdderIns_p6[14]}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, AdderIns_s2_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_14_a1_U1 ( .a ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, AdderIns_g1[15]}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, AdderIns_s2_bc_14_a1_t}), .c ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, AdderIns_g2[15]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, AdderIns_g1[14]}), .b ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, AdderIns_p6[15]}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, AdderIns_s2_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_15_a1_U1 ( .a ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, AdderIns_g1[16]}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, AdderIns_s2_bc_15_a1_t}), .c ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, AdderIns_g2[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, AdderIns_g1[15]}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, AdderIns_p6[16]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, AdderIns_s2_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_16_a1_U1 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, AdderIns_g1[17]}), .b ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, AdderIns_s2_bc_16_a1_t}), .c ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, AdderIns_g2[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_16_a1_a1_U1 ( .a ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, AdderIns_g1[16]}), .b ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, AdderIns_p6[17]}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, AdderIns_s2_bc_16_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_17_a1_U1 ( .a ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, AdderIns_g1[18]}), .b ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, AdderIns_s2_bc_17_a1_t}), .c ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, AdderIns_g2[18]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_17_a1_a1_U1 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, AdderIns_g1[17]}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, AdderIns_p6[18]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, AdderIns_s2_bc_17_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_18_a1_U1 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, AdderIns_g1[19]}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, AdderIns_s2_bc_18_a1_t}), .c ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, AdderIns_g2[19]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_18_a1_a1_U1 ( .a ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, AdderIns_g1[18]}), .b ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, AdderIns_p6[19]}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, AdderIns_s2_bc_18_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_19_a1_U1 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, AdderIns_g1[20]}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, AdderIns_s2_bc_19_a1_t}), .c ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, AdderIns_g2[20]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_19_a1_a1_U1 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, AdderIns_g1[19]}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, AdderIns_p6[20]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, AdderIns_s2_bc_19_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_20_a1_U1 ( .a ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, AdderIns_g1[21]}), .b ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, AdderIns_s2_bc_20_a1_t}), .c ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, AdderIns_g2[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_20_a1_a1_U1 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, AdderIns_g1[20]}), .b ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, AdderIns_p6[21]}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, AdderIns_s2_bc_20_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_21_a1_U1 ( .a ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, AdderIns_g1[22]}), .b ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, AdderIns_s2_bc_21_a1_t}), .c ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, AdderIns_g2[22]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_21_a1_a1_U1 ( .a ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, AdderIns_g1[21]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, AdderIns_p6[22]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, AdderIns_s2_bc_21_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_22_a1_U1 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, AdderIns_g1[23]}), .b ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, AdderIns_s2_bc_22_a1_t}), .c ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, AdderIns_g2[23]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_22_a1_a1_U1 ( .a ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, AdderIns_g1[22]}), .b ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, AdderIns_p6[23]}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, AdderIns_s2_bc_22_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_23_a1_U1 ( .a ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, AdderIns_g1[24]}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, AdderIns_s2_bc_23_a1_t}), .c ({new_AGEMA_signal_1443, new_AGEMA_signal_1442, AdderIns_g2[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_23_a1_a1_U1 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, AdderIns_g1[23]}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, AdderIns_p6[24]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, AdderIns_s2_bc_23_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_24_a1_U1 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, AdderIns_g1[25]}), .b ({new_AGEMA_signal_1371, new_AGEMA_signal_1370, AdderIns_s2_bc_24_a1_t}), .c ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, AdderIns_g2[25]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_24_a1_a1_U1 ( .a ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, AdderIns_g1[24]}), .b ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, AdderIns_p6[25]}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1371, new_AGEMA_signal_1370, AdderIns_s2_bc_24_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_25_a1_U1 ( .a ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, AdderIns_g1[26]}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, AdderIns_s2_bc_25_a1_t}), .c ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, AdderIns_g2[26]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_25_a1_a1_U1 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, AdderIns_g1[25]}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, AdderIns_p6[26]}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, AdderIns_s2_bc_25_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_26_a1_U1 ( .a ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, AdderIns_g1[27]}), .b ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, AdderIns_s2_bc_26_a1_t}), .c ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, AdderIns_g2[27]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_26_a1_a1_U1 ( .a ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, AdderIns_g1[26]}), .b ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, AdderIns_p6[27]}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, AdderIns_s2_bc_26_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_27_a1_U1 ( .a ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, AdderIns_g1[28]}), .b ({new_AGEMA_signal_1383, new_AGEMA_signal_1382, AdderIns_s2_bc_27_a1_t}), .c ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, AdderIns_g2[28]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_27_a1_a1_U1 ( .a ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, AdderIns_g1[27]}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, AdderIns_p6[28]}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_1383, new_AGEMA_signal_1382, AdderIns_s2_bc_27_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_28_a1_U1 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, AdderIns_g1[29]}), .b ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, AdderIns_s2_bc_28_a1_t}), .c ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, AdderIns_g2[29]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_28_a1_a1_U1 ( .a ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, AdderIns_g1[28]}), .b ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, AdderIns_p6[29]}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, AdderIns_s2_bc_28_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_29_a1_U1 ( .a ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, AdderIns_g1[30]}), .b ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, AdderIns_s2_bc_29_a1_t}), .c ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, AdderIns_g2[30]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s2_bc_29_a1_a1_U1 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, AdderIns_g1[29]}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, AdderIns_p6[30]}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, AdderIns_s2_bc_29_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_gc_0_a1_U1 ( .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, AdderIns_g2[1]}), .b ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, AdderIns_s3_gc_0_a1_t}), .c ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, AdderIns_g6[1]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, AdderIns_p2[0]}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, AdderIns_s3_gc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_gc_1_a1_U1 ( .a ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, AdderIns_g2[2]}), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, AdderIns_s3_gc_1_a1_t}), .c ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, AdderIns_g6[2]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, AdderIns_p2[1]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, AdderIns_s3_gc_1_a1_t}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_0_a2_U1 ( .a ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, AdderIns_p2[0]}), .b ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, AdderIns_p2[2]}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, AdderIns_p3[0]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, AdderIns_p2[1]}), .b ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, AdderIns_p2[3]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, AdderIns_p3[1]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, AdderIns_p2[2]}), .b ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, AdderIns_p2[4]}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, AdderIns_p3[2]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, AdderIns_p2[3]}), .b ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, AdderIns_p2[5]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, AdderIns_p3[3]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, AdderIns_p2[4]}), .b ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, AdderIns_p2[6]}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, AdderIns_p3[4]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, AdderIns_p2[5]}), .b ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, AdderIns_p2[7]}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, AdderIns_p3[5]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, AdderIns_p2[6]}), .b ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, AdderIns_p2[8]}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, AdderIns_p3[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, AdderIns_p2[7]}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, AdderIns_p2[9]}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, AdderIns_p3[7]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, AdderIns_p2[8]}), .b ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, AdderIns_p2[10]}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, AdderIns_p3[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, AdderIns_p2[9]}), .b ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, AdderIns_p2[11]}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, AdderIns_p3[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, AdderIns_p2[10]}), .b ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, AdderIns_p2[12]}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, AdderIns_p3[10]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, AdderIns_p2[11]}), .b ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, AdderIns_p2[13]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, AdderIns_p3[11]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, AdderIns_p2[12]}), .b ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, AdderIns_p2[14]}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, AdderIns_p3[12]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, AdderIns_p2[13]}), .b ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, AdderIns_p2[15]}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, AdderIns_p3[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, AdderIns_p2[14]}), .b ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, AdderIns_p2[16]}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, AdderIns_p3[14]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_15_a2_U1 ( .a ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, AdderIns_p2[15]}), .b ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, AdderIns_p2[17]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, AdderIns_p3[15]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_16_a2_U1 ( .a ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, AdderIns_p2[16]}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, AdderIns_p2[18]}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, AdderIns_p3[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_17_a2_U1 ( .a ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, AdderIns_p2[17]}), .b ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, AdderIns_p2[19]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, AdderIns_p3[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_18_a2_U1 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, AdderIns_p2[18]}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, AdderIns_p2[20]}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, AdderIns_p3[18]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_19_a2_U1 ( .a ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, AdderIns_p2[19]}), .b ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, AdderIns_p2[21]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, AdderIns_p3[19]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_20_a2_U1 ( .a ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, AdderIns_p2[20]}), .b ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, AdderIns_p2[22]}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, AdderIns_p3[20]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_21_a2_U1 ( .a ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, AdderIns_p2[21]}), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, AdderIns_p2[23]}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, AdderIns_p3[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_22_a2_U1 ( .a ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, AdderIns_p2[22]}), .b ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, AdderIns_p2[24]}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, AdderIns_p3[22]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_23_a2_U1 ( .a ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, AdderIns_p2[23]}), .b ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, AdderIns_p2[25]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, AdderIns_p3[23]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_24_a2_U1 ( .a ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, AdderIns_p2[24]}), .b ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, AdderIns_p2[26]}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, AdderIns_p3[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_25_a2_U1 ( .a ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, AdderIns_p2[25]}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, AdderIns_p2[27]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, AdderIns_p3[25]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_26_a2_U1 ( .a ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, AdderIns_p2[26]}), .b ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, AdderIns_p2[28]}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, AdderIns_p3[26]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_27_a2_U1 ( .a ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, AdderIns_p2[27]}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, AdderIns_p2[29]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, AdderIns_p3[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U25 ( .a ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, AdderIns_g6[2]}), .b ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, AdderIns_p6[3]}), .c ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, sum[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U22 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, AdderIns_g6[1]}), .b ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, AdderIns_p6[2]}), .c ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, sum[2]}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) U155 ( .a ({1'b0, 1'b0, round_constant[4]}), .b ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, sum[4]}), .c ({x_round_out_s2[4], x_round_out_s1[4], x_round_out_s0[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U156 ( .a ({1'b0, 1'b0, round_constant[5]}), .b ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, sum[5]}), .c ({x_round_out_s2[5], x_round_out_s1[5], x_round_out_s0[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U157 ( .a ({1'b0, 1'b0, round_constant[6]}), .b ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, sum[6]}), .c ({x_round_out_s2[6], x_round_out_s1[6], x_round_out_s0[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U158 ( .a ({1'b0, 1'b0, round_constant[7]}), .b ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, sum[7]}), .c ({x_round_out_s2[7], x_round_out_s1[7], x_round_out_s0[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_0_a1_U1 ( .a ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, AdderIns_g2[3]}), .b ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, AdderIns_s3_bc_0_a1_t}), .c ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, AdderIns_g3[3]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, AdderIns_g2[1]}), .b ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, AdderIns_p2[2]}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, AdderIns_s3_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_1_a1_U1 ( .a ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, AdderIns_g2[4]}), .b ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, AdderIns_s3_bc_1_a1_t}), .c ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, AdderIns_g3[4]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, AdderIns_g2[2]}), .b ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, AdderIns_p2[3]}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, AdderIns_s3_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_2_a1_U1 ( .a ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, AdderIns_g2[5]}), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, AdderIns_s3_bc_2_a1_t}), .c ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, AdderIns_g3[5]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, AdderIns_g2[3]}), .b ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, AdderIns_p2[4]}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, AdderIns_s3_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_3_a1_U1 ( .a ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, AdderIns_g2[6]}), .b ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, AdderIns_s3_bc_3_a1_t}), .c ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, AdderIns_g3[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, AdderIns_g2[4]}), .b ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, AdderIns_p2[5]}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, AdderIns_s3_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_4_a1_U1 ( .a ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, AdderIns_g2[7]}), .b ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, AdderIns_s3_bc_4_a1_t}), .c ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, AdderIns_g3[7]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, AdderIns_g2[5]}), .b ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, AdderIns_p2[6]}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, AdderIns_s3_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_5_a1_U1 ( .a ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, AdderIns_g2[8]}), .b ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, AdderIns_s3_bc_5_a1_t}), .c ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, AdderIns_g3[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, AdderIns_g2[6]}), .b ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, AdderIns_p2[7]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, AdderIns_s3_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_6_a1_U1 ( .a ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, AdderIns_g2[9]}), .b ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, AdderIns_s3_bc_6_a1_t}), .c ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, AdderIns_g3[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, AdderIns_g2[7]}), .b ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, AdderIns_p2[8]}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, AdderIns_s3_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_7_a1_U1 ( .a ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, AdderIns_g2[10]}), .b ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, AdderIns_s3_bc_7_a1_t}), .c ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, AdderIns_g3[10]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, AdderIns_g2[8]}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, AdderIns_p2[9]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, AdderIns_s3_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_8_a1_U1 ( .a ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, AdderIns_g2[11]}), .b ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, AdderIns_s3_bc_8_a1_t}), .c ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, AdderIns_g3[11]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, AdderIns_g2[9]}), .b ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, AdderIns_p2[10]}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, AdderIns_s3_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_9_a1_U1 ( .a ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, AdderIns_g2[12]}), .b ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, AdderIns_s3_bc_9_a1_t}), .c ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, AdderIns_g3[12]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, AdderIns_g2[10]}), .b ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, AdderIns_p2[11]}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, AdderIns_s3_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_10_a1_U1 ( .a ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, AdderIns_g2[13]}), .b ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, AdderIns_s3_bc_10_a1_t}), .c ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, AdderIns_g3[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, AdderIns_g2[11]}), .b ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, AdderIns_p2[12]}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, AdderIns_s3_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_11_a1_U1 ( .a ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, AdderIns_g2[14]}), .b ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, AdderIns_s3_bc_11_a1_t}), .c ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, AdderIns_g3[14]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, AdderIns_g2[12]}), .b ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, AdderIns_p2[13]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, AdderIns_s3_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_12_a1_U1 ( .a ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, AdderIns_g2[15]}), .b ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, AdderIns_s3_bc_12_a1_t}), .c ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, AdderIns_g3[15]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, AdderIns_g2[13]}), .b ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, AdderIns_p2[14]}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, AdderIns_s3_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_13_a1_U1 ( .a ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, AdderIns_g2[16]}), .b ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, AdderIns_s3_bc_13_a1_t}), .c ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, AdderIns_g3[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, AdderIns_g2[14]}), .b ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, AdderIns_p2[15]}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, AdderIns_s3_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_14_a1_U1 ( .a ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, AdderIns_g2[17]}), .b ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, AdderIns_s3_bc_14_a1_t}), .c ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, AdderIns_g3[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, AdderIns_g2[15]}), .b ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, AdderIns_p2[16]}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, AdderIns_s3_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_15_a1_U1 ( .a ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, AdderIns_g2[18]}), .b ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, AdderIns_s3_bc_15_a1_t}), .c ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, AdderIns_g3[18]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, AdderIns_g2[16]}), .b ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, AdderIns_p2[17]}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, AdderIns_s3_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_16_a1_U1 ( .a ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, AdderIns_g2[19]}), .b ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, AdderIns_s3_bc_16_a1_t}), .c ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, AdderIns_g3[19]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_16_a1_a1_U1 ( .a ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, AdderIns_g2[17]}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, AdderIns_p2[18]}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, AdderIns_s3_bc_16_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_17_a1_U1 ( .a ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, AdderIns_g2[20]}), .b ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, AdderIns_s3_bc_17_a1_t}), .c ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, AdderIns_g3[20]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_17_a1_a1_U1 ( .a ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, AdderIns_g2[18]}), .b ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, AdderIns_p2[19]}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, AdderIns_s3_bc_17_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_18_a1_U1 ( .a ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, AdderIns_g2[21]}), .b ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, AdderIns_s3_bc_18_a1_t}), .c ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, AdderIns_g3[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_18_a1_a1_U1 ( .a ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, AdderIns_g2[19]}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, AdderIns_p2[20]}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, AdderIns_s3_bc_18_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_19_a1_U1 ( .a ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, AdderIns_g2[22]}), .b ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, AdderIns_s3_bc_19_a1_t}), .c ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, AdderIns_g3[22]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_19_a1_a1_U1 ( .a ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, AdderIns_g2[20]}), .b ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, AdderIns_p2[21]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, AdderIns_s3_bc_19_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_20_a1_U1 ( .a ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, AdderIns_g2[23]}), .b ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, AdderIns_s3_bc_20_a1_t}), .c ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, AdderIns_g3[23]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_20_a1_a1_U1 ( .a ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, AdderIns_g2[21]}), .b ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, AdderIns_p2[22]}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, AdderIns_s3_bc_20_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_21_a1_U1 ( .a ({new_AGEMA_signal_1443, new_AGEMA_signal_1442, AdderIns_g2[24]}), .b ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, AdderIns_s3_bc_21_a1_t}), .c ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, AdderIns_g3[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_21_a1_a1_U1 ( .a ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, AdderIns_g2[22]}), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, AdderIns_p2[23]}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, AdderIns_s3_bc_21_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_22_a1_U1 ( .a ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, AdderIns_g2[25]}), .b ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, AdderIns_s3_bc_22_a1_t}), .c ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, AdderIns_g3[25]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_22_a1_a1_U1 ( .a ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, AdderIns_g2[23]}), .b ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, AdderIns_p2[24]}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, AdderIns_s3_bc_22_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_23_a1_U1 ( .a ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, AdderIns_g2[26]}), .b ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, AdderIns_s3_bc_23_a1_t}), .c ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, AdderIns_g3[26]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_23_a1_a1_U1 ( .a ({new_AGEMA_signal_1443, new_AGEMA_signal_1442, AdderIns_g2[24]}), .b ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, AdderIns_p2[25]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, AdderIns_s3_bc_23_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_24_a1_U1 ( .a ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, AdderIns_g2[27]}), .b ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, AdderIns_s3_bc_24_a1_t}), .c ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, AdderIns_g3[27]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_24_a1_a1_U1 ( .a ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, AdderIns_g2[25]}), .b ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, AdderIns_p2[26]}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, AdderIns_s3_bc_24_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_25_a1_U1 ( .a ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, AdderIns_g2[28]}), .b ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, AdderIns_s3_bc_25_a1_t}), .c ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, AdderIns_g3[28]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_25_a1_a1_U1 ( .a ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, AdderIns_g2[26]}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, AdderIns_p2[27]}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, AdderIns_s3_bc_25_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_26_a1_U1 ( .a ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, AdderIns_g2[29]}), .b ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, AdderIns_s3_bc_26_a1_t}), .c ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, AdderIns_g3[29]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_26_a1_a1_U1 ( .a ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, AdderIns_g2[27]}), .b ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, AdderIns_p2[28]}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, AdderIns_s3_bc_26_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_27_a1_U1 ( .a ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, AdderIns_g2[30]}), .b ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, AdderIns_s3_bc_27_a1_t}), .c ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, AdderIns_g3[30]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s3_bc_27_a1_a1_U1 ( .a ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, AdderIns_g2[28]}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, AdderIns_p2[29]}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, AdderIns_s3_bc_27_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_gc_0_a1_U1 ( .a ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, AdderIns_g3[3]}), .b ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, AdderIns_s4_gc_0_a1_t}), .c ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, AdderIns_g6[3]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, AdderIns_p3[0]}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, AdderIns_s4_gc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_gc_1_a1_U1 ( .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, AdderIns_g3[4]}), .b ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, AdderIns_s4_gc_1_a1_t}), .c ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, AdderIns_g6[4]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, AdderIns_p3[1]}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, AdderIns_s4_gc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_gc_2_a1_U1 ( .a ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, AdderIns_g3[5]}), .b ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, AdderIns_s4_gc_2_a1_t}), .c ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, AdderIns_g6[5]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_gc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, AdderIns_g6[1]}), .b ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, AdderIns_p3[2]}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, AdderIns_s4_gc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_gc_3_a1_U1 ( .a ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, AdderIns_g3[6]}), .b ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, AdderIns_s4_gc_3_a1_t}), .c ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, AdderIns_g6[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_gc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, AdderIns_g6[2]}), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, AdderIns_p3[3]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, AdderIns_s4_gc_3_a1_t}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_0_a2_U1 ( .a ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, AdderIns_p3[0]}), .b ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, AdderIns_p3[4]}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, AdderIns_p4[0]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, AdderIns_p3[1]}), .b ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, AdderIns_p3[5]}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, AdderIns_p4[1]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, AdderIns_p3[2]}), .b ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, AdderIns_p3[6]}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, AdderIns_p4[2]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, AdderIns_p3[3]}), .b ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, AdderIns_p3[7]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, AdderIns_p4[3]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, AdderIns_p3[4]}), .b ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, AdderIns_p3[8]}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, AdderIns_p4[4]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, AdderIns_p3[5]}), .b ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, AdderIns_p3[9]}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, AdderIns_p4[5]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, AdderIns_p3[6]}), .b ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, AdderIns_p3[10]}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, AdderIns_p4[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, AdderIns_p3[7]}), .b ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, AdderIns_p3[11]}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, AdderIns_p4[7]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, AdderIns_p3[8]}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, AdderIns_p3[12]}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, AdderIns_p4[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, AdderIns_p3[9]}), .b ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, AdderIns_p3[13]}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, AdderIns_p4[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, AdderIns_p3[10]}), .b ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, AdderIns_p3[14]}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, AdderIns_p4[10]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, AdderIns_p3[11]}), .b ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, AdderIns_p3[15]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, AdderIns_p4[11]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, AdderIns_p3[12]}), .b ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, AdderIns_p3[16]}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, AdderIns_p4[12]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, AdderIns_p3[13]}), .b ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, AdderIns_p3[17]}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, AdderIns_p4[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, AdderIns_p3[14]}), .b ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, AdderIns_p3[18]}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, AdderIns_p4[14]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_15_a2_U1 ( .a ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, AdderIns_p3[15]}), .b ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, AdderIns_p3[19]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, AdderIns_p4[15]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_16_a2_U1 ( .a ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, AdderIns_p3[16]}), .b ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, AdderIns_p3[20]}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, AdderIns_p4[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_17_a2_U1 ( .a ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, AdderIns_p3[17]}), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, AdderIns_p3[21]}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, AdderIns_p4[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_18_a2_U1 ( .a ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, AdderIns_p3[18]}), .b ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, AdderIns_p3[22]}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, AdderIns_p4[18]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_19_a2_U1 ( .a ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, AdderIns_p3[19]}), .b ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, AdderIns_p3[23]}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, AdderIns_p4[19]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_20_a2_U1 ( .a ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, AdderIns_p3[20]}), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, AdderIns_p3[24]}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, AdderIns_p4[20]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_21_a2_U1 ( .a ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, AdderIns_p3[21]}), .b ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, AdderIns_p3[25]}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, AdderIns_p4[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_22_a2_U1 ( .a ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, AdderIns_p3[22]}), .b ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, AdderIns_p3[26]}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, AdderIns_p4[22]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_23_a2_U1 ( .a ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, AdderIns_p3[23]}), .b ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, AdderIns_p3[27]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, AdderIns_p4[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U29 ( .a ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, AdderIns_g6[6]}), .b ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, AdderIns_p6[7]}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, sum[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U28 ( .a ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, AdderIns_g6[5]}), .b ({new_AGEMA_signal_1119, new_AGEMA_signal_1118, AdderIns_p6[6]}), .c ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, sum[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U27 ( .a ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, AdderIns_g6[4]}), .b ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, AdderIns_p6[5]}), .c ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, sum[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U26 ( .a ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, AdderIns_g6[3]}), .b ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, AdderIns_p6[4]}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, sum[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_15_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, sum[7]}), .a ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, sum[0]}), .c ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, sum_rotated01[15]}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) U130 ( .a ({1'b0, 1'b0, round_constant[10]}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, sum[10]}), .c ({x_round_out_s2[10], x_round_out_s1[10], x_round_out_s0[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U131 ( .a ({1'b0, 1'b0, round_constant[11]}), .b ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, sum[11]}), .c ({x_round_out_s2[11], x_round_out_s1[11], x_round_out_s0[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U132 ( .a ({1'b0, 1'b0, round_constant[12]}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, sum[12]}), .c ({x_round_out_s2[12], x_round_out_s1[12], x_round_out_s0[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U133 ( .a ({1'b0, 1'b0, round_constant[13]}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, sum[13]}), .c ({x_round_out_s2[13], x_round_out_s1[13], x_round_out_s0[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U134 ( .a ({1'b0, 1'b0, round_constant[14]}), .b ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, sum[14]}), .c ({x_round_out_s2[14], x_round_out_s1[14], x_round_out_s0[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U135 ( .a ({1'b0, 1'b0, round_constant[15]}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, sum[15]}), .c ({x_round_out_s2[15], x_round_out_s1[15], x_round_out_s0[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U159 ( .a ({1'b0, 1'b0, round_constant[8]}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, sum[8]}), .c ({x_round_out_s2[8], x_round_out_s1[8], x_round_out_s0[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U160 ( .a ({1'b0, 1'b0, round_constant[9]}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, sum[9]}), .c ({x_round_out_s2[9], x_round_out_s1[9], x_round_out_s0[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U168 ( .a ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, sum_rotated[16]}), .b ({y_round_in_s2[16], y_round_in_s1[16], y_round_in_s0[16]}), .c ({y_round_out_s2[16], y_round_out_s1[16], y_round_out_s0[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_0_a1_U1 ( .a ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, AdderIns_g3[7]}), .b ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, AdderIns_s4_bc_0_a1_t}), .c ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, AdderIns_g4[7]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, AdderIns_g3[3]}), .b ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, AdderIns_p3[4]}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, AdderIns_s4_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_1_a1_U1 ( .a ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, AdderIns_g3[8]}), .b ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, AdderIns_s4_bc_1_a1_t}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, AdderIns_g4[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, AdderIns_g3[4]}), .b ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, AdderIns_p3[5]}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, AdderIns_s4_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_2_a1_U1 ( .a ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, AdderIns_g3[9]}), .b ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, AdderIns_s4_bc_2_a1_t}), .c ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, AdderIns_g4[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, AdderIns_g3[5]}), .b ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, AdderIns_p3[6]}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, AdderIns_s4_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_3_a1_U1 ( .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, AdderIns_g3[10]}), .b ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, AdderIns_s4_bc_3_a1_t}), .c ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, AdderIns_g4[10]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, AdderIns_g3[6]}), .b ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, AdderIns_p3[7]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, AdderIns_s4_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_4_a1_U1 ( .a ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, AdderIns_g3[11]}), .b ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, AdderIns_s4_bc_4_a1_t}), .c ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, AdderIns_g4[11]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, AdderIns_g3[7]}), .b ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, AdderIns_p3[8]}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, AdderIns_s4_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_5_a1_U1 ( .a ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, AdderIns_g3[12]}), .b ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, AdderIns_s4_bc_5_a1_t}), .c ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, AdderIns_g4[12]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, AdderIns_g3[8]}), .b ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, AdderIns_p3[9]}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, AdderIns_s4_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_6_a1_U1 ( .a ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, AdderIns_g3[13]}), .b ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, AdderIns_s4_bc_6_a1_t}), .c ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, AdderIns_g4[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, AdderIns_g3[9]}), .b ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, AdderIns_p3[10]}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, AdderIns_s4_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_7_a1_U1 ( .a ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, AdderIns_g3[14]}), .b ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, AdderIns_s4_bc_7_a1_t}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, AdderIns_g4[14]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, AdderIns_g3[10]}), .b ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, AdderIns_p3[11]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, AdderIns_s4_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_8_a1_U1 ( .a ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, AdderIns_g3[15]}), .b ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, AdderIns_s4_bc_8_a1_t}), .c ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, AdderIns_g4[15]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, AdderIns_g3[11]}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, AdderIns_p3[12]}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, AdderIns_s4_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_9_a1_U1 ( .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, AdderIns_g3[16]}), .b ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, AdderIns_s4_bc_9_a1_t}), .c ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, AdderIns_g4[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, AdderIns_g3[12]}), .b ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, AdderIns_p3[13]}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, AdderIns_s4_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_10_a1_U1 ( .a ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, AdderIns_g3[17]}), .b ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, AdderIns_s4_bc_10_a1_t}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, AdderIns_g4[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, AdderIns_g3[13]}), .b ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, AdderIns_p3[14]}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, AdderIns_s4_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_11_a1_U1 ( .a ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, AdderIns_g3[18]}), .b ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, AdderIns_s4_bc_11_a1_t}), .c ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, AdderIns_g4[18]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, AdderIns_g3[14]}), .b ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, AdderIns_p3[15]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, AdderIns_s4_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_12_a1_U1 ( .a ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, AdderIns_g3[19]}), .b ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, AdderIns_s4_bc_12_a1_t}), .c ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, AdderIns_g4[19]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, AdderIns_g3[15]}), .b ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, AdderIns_p3[16]}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, AdderIns_s4_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_13_a1_U1 ( .a ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, AdderIns_g3[20]}), .b ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, AdderIns_s4_bc_13_a1_t}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, AdderIns_g4[20]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, AdderIns_g3[16]}), .b ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, AdderIns_p3[17]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, AdderIns_s4_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_14_a1_U1 ( .a ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, AdderIns_g3[21]}), .b ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, AdderIns_s4_bc_14_a1_t}), .c ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, AdderIns_g4[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, AdderIns_g3[17]}), .b ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, AdderIns_p3[18]}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, AdderIns_s4_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_15_a1_U1 ( .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, AdderIns_g3[22]}), .b ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, AdderIns_s4_bc_15_a1_t}), .c ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, AdderIns_g4[22]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, AdderIns_g3[18]}), .b ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, AdderIns_p3[19]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, AdderIns_s4_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_16_a1_U1 ( .a ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, AdderIns_g3[23]}), .b ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, AdderIns_s4_bc_16_a1_t}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, AdderIns_g4[23]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_16_a1_a1_U1 ( .a ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, AdderIns_g3[19]}), .b ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, AdderIns_p3[20]}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, AdderIns_s4_bc_16_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_17_a1_U1 ( .a ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, AdderIns_g3[24]}), .b ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, AdderIns_s4_bc_17_a1_t}), .c ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, AdderIns_g4[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_17_a1_a1_U1 ( .a ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, AdderIns_g3[20]}), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, AdderIns_p3[21]}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, AdderIns_s4_bc_17_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_18_a1_U1 ( .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, AdderIns_g3[25]}), .b ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, AdderIns_s4_bc_18_a1_t}), .c ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, AdderIns_g4[25]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_18_a1_a1_U1 ( .a ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, AdderIns_g3[21]}), .b ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, AdderIns_p3[22]}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, AdderIns_s4_bc_18_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_19_a1_U1 ( .a ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, AdderIns_g3[26]}), .b ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, AdderIns_s4_bc_19_a1_t}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, AdderIns_g4[26]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_19_a1_a1_U1 ( .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, AdderIns_g3[22]}), .b ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, AdderIns_p3[23]}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, AdderIns_s4_bc_19_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_20_a1_U1 ( .a ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, AdderIns_g3[27]}), .b ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, AdderIns_s4_bc_20_a1_t}), .c ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, AdderIns_g4[27]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_20_a1_a1_U1 ( .a ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, AdderIns_g3[23]}), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, AdderIns_p3[24]}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, AdderIns_s4_bc_20_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_21_a1_U1 ( .a ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, AdderIns_g3[28]}), .b ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, AdderIns_s4_bc_21_a1_t}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, AdderIns_g4[28]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_21_a1_a1_U1 ( .a ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, AdderIns_g3[24]}), .b ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, AdderIns_p3[25]}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, AdderIns_s4_bc_21_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_22_a1_U1 ( .a ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, AdderIns_g3[29]}), .b ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, AdderIns_s4_bc_22_a1_t}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, AdderIns_g4[29]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_22_a1_a1_U1 ( .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, AdderIns_g3[25]}), .b ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, AdderIns_p3[26]}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, AdderIns_s4_bc_22_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_23_a1_U1 ( .a ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, AdderIns_g3[30]}), .b ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, AdderIns_s4_bc_23_a1_t}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, AdderIns_g4[30]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s4_bc_23_a1_a1_U1 ( .a ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, AdderIns_g3[26]}), .b ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, AdderIns_p3[27]}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, AdderIns_s4_bc_23_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_0_a1_U1 ( .a ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, AdderIns_g4[7]}), .b ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, AdderIns_s5_gc_0_a1_t}), .c ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, AdderIns_g6[7]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, AdderIns_p4[0]}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, AdderIns_s5_gc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_1_a1_U1 ( .a ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, AdderIns_g4[8]}), .b ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, AdderIns_s5_gc_1_a1_t}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, AdderIns_g6[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, AdderIns_p4[1]}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, AdderIns_s5_gc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_2_a1_U1 ( .a ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, AdderIns_g4[9]}), .b ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, AdderIns_s5_gc_2_a1_t}), .c ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, AdderIns_g6[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, AdderIns_g6[1]}), .b ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, AdderIns_p4[2]}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, AdderIns_s5_gc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_3_a1_U1 ( .a ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, AdderIns_g4[10]}), .b ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, AdderIns_s5_gc_3_a1_t}), .c ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, AdderIns_g6[10]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, AdderIns_g6[2]}), .b ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, AdderIns_p4[3]}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, AdderIns_s5_gc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_4_a1_U1 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, AdderIns_g4[11]}), .b ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, AdderIns_s5_gc_4_a1_t}), .c ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, AdderIns_g6[11]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, AdderIns_g6[3]}), .b ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, AdderIns_p4[4]}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, AdderIns_s5_gc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_5_a1_U1 ( .a ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, AdderIns_g4[12]}), .b ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, AdderIns_s5_gc_5_a1_t}), .c ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, AdderIns_g6[12]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, AdderIns_g6[4]}), .b ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, AdderIns_p4[5]}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, AdderIns_s5_gc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_6_a1_U1 ( .a ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, AdderIns_g4[13]}), .b ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, AdderIns_s5_gc_6_a1_t}), .c ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, AdderIns_g6[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, AdderIns_g6[5]}), .b ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, AdderIns_p4[6]}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, AdderIns_s5_gc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_7_a1_U1 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, AdderIns_g4[14]}), .b ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, AdderIns_s5_gc_7_a1_t}), .c ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, AdderIns_g6[14]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_gc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, AdderIns_g6[6]}), .b ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, AdderIns_p4[7]}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, AdderIns_s5_gc_7_a1_t}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, AdderIns_p4[1]}), .b ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, AdderIns_p4[9]}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, AdderIns_p5[1]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, AdderIns_p4[2]}), .b ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, AdderIns_p4[10]}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, AdderIns_p5[2]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, AdderIns_p4[3]}), .b ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, AdderIns_p4[11]}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, AdderIns_p5[3]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, AdderIns_p4[4]}), .b ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, AdderIns_p4[12]}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, AdderIns_p5[4]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, AdderIns_p4[5]}), .b ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, AdderIns_p4[13]}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, AdderIns_p5[5]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, AdderIns_p4[6]}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, AdderIns_p4[14]}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, AdderIns_p5[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, AdderIns_p4[7]}), .b ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, AdderIns_p4[15]}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, AdderIns_p5[7]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, AdderIns_p4[8]}), .b ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, AdderIns_p4[16]}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, AdderIns_p5[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, AdderIns_p4[9]}), .b ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, AdderIns_p4[17]}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, AdderIns_p5[9]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, AdderIns_p4[10]}), .b ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, AdderIns_p4[18]}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, AdderIns_p5[10]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, AdderIns_p4[11]}), .b ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, AdderIns_p4[19]}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, AdderIns_p5[11]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, AdderIns_p4[12]}), .b ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, AdderIns_p4[20]}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, AdderIns_p5[12]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, AdderIns_p4[13]}), .b ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, AdderIns_p4[21]}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, AdderIns_p5[13]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, AdderIns_p4[14]}), .b ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, AdderIns_p4[22]}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, AdderIns_p5[14]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_15_a2_U1 ( .a ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, AdderIns_p4[15]}), .b ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, AdderIns_p4[23]}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, AdderIns_p5[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U31 ( .a ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, AdderIns_g6[8]}), .b ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, AdderIns_p6[9]}), .c ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, sum[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U30 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, AdderIns_g6[7]}), .b ({new_AGEMA_signal_1131, new_AGEMA_signal_1130, AdderIns_p6[8]}), .c ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, sum[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U6 ( .a ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, AdderIns_g6[14]}), .b ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, AdderIns_p6[15]}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, sum[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U5 ( .a ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, AdderIns_g6[13]}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, AdderIns_p6[14]}), .c ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, sum[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U4 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, AdderIns_g6[12]}), .b ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, AdderIns_p6[13]}), .c ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, sum[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U3 ( .a ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, AdderIns_g6[11]}), .b ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, AdderIns_p6[12]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, sum[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U2 ( .a ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, AdderIns_g6[10]}), .b ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, AdderIns_p6[11]}), .c ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, sum[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U1 ( .a ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, AdderIns_g6[9]}), .b ({new_AGEMA_signal_1143, new_AGEMA_signal_1142, AdderIns_p6[10]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, sum[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_16_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, sum[8]}), .a ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, sum[1]}), .c ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, sum_rotated01[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_17_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, sum[9]}), .a ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, sum[2]}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, sum_rotated01[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_18_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, sum[10]}), .a ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, sum[3]}), .c ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, sum_rotated01[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_19_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, sum[11]}), .a ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, sum[4]}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, sum_rotated01[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_20_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, sum[12]}), .a ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, sum[5]}), .c ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, sum_rotated01[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_21_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, sum[13]}), .a ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, sum[6]}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, sum_rotated01[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_22_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, sum[14]}), .a ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, sum[7]}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, sum_rotated01[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_23_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, sum[15]}), .a ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, sum[8]}), .c ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, sum_rotated01[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_16_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, sum[15]}), .a ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, sum[0]}), .c ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, sum_rotated23[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_16_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, sum_rotated01[16]}), .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, sum_rotated23[16]}), .c ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, sum_rotated[16]}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) U136 ( .a ({1'b0, 1'b0, round_constant[16]}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, sum[16]}), .c ({x_round_out_s2[16], x_round_out_s1[16], x_round_out_s0[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U137 ( .a ({1'b0, 1'b0, round_constant[17]}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, sum[17]}), .c ({x_round_out_s2[17], x_round_out_s1[17], x_round_out_s0[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U138 ( .a ({1'b0, 1'b0, round_constant[18]}), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, sum[18]}), .c ({x_round_out_s2[18], x_round_out_s1[18], x_round_out_s0[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U139 ( .a ({1'b0, 1'b0, round_constant[19]}), .b ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, sum[19]}), .c ({x_round_out_s2[19], x_round_out_s1[19], x_round_out_s0[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U141 ( .a ({1'b0, 1'b0, round_constant[20]}), .b ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, sum[20]}), .c ({x_round_out_s2[20], x_round_out_s1[20], x_round_out_s0[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U142 ( .a ({1'b0, 1'b0, round_constant[21]}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, sum[21]}), .c ({x_round_out_s2[21], x_round_out_s1[21], x_round_out_s0[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U143 ( .a ({1'b0, 1'b0, round_constant[22]}), .b ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, sum[22]}), .c ({x_round_out_s2[22], x_round_out_s1[22], x_round_out_s0[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U144 ( .a ({1'b0, 1'b0, round_constant[23]}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, sum[23]}), .c ({x_round_out_s2[23], x_round_out_s1[23], x_round_out_s0[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U145 ( .a ({1'b0, 1'b0, round_constant[24]}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, sum[24]}), .c ({x_round_out_s2[24], x_round_out_s1[24], x_round_out_s0[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U146 ( .a ({1'b0, 1'b0, round_constant[25]}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, sum[25]}), .c ({x_round_out_s2[25], x_round_out_s1[25], x_round_out_s0[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U147 ( .a ({1'b0, 1'b0, round_constant[26]}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, sum[26]}), .c ({x_round_out_s2[26], x_round_out_s1[26], x_round_out_s0[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U148 ( .a ({1'b0, 1'b0, round_constant[27]}), .b ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, sum[27]}), .c ({x_round_out_s2[27], x_round_out_s1[27], x_round_out_s0[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U149 ( .a ({1'b0, 1'b0, round_constant[28]}), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, sum[28]}), .c ({x_round_out_s2[28], x_round_out_s1[28], x_round_out_s0[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U150 ( .a ({1'b0, 1'b0, round_constant[29]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, sum[29]}), .c ({x_round_out_s2[29], x_round_out_s1[29], x_round_out_s0[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U152 ( .a ({1'b0, 1'b0, round_constant[30]}), .b ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, sum[30]}), .c ({x_round_out_s2[30], x_round_out_s1[30], x_round_out_s0[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U153 ( .a ({1'b0, 1'b0, round_constant[31]}), .b ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, sum[31]}), .c ({x_round_out_s2[31], x_round_out_s1[31], x_round_out_s0[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U161 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, sum_rotated[0]}), .b ({y_round_in_s2[0], y_round_in_s1[0], y_round_in_s0[0]}), .c ({y_round_out_s2[0], y_round_out_s1[0], y_round_out_s0[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U162 ( .a ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, sum_rotated[10]}), .b ({y_round_in_s2[10], y_round_in_s1[10], y_round_in_s0[10]}), .c ({y_round_out_s2[10], y_round_out_s1[10], y_round_out_s0[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U163 ( .a ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, sum_rotated[11]}), .b ({y_round_in_s2[11], y_round_in_s1[11], y_round_in_s0[11]}), .c ({y_round_out_s2[11], y_round_out_s1[11], y_round_out_s0[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U164 ( .a ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, sum_rotated[12]}), .b ({y_round_in_s2[12], y_round_in_s1[12], y_round_in_s0[12]}), .c ({y_round_out_s2[12], y_round_out_s1[12], y_round_out_s0[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U165 ( .a ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, sum_rotated[13]}), .b ({y_round_in_s2[13], y_round_in_s1[13], y_round_in_s0[13]}), .c ({y_round_out_s2[13], y_round_out_s1[13], y_round_out_s0[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U166 ( .a ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, sum_rotated[14]}), .b ({y_round_in_s2[14], y_round_in_s1[14], y_round_in_s0[14]}), .c ({y_round_out_s2[14], y_round_out_s1[14], y_round_out_s0[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U167 ( .a ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, sum_rotated[15]}), .b ({y_round_in_s2[15], y_round_in_s1[15], y_round_in_s0[15]}), .c ({y_round_out_s2[15], y_round_out_s1[15], y_round_out_s0[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U169 ( .a ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, sum_rotated[17]}), .b ({y_round_in_s2[17], y_round_in_s1[17], y_round_in_s0[17]}), .c ({y_round_out_s2[17], y_round_out_s1[17], y_round_out_s0[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U170 ( .a ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, sum_rotated[18]}), .b ({y_round_in_s2[18], y_round_in_s1[18], y_round_in_s0[18]}), .c ({y_round_out_s2[18], y_round_out_s1[18], y_round_out_s0[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U171 ( .a ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, sum_rotated[19]}), .b ({y_round_in_s2[19], y_round_in_s1[19], y_round_in_s0[19]}), .c ({y_round_out_s2[19], y_round_out_s1[19], y_round_out_s0[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U172 ( .a ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, sum_rotated[1]}), .b ({y_round_in_s2[1], y_round_in_s1[1], y_round_in_s0[1]}), .c ({y_round_out_s2[1], y_round_out_s1[1], y_round_out_s0[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U173 ( .a ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, sum_rotated[20]}), .b ({y_round_in_s2[20], y_round_in_s1[20], y_round_in_s0[20]}), .c ({y_round_out_s2[20], y_round_out_s1[20], y_round_out_s0[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U174 ( .a ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, sum_rotated[21]}), .b ({y_round_in_s2[21], y_round_in_s1[21], y_round_in_s0[21]}), .c ({y_round_out_s2[21], y_round_out_s1[21], y_round_out_s0[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U175 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, sum_rotated[22]}), .b ({y_round_in_s2[22], y_round_in_s1[22], y_round_in_s0[22]}), .c ({y_round_out_s2[22], y_round_out_s1[22], y_round_out_s0[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U176 ( .a ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, sum_rotated[23]}), .b ({y_round_in_s2[23], y_round_in_s1[23], y_round_in_s0[23]}), .c ({y_round_out_s2[23], y_round_out_s1[23], y_round_out_s0[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U177 ( .a ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, sum_rotated[24]}), .b ({y_round_in_s2[24], y_round_in_s1[24], y_round_in_s0[24]}), .c ({y_round_out_s2[24], y_round_out_s1[24], y_round_out_s0[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U178 ( .a ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, sum_rotated[25]}), .b ({y_round_in_s2[25], y_round_in_s1[25], y_round_in_s0[25]}), .c ({y_round_out_s2[25], y_round_out_s1[25], y_round_out_s0[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U179 ( .a ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, sum_rotated[26]}), .b ({y_round_in_s2[26], y_round_in_s1[26], y_round_in_s0[26]}), .c ({y_round_out_s2[26], y_round_out_s1[26], y_round_out_s0[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U180 ( .a ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, sum_rotated[27]}), .b ({y_round_in_s2[27], y_round_in_s1[27], y_round_in_s0[27]}), .c ({y_round_out_s2[27], y_round_out_s1[27], y_round_out_s0[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U181 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, sum_rotated[28]}), .b ({y_round_in_s2[28], y_round_in_s1[28], y_round_in_s0[28]}), .c ({y_round_out_s2[28], y_round_out_s1[28], y_round_out_s0[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U182 ( .a ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, sum_rotated[29]}), .b ({y_round_in_s2[29], y_round_in_s1[29], y_round_in_s0[29]}), .c ({y_round_out_s2[29], y_round_out_s1[29], y_round_out_s0[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U183 ( .a ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, sum_rotated[2]}), .b ({y_round_in_s2[2], y_round_in_s1[2], y_round_in_s0[2]}), .c ({y_round_out_s2[2], y_round_out_s1[2], y_round_out_s0[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U184 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, sum_rotated[30]}), .b ({y_round_in_s2[30], y_round_in_s1[30], y_round_in_s0[30]}), .c ({y_round_out_s2[30], y_round_out_s1[30], y_round_out_s0[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U185 ( .a ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, sum_rotated[31]}), .b ({y_round_in_s2[31], y_round_in_s1[31], y_round_in_s0[31]}), .c ({y_round_out_s2[31], y_round_out_s1[31], y_round_out_s0[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U186 ( .a ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, sum_rotated[3]}), .b ({y_round_in_s2[3], y_round_in_s1[3], y_round_in_s0[3]}), .c ({y_round_out_s2[3], y_round_out_s1[3], y_round_out_s0[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U187 ( .a ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, sum_rotated[4]}), .b ({y_round_in_s2[4], y_round_in_s1[4], y_round_in_s0[4]}), .c ({y_round_out_s2[4], y_round_out_s1[4], y_round_out_s0[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U188 ( .a ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, sum_rotated[5]}), .b ({y_round_in_s2[5], y_round_in_s1[5], y_round_in_s0[5]}), .c ({y_round_out_s2[5], y_round_out_s1[5], y_round_out_s0[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U189 ( .a ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, sum_rotated[6]}), .b ({y_round_in_s2[6], y_round_in_s1[6], y_round_in_s0[6]}), .c ({y_round_out_s2[6], y_round_out_s1[6], y_round_out_s0[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U190 ( .a ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, sum_rotated[7]}), .b ({y_round_in_s2[7], y_round_in_s1[7], y_round_in_s0[7]}), .c ({y_round_out_s2[7], y_round_out_s1[7], y_round_out_s0[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U191 ( .a ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, sum_rotated[8]}), .b ({y_round_in_s2[8], y_round_in_s1[8], y_round_in_s0[8]}), .c ({y_round_out_s2[8], y_round_out_s1[8], y_round_out_s0[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U192 ( .a ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, sum_rotated[9]}), .b ({y_round_in_s2[9], y_round_in_s1[9], y_round_in_s0[9]}), .c ({y_round_out_s2[9], y_round_out_s1[9], y_round_out_s0[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_0_a1_U1 ( .a ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, AdderIns_g4[15]}), .b ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, AdderIns_s5_bc_0_a1_t}), .c ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, AdderIns_g6[15]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, AdderIns_g4[7]}), .b ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, AdderIns_p4[8]}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, AdderIns_s5_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_1_a1_U1 ( .a ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, AdderIns_g4[16]}), .b ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, AdderIns_s5_bc_1_a1_t}), .c ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, AdderIns_g5[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, AdderIns_g4[8]}), .b ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, AdderIns_p4[9]}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, AdderIns_s5_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_2_a1_U1 ( .a ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, AdderIns_g4[17]}), .b ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, AdderIns_s5_bc_2_a1_t}), .c ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, AdderIns_g5[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, AdderIns_g4[9]}), .b ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, AdderIns_p4[10]}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, AdderIns_s5_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_3_a1_U1 ( .a ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, AdderIns_g4[18]}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, AdderIns_s5_bc_3_a1_t}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, AdderIns_g5[18]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, AdderIns_g4[10]}), .b ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, AdderIns_p4[11]}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, AdderIns_s5_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_4_a1_U1 ( .a ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, AdderIns_g4[19]}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, AdderIns_s5_bc_4_a1_t}), .c ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, AdderIns_g5[19]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, AdderIns_g4[11]}), .b ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, AdderIns_p4[12]}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, AdderIns_s5_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_5_a1_U1 ( .a ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, AdderIns_g4[20]}), .b ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, AdderIns_s5_bc_5_a1_t}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, AdderIns_g5[20]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, AdderIns_g4[12]}), .b ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, AdderIns_p4[13]}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, AdderIns_s5_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_6_a1_U1 ( .a ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, AdderIns_g4[21]}), .b ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, AdderIns_s5_bc_6_a1_t}), .c ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, AdderIns_g5[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, AdderIns_g4[13]}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, AdderIns_p4[14]}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, AdderIns_s5_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_7_a1_U1 ( .a ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, AdderIns_g4[22]}), .b ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, AdderIns_s5_bc_7_a1_t}), .c ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, AdderIns_g5[22]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, AdderIns_g4[14]}), .b ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, AdderIns_p4[15]}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, AdderIns_s5_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_8_a1_U1 ( .a ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, AdderIns_g4[23]}), .b ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, AdderIns_s5_bc_8_a1_t}), .c ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, AdderIns_g5[23]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, AdderIns_g4[15]}), .b ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, AdderIns_p4[16]}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, AdderIns_s5_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_9_a1_U1 ( .a ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, AdderIns_g4[24]}), .b ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, AdderIns_s5_bc_9_a1_t}), .c ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, AdderIns_g5[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, AdderIns_g4[16]}), .b ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, AdderIns_p4[17]}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, AdderIns_s5_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_10_a1_U1 ( .a ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, AdderIns_g4[25]}), .b ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, AdderIns_s5_bc_10_a1_t}), .c ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, AdderIns_g5[25]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, AdderIns_g4[17]}), .b ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, AdderIns_p4[18]}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, AdderIns_s5_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_11_a1_U1 ( .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, AdderIns_g4[26]}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, AdderIns_s5_bc_11_a1_t}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, AdderIns_g5[26]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, AdderIns_g4[18]}), .b ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, AdderIns_p4[19]}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, AdderIns_s5_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_12_a1_U1 ( .a ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, AdderIns_g4[27]}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, AdderIns_s5_bc_12_a1_t}), .c ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, AdderIns_g5[27]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, AdderIns_g4[19]}), .b ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, AdderIns_p4[20]}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, AdderIns_s5_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_13_a1_U1 ( .a ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, AdderIns_g4[28]}), .b ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, AdderIns_s5_bc_13_a1_t}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, AdderIns_g5[28]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, AdderIns_g4[20]}), .b ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, AdderIns_p4[21]}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, AdderIns_s5_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_14_a1_U1 ( .a ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, AdderIns_g4[29]}), .b ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, AdderIns_s5_bc_14_a1_t}), .c ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, AdderIns_g5[29]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, AdderIns_g4[21]}), .b ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, AdderIns_p4[22]}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, AdderIns_s5_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_15_a1_U1 ( .a ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, AdderIns_g4[30]}), .b ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, AdderIns_s5_bc_15_a1_t}), .c ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, AdderIns_g5[30]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s5_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, AdderIns_g4[22]}), .b ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, AdderIns_p4[23]}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, AdderIns_s5_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_1_a1_U1 ( .a ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, AdderIns_g5[16]}), .b ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, AdderIns_s6_gc_1_a1_t}), .c ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, AdderIns_g6[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, AdderIns_p5[1]}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, AdderIns_s6_gc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_2_a1_U1 ( .a ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, AdderIns_g5[17]}), .b ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, AdderIns_s6_gc_2_a1_t}), .c ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, AdderIns_g6[17]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, AdderIns_g6[1]}), .b ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, AdderIns_p5[2]}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, AdderIns_s6_gc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_3_a1_U1 ( .a ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, AdderIns_g5[18]}), .b ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, AdderIns_s6_gc_3_a1_t}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, AdderIns_g6[18]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, AdderIns_g6[2]}), .b ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, AdderIns_p5[3]}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, AdderIns_s6_gc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_4_a1_U1 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, AdderIns_g5[19]}), .b ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, AdderIns_s6_gc_4_a1_t}), .c ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, AdderIns_g6[19]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, AdderIns_g6[3]}), .b ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, AdderIns_p5[4]}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, AdderIns_s6_gc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_5_a1_U1 ( .a ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, AdderIns_g5[20]}), .b ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, AdderIns_s6_gc_5_a1_t}), .c ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, AdderIns_g6[20]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, AdderIns_g6[4]}), .b ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, AdderIns_p5[5]}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, AdderIns_s6_gc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_6_a1_U1 ( .a ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, AdderIns_g5[21]}), .b ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, AdderIns_s6_gc_6_a1_t}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, AdderIns_g6[21]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, AdderIns_g6[5]}), .b ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, AdderIns_p5[6]}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, AdderIns_s6_gc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_7_a1_U1 ( .a ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, AdderIns_g5[22]}), .b ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, AdderIns_s6_gc_7_a1_t}), .c ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, AdderIns_g6[22]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, AdderIns_g6[6]}), .b ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, AdderIns_p5[7]}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, AdderIns_s6_gc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_8_a1_U1 ( .a ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, AdderIns_g5[23]}), .b ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, AdderIns_s6_gc_8_a1_t}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, AdderIns_g6[23]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, AdderIns_g6[7]}), .b ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, AdderIns_p5[8]}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, AdderIns_s6_gc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_9_a1_U1 ( .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, AdderIns_g5[24]}), .b ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, AdderIns_s6_gc_9_a1_t}), .c ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, AdderIns_g6[24]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, AdderIns_g6[8]}), .b ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, AdderIns_p5[9]}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, AdderIns_s6_gc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_10_a1_U1 ( .a ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, AdderIns_g5[25]}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, AdderIns_s6_gc_10_a1_t}), .c ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, AdderIns_g6[25]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, AdderIns_g6[9]}), .b ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, AdderIns_p5[10]}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, AdderIns_s6_gc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_11_a1_U1 ( .a ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, AdderIns_g5[26]}), .b ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, AdderIns_s6_gc_11_a1_t}), .c ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, AdderIns_g6[26]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, AdderIns_g6[10]}), .b ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, AdderIns_p5[11]}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, AdderIns_s6_gc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_12_a1_U1 ( .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, AdderIns_g5[27]}), .b ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, AdderIns_s6_gc_12_a1_t}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, AdderIns_g6[27]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, AdderIns_g6[11]}), .b ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, AdderIns_p5[12]}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, AdderIns_s6_gc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_13_a1_U1 ( .a ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, AdderIns_g5[28]}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, AdderIns_s6_gc_13_a1_t}), .c ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, AdderIns_g6[28]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, AdderIns_g6[12]}), .b ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, AdderIns_p5[13]}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, AdderIns_s6_gc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_14_a1_U1 ( .a ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, AdderIns_g5[29]}), .b ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, AdderIns_s6_gc_14_a1_t}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, AdderIns_g6[29]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, AdderIns_g6[13]}), .b ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, AdderIns_p5[14]}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, AdderIns_s6_gc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_15_a1_U1 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, AdderIns_g5[30]}), .b ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, AdderIns_s6_gc_15_a1_t}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, AdderIns_g6[30]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s6_gc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, AdderIns_g6[14]}), .b ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, AdderIns_p5[15]}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, AdderIns_s6_gc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U24 ( .a ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, AdderIns_g6[30]}), .b ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, AdderIns_p6[31]}), .c ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, sum[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U23 ( .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, AdderIns_g6[29]}), .b ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, AdderIns_p6[30]}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, sum[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U21 ( .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, AdderIns_g6[28]}), .b ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, AdderIns_p6[29]}), .c ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, sum[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U20 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, AdderIns_g6[27]}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, AdderIns_p6[28]}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, sum[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U19 ( .a ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, AdderIns_g6[26]}), .b ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, AdderIns_p6[27]}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, sum[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U18 ( .a ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, AdderIns_g6[25]}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, AdderIns_p6[26]}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, sum[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U17 ( .a ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, AdderIns_g6[24]}), .b ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, AdderIns_p6[25]}), .c ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, sum[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U16 ( .a ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, AdderIns_g6[23]}), .b ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, AdderIns_p6[24]}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, sum[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U15 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, AdderIns_g6[22]}), .b ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, AdderIns_p6[23]}), .c ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, sum[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U14 ( .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, AdderIns_g6[21]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, AdderIns_p6[22]}), .c ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, sum[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U13 ( .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, AdderIns_g6[20]}), .b ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, AdderIns_p6[21]}), .c ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, sum[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U12 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, AdderIns_g6[19]}), .b ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, AdderIns_p6[20]}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, sum[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U10 ( .a ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, AdderIns_g6[18]}), .b ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, AdderIns_p6[19]}), .c ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, sum[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U9 ( .a ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, AdderIns_g6[17]}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, AdderIns_p6[18]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, sum[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U8 ( .a ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, AdderIns_g6[16]}), .b ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, AdderIns_p6[17]}), .c ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, sum[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) AdderIns_s7_U7 ( .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, AdderIns_g6[15]}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, AdderIns_p6[16]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, sum[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_0_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, sum[24]}), .a ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, sum[17]}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, sum_rotated01[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_1_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, sum[25]}), .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, sum[18]}), .c ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, sum_rotated01[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_2_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, sum[26]}), .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, sum[19]}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, sum_rotated01[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_3_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, sum[27]}), .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, sum[20]}), .c ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, sum_rotated01[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_4_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, sum[28]}), .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, sum[21]}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, sum_rotated01[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_5_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, sum[29]}), .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, sum[22]}), .c ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, sum_rotated01[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_6_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, sum[30]}), .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, sum[23]}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, sum_rotated01[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_7_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, sum[31]}), .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, sum[24]}), .c ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, sum_rotated01[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_8_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, sum[0]}), .a ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, sum[25]}), .c ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, sum_rotated01[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_9_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, sum[1]}), .a ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, sum[26]}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, sum_rotated01[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_10_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, sum[2]}), .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, sum[27]}), .c ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, sum_rotated01[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_11_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, sum[3]}), .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, sum[28]}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, sum_rotated01[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_12_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, sum[4]}), .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, sum[29]}), .c ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, sum_rotated01[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_13_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, sum[5]}), .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, sum[30]}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, sum_rotated01[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_14_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, sum[6]}), .a ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, sum[31]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, sum_rotated01[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_24_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, sum[16]}), .a ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, sum[9]}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, sum_rotated01[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_25_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, sum[17]}), .a ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, sum[10]}), .c ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, sum_rotated01[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_26_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, sum[18]}), .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, sum[11]}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, sum_rotated01[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_27_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, sum[19]}), .a ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, sum[12]}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, sum_rotated01[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_28_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, sum[20]}), .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, sum[13]}), .c ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, sum_rotated01[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_29_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, sum[21]}), .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, sum[14]}), .c ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, sum_rotated01[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_30_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, sum[22]}), .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, sum[15]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, sum_rotated01[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M4_mux_inst_31_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, sum[23]}), .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, sum[16]}), .c ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, sum_rotated01[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_0_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, sum[31]}), .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, sum[16]}), .c ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, sum_rotated23[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_1_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, sum[0]}), .a ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, sum[17]}), .c ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, sum_rotated23[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_2_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, sum[1]}), .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, sum[18]}), .c ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, sum_rotated23[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_3_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, sum[2]}), .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, sum[19]}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, sum_rotated23[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_4_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, sum[3]}), .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, sum[20]}), .c ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, sum_rotated23[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_5_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, sum[4]}), .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, sum[21]}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, sum_rotated23[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_6_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, sum[5]}), .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, sum[22]}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, sum_rotated23[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_7_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, sum[6]}), .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, sum[23]}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, sum_rotated23[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_8_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, sum[7]}), .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, sum[24]}), .c ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, sum_rotated23[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_9_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, sum[8]}), .a ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, sum[25]}), .c ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, sum_rotated23[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_10_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, sum[9]}), .a ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, sum[26]}), .c ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, sum_rotated23[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_11_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, sum[10]}), .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, sum[27]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, sum_rotated23[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_12_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, sum[11]}), .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, sum[28]}), .c ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, sum_rotated23[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_13_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, sum[12]}), .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, sum[29]}), .c ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, sum_rotated23[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_14_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, sum[13]}), .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, sum[30]}), .c ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, sum_rotated23[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_15_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, sum[14]}), .a ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, sum[31]}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, sum_rotated23[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_17_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, sum[16]}), .a ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, sum[1]}), .c ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, sum_rotated23[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_18_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, sum[17]}), .a ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, sum[2]}), .c ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, sum_rotated23[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_19_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, sum[18]}), .a ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, sum[3]}), .c ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, sum_rotated23[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_20_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, sum[19]}), .a ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, sum[4]}), .c ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, sum_rotated23[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_21_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, sum[20]}), .a ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, sum[5]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, sum_rotated23[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_22_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, sum[21]}), .a ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, sum[6]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, sum_rotated23[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_23_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, sum[22]}), .a ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, sum[7]}), .c ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, sum_rotated23[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_24_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, sum[23]}), .a ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, sum[8]}), .c ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, sum_rotated23[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_25_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, sum[24]}), .a ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, sum[9]}), .c ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, sum_rotated23[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_26_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, sum[25]}), .a ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, sum[10]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, sum_rotated23[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_27_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, sum[26]}), .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, sum[11]}), .c ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, sum_rotated23[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_28_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, sum[27]}), .a ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, sum[12]}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, sum_rotated23[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_29_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, sum[28]}), .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, sum[13]}), .c ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, sum_rotated23[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_30_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, sum[29]}), .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, sum[14]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, sum_rotated23[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M5_mux_inst_31_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, sum[30]}), .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, sum[15]}), .c ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, sum_rotated23[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_0_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, sum_rotated01[0]}), .a ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, sum_rotated23[0]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, sum_rotated[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_1_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, sum_rotated01[1]}), .a ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, sum_rotated23[1]}), .c ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, sum_rotated[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_2_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, sum_rotated01[2]}), .a ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, sum_rotated23[2]}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, sum_rotated[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_3_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, sum_rotated01[3]}), .a ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, sum_rotated23[3]}), .c ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, sum_rotated[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_4_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, sum_rotated01[4]}), .a ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, sum_rotated23[4]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, sum_rotated[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_5_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, sum_rotated01[5]}), .a ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, sum_rotated23[5]}), .c ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, sum_rotated[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_6_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, sum_rotated01[6]}), .a ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, sum_rotated23[6]}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, sum_rotated[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_7_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, sum_rotated01[7]}), .a ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, sum_rotated23[7]}), .c ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, sum_rotated[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_8_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, sum_rotated01[8]}), .a ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, sum_rotated23[8]}), .c ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, sum_rotated[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_9_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, sum_rotated01[9]}), .a ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, sum_rotated23[9]}), .c ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, sum_rotated[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_10_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, sum_rotated01[10]}), .a ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, sum_rotated23[10]}), .c ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, sum_rotated[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_11_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, sum_rotated01[11]}), .a ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, sum_rotated23[11]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, sum_rotated[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_12_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, sum_rotated01[12]}), .a ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, sum_rotated23[12]}), .c ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, sum_rotated[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_13_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, sum_rotated01[13]}), .a ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, sum_rotated23[13]}), .c ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, sum_rotated[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_14_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, sum_rotated01[14]}), .a ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, sum_rotated23[14]}), .c ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, sum_rotated[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_15_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, sum_rotated01[15]}), .a ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, sum_rotated23[15]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, sum_rotated[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_17_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, sum_rotated01[17]}), .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, sum_rotated23[17]}), .c ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, sum_rotated[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_18_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, sum_rotated01[18]}), .a ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, sum_rotated23[18]}), .c ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, sum_rotated[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_19_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, sum_rotated01[19]}), .a ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, sum_rotated23[19]}), .c ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, sum_rotated[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_20_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, sum_rotated01[20]}), .a ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, sum_rotated23[20]}), .c ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, sum_rotated[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_21_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, sum_rotated01[21]}), .a ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, sum_rotated23[21]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, sum_rotated[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_22_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, sum_rotated01[22]}), .a ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, sum_rotated23[22]}), .c ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, sum_rotated[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_23_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, sum_rotated01[23]}), .a ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, sum_rotated23[23]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, sum_rotated[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_24_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, sum_rotated01[24]}), .a ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, sum_rotated23[24]}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, sum_rotated[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_25_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, sum_rotated01[25]}), .a ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, sum_rotated23[25]}), .c ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, sum_rotated[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_26_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, sum_rotated01[26]}), .a ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, sum_rotated23[26]}), .c ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, sum_rotated[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_27_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, sum_rotated01[27]}), .a ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, sum_rotated23[27]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, sum_rotated[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_28_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, sum_rotated01[28]}), .a ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, sum_rotated23[28]}), .c ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, sum_rotated[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_29_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, sum_rotated01[29]}), .a ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, sum_rotated23[29]}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, sum_rotated[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_30_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, sum_rotated01[30]}), .a ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, sum_rotated23[30]}), .c ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, sum_rotated[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) M6_mux_inst_31_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, sum_rotated01[31]}), .a ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, sum_rotated23[31]}), .c ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, sum_rotated[31]}) ) ;

endmodule
