/* modified netlist. Source: module elephant_perm in file ./test/elephant_perm.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module elephant_perm_HPC2_ClockGating_d1 (input0_s0, lfsr, rev_lfsr, clk, input0_s1, Fresh, /*rst,*/ output0_s0, output0_s1/*, Synch*/);
    input [159:0] input0_s0 ;
    input [6:0] lfsr ;
    input [6:0] rev_lfsr ;
    input clk ;
    input [159:0] input0_s1 ;
    //input rst ;
    input [279:0] Fresh ;
    output [159:0] output0_s0 ;
    output [159:0] output0_s1 ;
    //output Synch ;
    wire input_array_6 ;
    wire input_array_5 ;
    wire input_array_4 ;
    wire input_array_3 ;
    wire input_array_2 ;
    wire input_array_1 ;
    wire input_array_0 ;
    wire sbox_inst_39_n20 ;
    wire sbox_inst_39_n19 ;
    wire sbox_inst_39_n18 ;
    wire sbox_inst_39_n17 ;
    wire sbox_inst_39_n16 ;
    wire sbox_inst_39_n15 ;
    wire sbox_inst_39_n14 ;
    wire sbox_inst_39_n13 ;
    wire sbox_inst_39_n12 ;
    wire sbox_inst_39_n11 ;
    wire sbox_inst_39_T6 ;
    wire sbox_inst_39_L0 ;
    wire sbox_inst_39_T5 ;
    wire sbox_inst_39_T4 ;
    wire sbox_inst_39_T3 ;
    wire sbox_inst_39_T2 ;
    wire sbox_inst_39_T1 ;
    wire sbox_inst_39_T0 ;
    wire sbox_inst_38_n20 ;
    wire sbox_inst_38_n19 ;
    wire sbox_inst_38_n18 ;
    wire sbox_inst_38_n17 ;
    wire sbox_inst_38_n16 ;
    wire sbox_inst_38_n15 ;
    wire sbox_inst_38_n14 ;
    wire sbox_inst_38_n13 ;
    wire sbox_inst_38_n12 ;
    wire sbox_inst_38_n11 ;
    wire sbox_inst_38_T6 ;
    wire sbox_inst_38_L0 ;
    wire sbox_inst_38_T5 ;
    wire sbox_inst_38_T4 ;
    wire sbox_inst_38_T3 ;
    wire sbox_inst_38_T2 ;
    wire sbox_inst_38_T1 ;
    wire sbox_inst_38_T0 ;
    wire sbox_inst_37_n20 ;
    wire sbox_inst_37_n19 ;
    wire sbox_inst_37_n18 ;
    wire sbox_inst_37_n17 ;
    wire sbox_inst_37_n16 ;
    wire sbox_inst_37_n15 ;
    wire sbox_inst_37_n14 ;
    wire sbox_inst_37_n13 ;
    wire sbox_inst_37_n12 ;
    wire sbox_inst_37_n11 ;
    wire sbox_inst_37_T6 ;
    wire sbox_inst_37_L0 ;
    wire sbox_inst_37_T5 ;
    wire sbox_inst_37_T4 ;
    wire sbox_inst_37_T3 ;
    wire sbox_inst_37_T2 ;
    wire sbox_inst_37_T1 ;
    wire sbox_inst_37_T0 ;
    wire sbox_inst_36_n20 ;
    wire sbox_inst_36_n19 ;
    wire sbox_inst_36_n18 ;
    wire sbox_inst_36_n17 ;
    wire sbox_inst_36_n16 ;
    wire sbox_inst_36_n15 ;
    wire sbox_inst_36_n14 ;
    wire sbox_inst_36_n13 ;
    wire sbox_inst_36_n12 ;
    wire sbox_inst_36_n11 ;
    wire sbox_inst_36_T6 ;
    wire sbox_inst_36_L0 ;
    wire sbox_inst_36_T5 ;
    wire sbox_inst_36_T4 ;
    wire sbox_inst_36_T3 ;
    wire sbox_inst_36_T2 ;
    wire sbox_inst_36_T1 ;
    wire sbox_inst_36_T0 ;
    wire sbox_inst_35_n20 ;
    wire sbox_inst_35_n19 ;
    wire sbox_inst_35_n18 ;
    wire sbox_inst_35_n17 ;
    wire sbox_inst_35_n16 ;
    wire sbox_inst_35_n15 ;
    wire sbox_inst_35_n14 ;
    wire sbox_inst_35_n13 ;
    wire sbox_inst_35_n12 ;
    wire sbox_inst_35_n11 ;
    wire sbox_inst_35_T6 ;
    wire sbox_inst_35_L0 ;
    wire sbox_inst_35_T5 ;
    wire sbox_inst_35_T4 ;
    wire sbox_inst_35_T3 ;
    wire sbox_inst_35_T2 ;
    wire sbox_inst_35_T1 ;
    wire sbox_inst_35_T0 ;
    wire sbox_inst_34_n20 ;
    wire sbox_inst_34_n19 ;
    wire sbox_inst_34_n18 ;
    wire sbox_inst_34_n17 ;
    wire sbox_inst_34_n16 ;
    wire sbox_inst_34_n15 ;
    wire sbox_inst_34_n14 ;
    wire sbox_inst_34_n13 ;
    wire sbox_inst_34_n12 ;
    wire sbox_inst_34_n11 ;
    wire sbox_inst_34_T6 ;
    wire sbox_inst_34_L0 ;
    wire sbox_inst_34_T5 ;
    wire sbox_inst_34_T4 ;
    wire sbox_inst_34_T3 ;
    wire sbox_inst_34_T2 ;
    wire sbox_inst_34_T1 ;
    wire sbox_inst_34_T0 ;
    wire sbox_inst_33_n20 ;
    wire sbox_inst_33_n19 ;
    wire sbox_inst_33_n18 ;
    wire sbox_inst_33_n17 ;
    wire sbox_inst_33_n16 ;
    wire sbox_inst_33_n15 ;
    wire sbox_inst_33_n14 ;
    wire sbox_inst_33_n13 ;
    wire sbox_inst_33_n12 ;
    wire sbox_inst_33_n11 ;
    wire sbox_inst_33_T6 ;
    wire sbox_inst_33_L0 ;
    wire sbox_inst_33_T5 ;
    wire sbox_inst_33_T4 ;
    wire sbox_inst_33_T3 ;
    wire sbox_inst_33_T2 ;
    wire sbox_inst_33_T1 ;
    wire sbox_inst_33_T0 ;
    wire sbox_inst_32_n20 ;
    wire sbox_inst_32_n19 ;
    wire sbox_inst_32_n18 ;
    wire sbox_inst_32_n17 ;
    wire sbox_inst_32_n16 ;
    wire sbox_inst_32_n15 ;
    wire sbox_inst_32_n14 ;
    wire sbox_inst_32_n13 ;
    wire sbox_inst_32_n12 ;
    wire sbox_inst_32_n11 ;
    wire sbox_inst_32_T6 ;
    wire sbox_inst_32_L0 ;
    wire sbox_inst_32_T5 ;
    wire sbox_inst_32_T4 ;
    wire sbox_inst_32_T3 ;
    wire sbox_inst_32_T2 ;
    wire sbox_inst_32_T1 ;
    wire sbox_inst_32_T0 ;
    wire sbox_inst_31_n20 ;
    wire sbox_inst_31_n19 ;
    wire sbox_inst_31_n18 ;
    wire sbox_inst_31_n17 ;
    wire sbox_inst_31_n16 ;
    wire sbox_inst_31_n15 ;
    wire sbox_inst_31_n14 ;
    wire sbox_inst_31_n13 ;
    wire sbox_inst_31_n12 ;
    wire sbox_inst_31_n11 ;
    wire sbox_inst_31_T6 ;
    wire sbox_inst_31_L0 ;
    wire sbox_inst_31_T5 ;
    wire sbox_inst_31_T4 ;
    wire sbox_inst_31_T3 ;
    wire sbox_inst_31_T2 ;
    wire sbox_inst_31_T1 ;
    wire sbox_inst_31_T0 ;
    wire sbox_inst_30_n20 ;
    wire sbox_inst_30_n19 ;
    wire sbox_inst_30_n18 ;
    wire sbox_inst_30_n17 ;
    wire sbox_inst_30_n16 ;
    wire sbox_inst_30_n15 ;
    wire sbox_inst_30_n14 ;
    wire sbox_inst_30_n13 ;
    wire sbox_inst_30_n12 ;
    wire sbox_inst_30_n11 ;
    wire sbox_inst_30_T6 ;
    wire sbox_inst_30_L0 ;
    wire sbox_inst_30_T5 ;
    wire sbox_inst_30_T4 ;
    wire sbox_inst_30_T3 ;
    wire sbox_inst_30_T2 ;
    wire sbox_inst_30_T1 ;
    wire sbox_inst_30_T0 ;
    wire sbox_inst_29_n20 ;
    wire sbox_inst_29_n19 ;
    wire sbox_inst_29_n18 ;
    wire sbox_inst_29_n17 ;
    wire sbox_inst_29_n16 ;
    wire sbox_inst_29_n15 ;
    wire sbox_inst_29_n14 ;
    wire sbox_inst_29_n13 ;
    wire sbox_inst_29_n12 ;
    wire sbox_inst_29_n11 ;
    wire sbox_inst_29_T6 ;
    wire sbox_inst_29_L0 ;
    wire sbox_inst_29_T5 ;
    wire sbox_inst_29_T4 ;
    wire sbox_inst_29_T3 ;
    wire sbox_inst_29_T2 ;
    wire sbox_inst_29_T1 ;
    wire sbox_inst_29_T0 ;
    wire sbox_inst_28_n20 ;
    wire sbox_inst_28_n19 ;
    wire sbox_inst_28_n18 ;
    wire sbox_inst_28_n17 ;
    wire sbox_inst_28_n16 ;
    wire sbox_inst_28_n15 ;
    wire sbox_inst_28_n14 ;
    wire sbox_inst_28_n13 ;
    wire sbox_inst_28_n12 ;
    wire sbox_inst_28_n11 ;
    wire sbox_inst_28_T6 ;
    wire sbox_inst_28_L0 ;
    wire sbox_inst_28_T5 ;
    wire sbox_inst_28_T4 ;
    wire sbox_inst_28_T3 ;
    wire sbox_inst_28_T2 ;
    wire sbox_inst_28_T1 ;
    wire sbox_inst_28_T0 ;
    wire sbox_inst_27_n20 ;
    wire sbox_inst_27_n19 ;
    wire sbox_inst_27_n18 ;
    wire sbox_inst_27_n17 ;
    wire sbox_inst_27_n16 ;
    wire sbox_inst_27_n15 ;
    wire sbox_inst_27_n14 ;
    wire sbox_inst_27_n13 ;
    wire sbox_inst_27_n12 ;
    wire sbox_inst_27_n11 ;
    wire sbox_inst_27_T6 ;
    wire sbox_inst_27_L0 ;
    wire sbox_inst_27_T5 ;
    wire sbox_inst_27_T4 ;
    wire sbox_inst_27_T3 ;
    wire sbox_inst_27_T2 ;
    wire sbox_inst_27_T1 ;
    wire sbox_inst_27_T0 ;
    wire sbox_inst_26_n20 ;
    wire sbox_inst_26_n19 ;
    wire sbox_inst_26_n18 ;
    wire sbox_inst_26_n17 ;
    wire sbox_inst_26_n16 ;
    wire sbox_inst_26_n15 ;
    wire sbox_inst_26_n14 ;
    wire sbox_inst_26_n13 ;
    wire sbox_inst_26_n12 ;
    wire sbox_inst_26_n11 ;
    wire sbox_inst_26_T6 ;
    wire sbox_inst_26_L0 ;
    wire sbox_inst_26_T5 ;
    wire sbox_inst_26_T4 ;
    wire sbox_inst_26_T3 ;
    wire sbox_inst_26_T2 ;
    wire sbox_inst_26_T1 ;
    wire sbox_inst_26_T0 ;
    wire sbox_inst_25_n20 ;
    wire sbox_inst_25_n19 ;
    wire sbox_inst_25_n18 ;
    wire sbox_inst_25_n17 ;
    wire sbox_inst_25_n16 ;
    wire sbox_inst_25_n15 ;
    wire sbox_inst_25_n14 ;
    wire sbox_inst_25_n13 ;
    wire sbox_inst_25_n12 ;
    wire sbox_inst_25_n11 ;
    wire sbox_inst_25_T6 ;
    wire sbox_inst_25_L0 ;
    wire sbox_inst_25_T5 ;
    wire sbox_inst_25_T4 ;
    wire sbox_inst_25_T3 ;
    wire sbox_inst_25_T2 ;
    wire sbox_inst_25_T1 ;
    wire sbox_inst_25_T0 ;
    wire sbox_inst_24_n20 ;
    wire sbox_inst_24_n19 ;
    wire sbox_inst_24_n18 ;
    wire sbox_inst_24_n17 ;
    wire sbox_inst_24_n16 ;
    wire sbox_inst_24_n15 ;
    wire sbox_inst_24_n14 ;
    wire sbox_inst_24_n13 ;
    wire sbox_inst_24_n12 ;
    wire sbox_inst_24_n11 ;
    wire sbox_inst_24_T6 ;
    wire sbox_inst_24_L0 ;
    wire sbox_inst_24_T5 ;
    wire sbox_inst_24_T4 ;
    wire sbox_inst_24_T3 ;
    wire sbox_inst_24_T2 ;
    wire sbox_inst_24_T1 ;
    wire sbox_inst_24_T0 ;
    wire sbox_inst_23_n20 ;
    wire sbox_inst_23_n19 ;
    wire sbox_inst_23_n18 ;
    wire sbox_inst_23_n17 ;
    wire sbox_inst_23_n16 ;
    wire sbox_inst_23_n15 ;
    wire sbox_inst_23_n14 ;
    wire sbox_inst_23_n13 ;
    wire sbox_inst_23_n12 ;
    wire sbox_inst_23_n11 ;
    wire sbox_inst_23_T6 ;
    wire sbox_inst_23_L0 ;
    wire sbox_inst_23_T5 ;
    wire sbox_inst_23_T4 ;
    wire sbox_inst_23_T3 ;
    wire sbox_inst_23_T2 ;
    wire sbox_inst_23_T1 ;
    wire sbox_inst_23_T0 ;
    wire sbox_inst_22_n20 ;
    wire sbox_inst_22_n19 ;
    wire sbox_inst_22_n18 ;
    wire sbox_inst_22_n17 ;
    wire sbox_inst_22_n16 ;
    wire sbox_inst_22_n15 ;
    wire sbox_inst_22_n14 ;
    wire sbox_inst_22_n13 ;
    wire sbox_inst_22_n12 ;
    wire sbox_inst_22_n11 ;
    wire sbox_inst_22_T6 ;
    wire sbox_inst_22_L0 ;
    wire sbox_inst_22_T5 ;
    wire sbox_inst_22_T4 ;
    wire sbox_inst_22_T3 ;
    wire sbox_inst_22_T2 ;
    wire sbox_inst_22_T1 ;
    wire sbox_inst_22_T0 ;
    wire sbox_inst_21_n20 ;
    wire sbox_inst_21_n19 ;
    wire sbox_inst_21_n18 ;
    wire sbox_inst_21_n17 ;
    wire sbox_inst_21_n16 ;
    wire sbox_inst_21_n15 ;
    wire sbox_inst_21_n14 ;
    wire sbox_inst_21_n13 ;
    wire sbox_inst_21_n12 ;
    wire sbox_inst_21_n11 ;
    wire sbox_inst_21_T6 ;
    wire sbox_inst_21_L0 ;
    wire sbox_inst_21_T5 ;
    wire sbox_inst_21_T4 ;
    wire sbox_inst_21_T3 ;
    wire sbox_inst_21_T2 ;
    wire sbox_inst_21_T1 ;
    wire sbox_inst_21_T0 ;
    wire sbox_inst_20_n20 ;
    wire sbox_inst_20_n19 ;
    wire sbox_inst_20_n18 ;
    wire sbox_inst_20_n17 ;
    wire sbox_inst_20_n16 ;
    wire sbox_inst_20_n15 ;
    wire sbox_inst_20_n14 ;
    wire sbox_inst_20_n13 ;
    wire sbox_inst_20_n12 ;
    wire sbox_inst_20_n11 ;
    wire sbox_inst_20_T6 ;
    wire sbox_inst_20_L0 ;
    wire sbox_inst_20_T5 ;
    wire sbox_inst_20_T4 ;
    wire sbox_inst_20_T3 ;
    wire sbox_inst_20_T2 ;
    wire sbox_inst_20_T1 ;
    wire sbox_inst_20_T0 ;
    wire sbox_inst_19_n20 ;
    wire sbox_inst_19_n19 ;
    wire sbox_inst_19_n18 ;
    wire sbox_inst_19_n17 ;
    wire sbox_inst_19_n16 ;
    wire sbox_inst_19_n15 ;
    wire sbox_inst_19_n14 ;
    wire sbox_inst_19_n13 ;
    wire sbox_inst_19_n12 ;
    wire sbox_inst_19_n11 ;
    wire sbox_inst_19_T6 ;
    wire sbox_inst_19_L0 ;
    wire sbox_inst_19_T5 ;
    wire sbox_inst_19_T4 ;
    wire sbox_inst_19_T3 ;
    wire sbox_inst_19_T2 ;
    wire sbox_inst_19_T1 ;
    wire sbox_inst_19_T0 ;
    wire sbox_inst_18_n20 ;
    wire sbox_inst_18_n19 ;
    wire sbox_inst_18_n18 ;
    wire sbox_inst_18_n17 ;
    wire sbox_inst_18_n16 ;
    wire sbox_inst_18_n15 ;
    wire sbox_inst_18_n14 ;
    wire sbox_inst_18_n13 ;
    wire sbox_inst_18_n12 ;
    wire sbox_inst_18_n11 ;
    wire sbox_inst_18_T6 ;
    wire sbox_inst_18_L0 ;
    wire sbox_inst_18_T5 ;
    wire sbox_inst_18_T4 ;
    wire sbox_inst_18_T3 ;
    wire sbox_inst_18_T2 ;
    wire sbox_inst_18_T1 ;
    wire sbox_inst_18_T0 ;
    wire sbox_inst_17_n20 ;
    wire sbox_inst_17_n19 ;
    wire sbox_inst_17_n18 ;
    wire sbox_inst_17_n17 ;
    wire sbox_inst_17_n16 ;
    wire sbox_inst_17_n15 ;
    wire sbox_inst_17_n14 ;
    wire sbox_inst_17_n13 ;
    wire sbox_inst_17_n12 ;
    wire sbox_inst_17_n11 ;
    wire sbox_inst_17_T6 ;
    wire sbox_inst_17_L0 ;
    wire sbox_inst_17_T5 ;
    wire sbox_inst_17_T4 ;
    wire sbox_inst_17_T3 ;
    wire sbox_inst_17_T2 ;
    wire sbox_inst_17_T1 ;
    wire sbox_inst_17_T0 ;
    wire sbox_inst_16_n20 ;
    wire sbox_inst_16_n19 ;
    wire sbox_inst_16_n18 ;
    wire sbox_inst_16_n17 ;
    wire sbox_inst_16_n16 ;
    wire sbox_inst_16_n15 ;
    wire sbox_inst_16_n14 ;
    wire sbox_inst_16_n13 ;
    wire sbox_inst_16_n12 ;
    wire sbox_inst_16_n11 ;
    wire sbox_inst_16_T6 ;
    wire sbox_inst_16_L0 ;
    wire sbox_inst_16_T5 ;
    wire sbox_inst_16_T4 ;
    wire sbox_inst_16_T3 ;
    wire sbox_inst_16_T2 ;
    wire sbox_inst_16_T1 ;
    wire sbox_inst_16_T0 ;
    wire sbox_inst_15_n20 ;
    wire sbox_inst_15_n19 ;
    wire sbox_inst_15_n18 ;
    wire sbox_inst_15_n17 ;
    wire sbox_inst_15_n16 ;
    wire sbox_inst_15_n15 ;
    wire sbox_inst_15_n14 ;
    wire sbox_inst_15_n13 ;
    wire sbox_inst_15_n12 ;
    wire sbox_inst_15_n11 ;
    wire sbox_inst_15_T6 ;
    wire sbox_inst_15_L0 ;
    wire sbox_inst_15_T5 ;
    wire sbox_inst_15_T4 ;
    wire sbox_inst_15_T3 ;
    wire sbox_inst_15_T2 ;
    wire sbox_inst_15_T1 ;
    wire sbox_inst_15_T0 ;
    wire sbox_inst_14_n20 ;
    wire sbox_inst_14_n19 ;
    wire sbox_inst_14_n18 ;
    wire sbox_inst_14_n17 ;
    wire sbox_inst_14_n16 ;
    wire sbox_inst_14_n15 ;
    wire sbox_inst_14_n14 ;
    wire sbox_inst_14_n13 ;
    wire sbox_inst_14_n12 ;
    wire sbox_inst_14_n11 ;
    wire sbox_inst_14_T6 ;
    wire sbox_inst_14_L0 ;
    wire sbox_inst_14_T5 ;
    wire sbox_inst_14_T4 ;
    wire sbox_inst_14_T3 ;
    wire sbox_inst_14_T2 ;
    wire sbox_inst_14_T1 ;
    wire sbox_inst_14_T0 ;
    wire sbox_inst_13_n20 ;
    wire sbox_inst_13_n19 ;
    wire sbox_inst_13_n18 ;
    wire sbox_inst_13_n17 ;
    wire sbox_inst_13_n16 ;
    wire sbox_inst_13_n15 ;
    wire sbox_inst_13_n14 ;
    wire sbox_inst_13_n13 ;
    wire sbox_inst_13_n12 ;
    wire sbox_inst_13_n11 ;
    wire sbox_inst_13_T6 ;
    wire sbox_inst_13_L0 ;
    wire sbox_inst_13_T5 ;
    wire sbox_inst_13_T4 ;
    wire sbox_inst_13_T3 ;
    wire sbox_inst_13_T2 ;
    wire sbox_inst_13_T1 ;
    wire sbox_inst_13_T0 ;
    wire sbox_inst_12_n20 ;
    wire sbox_inst_12_n19 ;
    wire sbox_inst_12_n18 ;
    wire sbox_inst_12_n17 ;
    wire sbox_inst_12_n16 ;
    wire sbox_inst_12_n15 ;
    wire sbox_inst_12_n14 ;
    wire sbox_inst_12_n13 ;
    wire sbox_inst_12_n12 ;
    wire sbox_inst_12_n11 ;
    wire sbox_inst_12_T6 ;
    wire sbox_inst_12_L0 ;
    wire sbox_inst_12_T5 ;
    wire sbox_inst_12_T4 ;
    wire sbox_inst_12_T3 ;
    wire sbox_inst_12_T2 ;
    wire sbox_inst_12_T1 ;
    wire sbox_inst_12_T0 ;
    wire sbox_inst_11_n20 ;
    wire sbox_inst_11_n19 ;
    wire sbox_inst_11_n18 ;
    wire sbox_inst_11_n17 ;
    wire sbox_inst_11_n16 ;
    wire sbox_inst_11_n15 ;
    wire sbox_inst_11_n14 ;
    wire sbox_inst_11_n13 ;
    wire sbox_inst_11_n12 ;
    wire sbox_inst_11_n11 ;
    wire sbox_inst_11_T6 ;
    wire sbox_inst_11_L0 ;
    wire sbox_inst_11_T5 ;
    wire sbox_inst_11_T4 ;
    wire sbox_inst_11_T3 ;
    wire sbox_inst_11_T2 ;
    wire sbox_inst_11_T1 ;
    wire sbox_inst_11_T0 ;
    wire sbox_inst_10_n20 ;
    wire sbox_inst_10_n19 ;
    wire sbox_inst_10_n18 ;
    wire sbox_inst_10_n17 ;
    wire sbox_inst_10_n16 ;
    wire sbox_inst_10_n15 ;
    wire sbox_inst_10_n14 ;
    wire sbox_inst_10_n13 ;
    wire sbox_inst_10_n12 ;
    wire sbox_inst_10_n11 ;
    wire sbox_inst_10_T6 ;
    wire sbox_inst_10_L0 ;
    wire sbox_inst_10_T5 ;
    wire sbox_inst_10_T4 ;
    wire sbox_inst_10_T3 ;
    wire sbox_inst_10_T2 ;
    wire sbox_inst_10_T1 ;
    wire sbox_inst_10_T0 ;
    wire sbox_inst_9_n20 ;
    wire sbox_inst_9_n19 ;
    wire sbox_inst_9_n18 ;
    wire sbox_inst_9_n17 ;
    wire sbox_inst_9_n16 ;
    wire sbox_inst_9_n15 ;
    wire sbox_inst_9_n14 ;
    wire sbox_inst_9_n13 ;
    wire sbox_inst_9_n12 ;
    wire sbox_inst_9_n11 ;
    wire sbox_inst_9_T6 ;
    wire sbox_inst_9_L0 ;
    wire sbox_inst_9_T5 ;
    wire sbox_inst_9_T4 ;
    wire sbox_inst_9_T3 ;
    wire sbox_inst_9_T2 ;
    wire sbox_inst_9_T1 ;
    wire sbox_inst_9_T0 ;
    wire sbox_inst_8_n20 ;
    wire sbox_inst_8_n19 ;
    wire sbox_inst_8_n18 ;
    wire sbox_inst_8_n17 ;
    wire sbox_inst_8_n16 ;
    wire sbox_inst_8_n15 ;
    wire sbox_inst_8_n14 ;
    wire sbox_inst_8_n13 ;
    wire sbox_inst_8_n12 ;
    wire sbox_inst_8_n11 ;
    wire sbox_inst_8_T6 ;
    wire sbox_inst_8_L0 ;
    wire sbox_inst_8_T5 ;
    wire sbox_inst_8_T4 ;
    wire sbox_inst_8_T3 ;
    wire sbox_inst_8_T2 ;
    wire sbox_inst_8_T1 ;
    wire sbox_inst_8_T0 ;
    wire sbox_inst_7_n20 ;
    wire sbox_inst_7_n19 ;
    wire sbox_inst_7_n18 ;
    wire sbox_inst_7_n17 ;
    wire sbox_inst_7_n16 ;
    wire sbox_inst_7_n15 ;
    wire sbox_inst_7_n14 ;
    wire sbox_inst_7_n13 ;
    wire sbox_inst_7_n12 ;
    wire sbox_inst_7_n11 ;
    wire sbox_inst_7_T6 ;
    wire sbox_inst_7_L0 ;
    wire sbox_inst_7_T5 ;
    wire sbox_inst_7_T4 ;
    wire sbox_inst_7_T3 ;
    wire sbox_inst_7_T2 ;
    wire sbox_inst_7_T1 ;
    wire sbox_inst_7_T0 ;
    wire sbox_inst_6_n20 ;
    wire sbox_inst_6_n19 ;
    wire sbox_inst_6_n18 ;
    wire sbox_inst_6_n17 ;
    wire sbox_inst_6_n16 ;
    wire sbox_inst_6_n15 ;
    wire sbox_inst_6_n14 ;
    wire sbox_inst_6_n13 ;
    wire sbox_inst_6_n12 ;
    wire sbox_inst_6_n11 ;
    wire sbox_inst_6_T6 ;
    wire sbox_inst_6_L0 ;
    wire sbox_inst_6_T5 ;
    wire sbox_inst_6_T4 ;
    wire sbox_inst_6_T3 ;
    wire sbox_inst_6_T2 ;
    wire sbox_inst_6_T1 ;
    wire sbox_inst_6_T0 ;
    wire sbox_inst_5_n20 ;
    wire sbox_inst_5_n19 ;
    wire sbox_inst_5_n18 ;
    wire sbox_inst_5_n17 ;
    wire sbox_inst_5_n16 ;
    wire sbox_inst_5_n15 ;
    wire sbox_inst_5_n14 ;
    wire sbox_inst_5_n13 ;
    wire sbox_inst_5_n12 ;
    wire sbox_inst_5_n11 ;
    wire sbox_inst_5_T6 ;
    wire sbox_inst_5_L0 ;
    wire sbox_inst_5_T5 ;
    wire sbox_inst_5_T4 ;
    wire sbox_inst_5_T3 ;
    wire sbox_inst_5_T2 ;
    wire sbox_inst_5_T1 ;
    wire sbox_inst_5_T0 ;
    wire sbox_inst_4_n20 ;
    wire sbox_inst_4_n19 ;
    wire sbox_inst_4_n18 ;
    wire sbox_inst_4_n17 ;
    wire sbox_inst_4_n16 ;
    wire sbox_inst_4_n15 ;
    wire sbox_inst_4_n14 ;
    wire sbox_inst_4_n13 ;
    wire sbox_inst_4_n12 ;
    wire sbox_inst_4_n11 ;
    wire sbox_inst_4_T6 ;
    wire sbox_inst_4_L0 ;
    wire sbox_inst_4_T5 ;
    wire sbox_inst_4_T4 ;
    wire sbox_inst_4_T3 ;
    wire sbox_inst_4_T2 ;
    wire sbox_inst_4_T1 ;
    wire sbox_inst_4_T0 ;
    wire sbox_inst_3_n20 ;
    wire sbox_inst_3_n19 ;
    wire sbox_inst_3_n18 ;
    wire sbox_inst_3_n17 ;
    wire sbox_inst_3_n16 ;
    wire sbox_inst_3_n15 ;
    wire sbox_inst_3_n14 ;
    wire sbox_inst_3_n13 ;
    wire sbox_inst_3_n12 ;
    wire sbox_inst_3_n11 ;
    wire sbox_inst_3_T6 ;
    wire sbox_inst_3_L0 ;
    wire sbox_inst_3_T5 ;
    wire sbox_inst_3_T4 ;
    wire sbox_inst_3_T3 ;
    wire sbox_inst_3_T2 ;
    wire sbox_inst_3_T1 ;
    wire sbox_inst_3_T0 ;
    wire sbox_inst_2_n20 ;
    wire sbox_inst_2_n19 ;
    wire sbox_inst_2_n18 ;
    wire sbox_inst_2_n17 ;
    wire sbox_inst_2_n16 ;
    wire sbox_inst_2_n15 ;
    wire sbox_inst_2_n14 ;
    wire sbox_inst_2_n13 ;
    wire sbox_inst_2_n12 ;
    wire sbox_inst_2_n11 ;
    wire sbox_inst_2_T6 ;
    wire sbox_inst_2_L0 ;
    wire sbox_inst_2_T5 ;
    wire sbox_inst_2_T4 ;
    wire sbox_inst_2_T3 ;
    wire sbox_inst_2_T2 ;
    wire sbox_inst_2_T1 ;
    wire sbox_inst_2_T0 ;
    wire sbox_inst_1_n20 ;
    wire sbox_inst_1_n19 ;
    wire sbox_inst_1_n18 ;
    wire sbox_inst_1_n17 ;
    wire sbox_inst_1_n16 ;
    wire sbox_inst_1_n15 ;
    wire sbox_inst_1_n14 ;
    wire sbox_inst_1_n13 ;
    wire sbox_inst_1_n12 ;
    wire sbox_inst_1_n11 ;
    wire sbox_inst_1_T6 ;
    wire sbox_inst_1_L0 ;
    wire sbox_inst_1_T5 ;
    wire sbox_inst_1_T4 ;
    wire sbox_inst_1_T3 ;
    wire sbox_inst_1_T2 ;
    wire sbox_inst_1_T1 ;
    wire sbox_inst_1_T0 ;
    wire sbox_inst_0_n20 ;
    wire sbox_inst_0_n19 ;
    wire sbox_inst_0_n18 ;
    wire sbox_inst_0_n17 ;
    wire sbox_inst_0_n16 ;
    wire sbox_inst_0_n15 ;
    wire sbox_inst_0_n14 ;
    wire sbox_inst_0_n13 ;
    wire sbox_inst_0_n12 ;
    wire sbox_inst_0_n11 ;
    wire sbox_inst_0_T6 ;
    wire sbox_inst_0_L0 ;
    wire sbox_inst_0_T5 ;
    wire sbox_inst_0_T4 ;
    wire sbox_inst_0_T3 ;
    wire sbox_inst_0_T2 ;
    wire sbox_inst_0_T1 ;
    wire sbox_inst_0_T0 ;
    wire [159:153] input_array ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2119 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) U29 ( .a ({input0_s1[1], input0_s0[1]}), .b ({1'b0, lfsr[1]}), .c ({new_AGEMA_signal_1076, input_array_1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U30 ( .a ({input0_s1[157], input0_s0[157]}), .b ({1'b0, rev_lfsr[4]}), .c ({new_AGEMA_signal_1078, input_array[157]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U31 ( .a ({input0_s1[153], input0_s0[153]}), .b ({1'b0, rev_lfsr[0]}), .c ({new_AGEMA_signal_1080, input_array[153]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U32 ( .a ({input0_s1[5], input0_s0[5]}), .b ({1'b0, lfsr[5]}), .c ({new_AGEMA_signal_1082, input_array_5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U33 ( .a ({input0_s1[6], input0_s0[6]}), .b ({1'b0, lfsr[6]}), .c ({new_AGEMA_signal_1084, input_array_6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U34 ( .a ({input0_s1[4], input0_s0[4]}), .b ({1'b0, lfsr[4]}), .c ({new_AGEMA_signal_1086, input_array_4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U35 ( .a ({input0_s1[3], input0_s0[3]}), .b ({1'b0, lfsr[3]}), .c ({new_AGEMA_signal_1088, input_array_3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U36 ( .a ({input0_s1[2], input0_s0[2]}), .b ({1'b0, lfsr[2]}), .c ({new_AGEMA_signal_1090, input_array_2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U37 ( .a ({input0_s1[0], input0_s0[0]}), .b ({1'b0, lfsr[0]}), .c ({new_AGEMA_signal_1092, input_array_0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U38 ( .a ({input0_s1[159], input0_s0[159]}), .b ({1'b0, rev_lfsr[6]}), .c ({new_AGEMA_signal_1094, input_array[159]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U39 ( .a ({input0_s1[158], input0_s0[158]}), .b ({1'b0, rev_lfsr[5]}), .c ({new_AGEMA_signal_1096, input_array[158]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U40 ( .a ({input0_s1[156], input0_s0[156]}), .b ({1'b0, rev_lfsr[3]}), .c ({new_AGEMA_signal_1098, input_array[156]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U41 ( .a ({input0_s1[155], input0_s0[155]}), .b ({1'b0, rev_lfsr[2]}), .c ({new_AGEMA_signal_1100, input_array[155]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U42 ( .a ({input0_s1[154], input0_s0[154]}), .b ({1'b0, rev_lfsr[1]}), .c ({new_AGEMA_signal_1102, input_array[154]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U1 ( .a ({new_AGEMA_signal_1096, input_array[158]}), .b ({new_AGEMA_signal_1078, input_array[157]}), .c ({new_AGEMA_signal_1463, sbox_inst_39_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U1 ( .a ({new_AGEMA_signal_1102, input_array[154]}), .b ({new_AGEMA_signal_1080, input_array[153]}), .c ({new_AGEMA_signal_1469, sbox_inst_38_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U1 ( .a ({input0_s1[150], input0_s0[150]}), .b ({input0_s1[149], input0_s0[149]}), .c ({new_AGEMA_signal_1105, sbox_inst_37_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U1 ( .a ({input0_s1[146], input0_s0[146]}), .b ({input0_s1[145], input0_s0[145]}), .c ({new_AGEMA_signal_1115, sbox_inst_36_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U1 ( .a ({input0_s1[142], input0_s0[142]}), .b ({input0_s1[141], input0_s0[141]}), .c ({new_AGEMA_signal_1125, sbox_inst_35_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U1 ( .a ({input0_s1[138], input0_s0[138]}), .b ({input0_s1[137], input0_s0[137]}), .c ({new_AGEMA_signal_1135, sbox_inst_34_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U1 ( .a ({input0_s1[134], input0_s0[134]}), .b ({input0_s1[133], input0_s0[133]}), .c ({new_AGEMA_signal_1145, sbox_inst_33_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U1 ( .a ({input0_s1[130], input0_s0[130]}), .b ({input0_s1[129], input0_s0[129]}), .c ({new_AGEMA_signal_1155, sbox_inst_32_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U1 ( .a ({input0_s1[126], input0_s0[126]}), .b ({input0_s1[125], input0_s0[125]}), .c ({new_AGEMA_signal_1165, sbox_inst_31_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U1 ( .a ({input0_s1[122], input0_s0[122]}), .b ({input0_s1[121], input0_s0[121]}), .c ({new_AGEMA_signal_1175, sbox_inst_30_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U1 ( .a ({input0_s1[118], input0_s0[118]}), .b ({input0_s1[117], input0_s0[117]}), .c ({new_AGEMA_signal_1185, sbox_inst_29_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U1 ( .a ({input0_s1[114], input0_s0[114]}), .b ({input0_s1[113], input0_s0[113]}), .c ({new_AGEMA_signal_1195, sbox_inst_28_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U1 ( .a ({input0_s1[110], input0_s0[110]}), .b ({input0_s1[109], input0_s0[109]}), .c ({new_AGEMA_signal_1205, sbox_inst_27_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U1 ( .a ({input0_s1[106], input0_s0[106]}), .b ({input0_s1[105], input0_s0[105]}), .c ({new_AGEMA_signal_1215, sbox_inst_26_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U1 ( .a ({input0_s1[102], input0_s0[102]}), .b ({input0_s1[101], input0_s0[101]}), .c ({new_AGEMA_signal_1225, sbox_inst_25_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U1 ( .a ({input0_s1[98], input0_s0[98]}), .b ({input0_s1[97], input0_s0[97]}), .c ({new_AGEMA_signal_1235, sbox_inst_24_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U1 ( .a ({input0_s1[94], input0_s0[94]}), .b ({input0_s1[93], input0_s0[93]}), .c ({new_AGEMA_signal_1245, sbox_inst_23_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U1 ( .a ({input0_s1[90], input0_s0[90]}), .b ({input0_s1[89], input0_s0[89]}), .c ({new_AGEMA_signal_1255, sbox_inst_22_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U1 ( .a ({input0_s1[86], input0_s0[86]}), .b ({input0_s1[85], input0_s0[85]}), .c ({new_AGEMA_signal_1265, sbox_inst_21_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U1 ( .a ({input0_s1[82], input0_s0[82]}), .b ({input0_s1[81], input0_s0[81]}), .c ({new_AGEMA_signal_1275, sbox_inst_20_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U1 ( .a ({input0_s1[78], input0_s0[78]}), .b ({input0_s1[77], input0_s0[77]}), .c ({new_AGEMA_signal_1285, sbox_inst_19_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U1 ( .a ({input0_s1[74], input0_s0[74]}), .b ({input0_s1[73], input0_s0[73]}), .c ({new_AGEMA_signal_1295, sbox_inst_18_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U1 ( .a ({input0_s1[70], input0_s0[70]}), .b ({input0_s1[69], input0_s0[69]}), .c ({new_AGEMA_signal_1305, sbox_inst_17_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U1 ( .a ({input0_s1[66], input0_s0[66]}), .b ({input0_s1[65], input0_s0[65]}), .c ({new_AGEMA_signal_1315, sbox_inst_16_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U1 ( .a ({input0_s1[62], input0_s0[62]}), .b ({input0_s1[61], input0_s0[61]}), .c ({new_AGEMA_signal_1325, sbox_inst_15_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U1 ( .a ({input0_s1[58], input0_s0[58]}), .b ({input0_s1[57], input0_s0[57]}), .c ({new_AGEMA_signal_1335, sbox_inst_14_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U1 ( .a ({input0_s1[54], input0_s0[54]}), .b ({input0_s1[53], input0_s0[53]}), .c ({new_AGEMA_signal_1345, sbox_inst_13_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U1 ( .a ({input0_s1[50], input0_s0[50]}), .b ({input0_s1[49], input0_s0[49]}), .c ({new_AGEMA_signal_1355, sbox_inst_12_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U1 ( .a ({input0_s1[46], input0_s0[46]}), .b ({input0_s1[45], input0_s0[45]}), .c ({new_AGEMA_signal_1365, sbox_inst_11_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U1 ( .a ({input0_s1[42], input0_s0[42]}), .b ({input0_s1[41], input0_s0[41]}), .c ({new_AGEMA_signal_1375, sbox_inst_10_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U1 ( .a ({input0_s1[38], input0_s0[38]}), .b ({input0_s1[37], input0_s0[37]}), .c ({new_AGEMA_signal_1385, sbox_inst_9_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U1 ( .a ({input0_s1[34], input0_s0[34]}), .b ({input0_s1[33], input0_s0[33]}), .c ({new_AGEMA_signal_1395, sbox_inst_8_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U1 ( .a ({input0_s1[30], input0_s0[30]}), .b ({input0_s1[29], input0_s0[29]}), .c ({new_AGEMA_signal_1405, sbox_inst_7_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U1 ( .a ({input0_s1[26], input0_s0[26]}), .b ({input0_s1[25], input0_s0[25]}), .c ({new_AGEMA_signal_1415, sbox_inst_6_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U1 ( .a ({input0_s1[22], input0_s0[22]}), .b ({input0_s1[21], input0_s0[21]}), .c ({new_AGEMA_signal_1425, sbox_inst_5_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U1 ( .a ({input0_s1[18], input0_s0[18]}), .b ({input0_s1[17], input0_s0[17]}), .c ({new_AGEMA_signal_1435, sbox_inst_4_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U1 ( .a ({input0_s1[14], input0_s0[14]}), .b ({input0_s1[13], input0_s0[13]}), .c ({new_AGEMA_signal_1445, sbox_inst_3_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U1 ( .a ({input0_s1[10], input0_s0[10]}), .b ({input0_s1[9], input0_s0[9]}), .c ({new_AGEMA_signal_1455, sbox_inst_2_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U1 ( .a ({new_AGEMA_signal_1084, input_array_6}), .b ({new_AGEMA_signal_1082, input_array_5}), .c ({new_AGEMA_signal_1656, sbox_inst_1_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U1 ( .a ({new_AGEMA_signal_1090, input_array_2}), .b ({new_AGEMA_signal_1076, input_array_1}), .c ({new_AGEMA_signal_1663, sbox_inst_0_L0}) ) ;
    //ClockGatingController #(4) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U12 ( .a ({new_AGEMA_signal_1467, sbox_inst_39_T3}), .b ({new_AGEMA_signal_1671, sbox_inst_39_n17}), .c ({new_AGEMA_signal_1870, sbox_inst_39_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U6 ( .a ({new_AGEMA_signal_1468, sbox_inst_39_T4}), .b ({new_AGEMA_signal_1466, sbox_inst_39_T2}), .c ({new_AGEMA_signal_1669, sbox_inst_39_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U5 ( .a ({new_AGEMA_signal_1465, sbox_inst_39_T1}), .b ({new_AGEMA_signal_1096, input_array[158]}), .c ({new_AGEMA_signal_1670, sbox_inst_39_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U4 ( .a ({new_AGEMA_signal_1873, sbox_inst_39_n11}), .b ({new_AGEMA_signal_1078, input_array[157]}), .c ({output0_s1[39], output0_s0[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U3 ( .a ({new_AGEMA_signal_1094, input_array[159]}), .b ({new_AGEMA_signal_1671, sbox_inst_39_n17}), .c ({new_AGEMA_signal_1873, sbox_inst_39_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U2 ( .a ({new_AGEMA_signal_1098, input_array[156]}), .b ({new_AGEMA_signal_1464, sbox_inst_39_T0}), .c ({new_AGEMA_signal_1671, sbox_inst_39_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_t0_AND_U1 ( .a ({new_AGEMA_signal_1078, input_array[157]}), .b ({new_AGEMA_signal_1096, input_array[158]}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_1464, sbox_inst_39_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_t1_AND_U1 ( .a ({new_AGEMA_signal_1098, input_array[156]}), .b ({new_AGEMA_signal_1094, input_array[159]}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_1465, sbox_inst_39_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_t2_AND_U1 ( .a ({new_AGEMA_signal_1078, input_array[157]}), .b ({new_AGEMA_signal_1094, input_array[159]}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_1466, sbox_inst_39_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_t3_AND_U1 ( .a ({new_AGEMA_signal_1096, input_array[158]}), .b ({new_AGEMA_signal_1094, input_array[159]}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_1467, sbox_inst_39_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_t4_AND_U1 ( .a ({new_AGEMA_signal_1098, input_array[156]}), .b ({new_AGEMA_signal_1078, input_array[157]}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_1468, sbox_inst_39_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U12 ( .a ({new_AGEMA_signal_1474, sbox_inst_38_T3}), .b ({new_AGEMA_signal_1676, sbox_inst_38_n17}), .c ({new_AGEMA_signal_1875, sbox_inst_38_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U6 ( .a ({new_AGEMA_signal_1475, sbox_inst_38_T4}), .b ({new_AGEMA_signal_1473, sbox_inst_38_T2}), .c ({new_AGEMA_signal_1674, sbox_inst_38_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U5 ( .a ({new_AGEMA_signal_1472, sbox_inst_38_T1}), .b ({new_AGEMA_signal_1102, input_array[154]}), .c ({new_AGEMA_signal_1675, sbox_inst_38_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U4 ( .a ({new_AGEMA_signal_1878, sbox_inst_38_n11}), .b ({new_AGEMA_signal_1080, input_array[153]}), .c ({output0_s1[38], output0_s0[38]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U3 ( .a ({new_AGEMA_signal_1100, input_array[155]}), .b ({new_AGEMA_signal_1676, sbox_inst_38_n17}), .c ({new_AGEMA_signal_1878, sbox_inst_38_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U2 ( .a ({input0_s1[152], input0_s0[152]}), .b ({new_AGEMA_signal_1470, sbox_inst_38_T0}), .c ({new_AGEMA_signal_1676, sbox_inst_38_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_t0_AND_U1 ( .a ({new_AGEMA_signal_1080, input_array[153]}), .b ({new_AGEMA_signal_1102, input_array[154]}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_1470, sbox_inst_38_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_t1_AND_U1 ( .a ({input0_s1[152], input0_s0[152]}), .b ({new_AGEMA_signal_1100, input_array[155]}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_1472, sbox_inst_38_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_t2_AND_U1 ( .a ({new_AGEMA_signal_1080, input_array[153]}), .b ({new_AGEMA_signal_1100, input_array[155]}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_1473, sbox_inst_38_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_t3_AND_U1 ( .a ({new_AGEMA_signal_1102, input_array[154]}), .b ({new_AGEMA_signal_1100, input_array[155]}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_1474, sbox_inst_38_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_t4_AND_U1 ( .a ({input0_s1[152], input0_s0[152]}), .b ({new_AGEMA_signal_1080, input_array[153]}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_1475, sbox_inst_38_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U12 ( .a ({new_AGEMA_signal_1111, sbox_inst_37_T3}), .b ({new_AGEMA_signal_1478, sbox_inst_37_n17}), .c ({new_AGEMA_signal_1680, sbox_inst_37_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U6 ( .a ({new_AGEMA_signal_1112, sbox_inst_37_T4}), .b ({new_AGEMA_signal_1110, sbox_inst_37_T2}), .c ({new_AGEMA_signal_1476, sbox_inst_37_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U5 ( .a ({new_AGEMA_signal_1109, sbox_inst_37_T1}), .b ({input0_s1[150], input0_s0[150]}), .c ({new_AGEMA_signal_1477, sbox_inst_37_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U4 ( .a ({new_AGEMA_signal_1683, sbox_inst_37_n11}), .b ({input0_s1[149], input0_s0[149]}), .c ({output0_s1[37], output0_s0[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U3 ( .a ({input0_s1[151], input0_s0[151]}), .b ({new_AGEMA_signal_1478, sbox_inst_37_n17}), .c ({new_AGEMA_signal_1683, sbox_inst_37_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U2 ( .a ({input0_s1[148], input0_s0[148]}), .b ({new_AGEMA_signal_1106, sbox_inst_37_T0}), .c ({new_AGEMA_signal_1478, sbox_inst_37_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_t0_AND_U1 ( .a ({input0_s1[149], input0_s0[149]}), .b ({input0_s1[150], input0_s0[150]}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_1106, sbox_inst_37_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_t1_AND_U1 ( .a ({input0_s1[148], input0_s0[148]}), .b ({input0_s1[151], input0_s0[151]}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_1109, sbox_inst_37_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_t2_AND_U1 ( .a ({input0_s1[149], input0_s0[149]}), .b ({input0_s1[151], input0_s0[151]}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_1110, sbox_inst_37_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_t3_AND_U1 ( .a ({input0_s1[150], input0_s0[150]}), .b ({input0_s1[151], input0_s0[151]}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_1111, sbox_inst_37_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_t4_AND_U1 ( .a ({input0_s1[148], input0_s0[148]}), .b ({input0_s1[149], input0_s0[149]}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_1112, sbox_inst_37_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U12 ( .a ({new_AGEMA_signal_1121, sbox_inst_36_T3}), .b ({new_AGEMA_signal_1483, sbox_inst_36_n17}), .c ({new_AGEMA_signal_1685, sbox_inst_36_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U6 ( .a ({new_AGEMA_signal_1122, sbox_inst_36_T4}), .b ({new_AGEMA_signal_1120, sbox_inst_36_T2}), .c ({new_AGEMA_signal_1481, sbox_inst_36_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U5 ( .a ({new_AGEMA_signal_1119, sbox_inst_36_T1}), .b ({input0_s1[146], input0_s0[146]}), .c ({new_AGEMA_signal_1482, sbox_inst_36_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U4 ( .a ({new_AGEMA_signal_1688, sbox_inst_36_n11}), .b ({input0_s1[145], input0_s0[145]}), .c ({output0_s1[36], output0_s0[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U3 ( .a ({input0_s1[147], input0_s0[147]}), .b ({new_AGEMA_signal_1483, sbox_inst_36_n17}), .c ({new_AGEMA_signal_1688, sbox_inst_36_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U2 ( .a ({input0_s1[144], input0_s0[144]}), .b ({new_AGEMA_signal_1116, sbox_inst_36_T0}), .c ({new_AGEMA_signal_1483, sbox_inst_36_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_t0_AND_U1 ( .a ({input0_s1[145], input0_s0[145]}), .b ({input0_s1[146], input0_s0[146]}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_1116, sbox_inst_36_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_t1_AND_U1 ( .a ({input0_s1[144], input0_s0[144]}), .b ({input0_s1[147], input0_s0[147]}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_1119, sbox_inst_36_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_t2_AND_U1 ( .a ({input0_s1[145], input0_s0[145]}), .b ({input0_s1[147], input0_s0[147]}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_1120, sbox_inst_36_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_t3_AND_U1 ( .a ({input0_s1[146], input0_s0[146]}), .b ({input0_s1[147], input0_s0[147]}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_1121, sbox_inst_36_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_t4_AND_U1 ( .a ({input0_s1[144], input0_s0[144]}), .b ({input0_s1[145], input0_s0[145]}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_1122, sbox_inst_36_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U12 ( .a ({new_AGEMA_signal_1131, sbox_inst_35_T3}), .b ({new_AGEMA_signal_1488, sbox_inst_35_n17}), .c ({new_AGEMA_signal_1690, sbox_inst_35_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U6 ( .a ({new_AGEMA_signal_1132, sbox_inst_35_T4}), .b ({new_AGEMA_signal_1130, sbox_inst_35_T2}), .c ({new_AGEMA_signal_1486, sbox_inst_35_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U5 ( .a ({new_AGEMA_signal_1129, sbox_inst_35_T1}), .b ({input0_s1[142], input0_s0[142]}), .c ({new_AGEMA_signal_1487, sbox_inst_35_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U4 ( .a ({new_AGEMA_signal_1693, sbox_inst_35_n11}), .b ({input0_s1[141], input0_s0[141]}), .c ({output0_s1[35], output0_s0[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U3 ( .a ({input0_s1[143], input0_s0[143]}), .b ({new_AGEMA_signal_1488, sbox_inst_35_n17}), .c ({new_AGEMA_signal_1693, sbox_inst_35_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U2 ( .a ({input0_s1[140], input0_s0[140]}), .b ({new_AGEMA_signal_1126, sbox_inst_35_T0}), .c ({new_AGEMA_signal_1488, sbox_inst_35_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_t0_AND_U1 ( .a ({input0_s1[141], input0_s0[141]}), .b ({input0_s1[142], input0_s0[142]}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_1126, sbox_inst_35_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_t1_AND_U1 ( .a ({input0_s1[140], input0_s0[140]}), .b ({input0_s1[143], input0_s0[143]}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_1129, sbox_inst_35_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_t2_AND_U1 ( .a ({input0_s1[141], input0_s0[141]}), .b ({input0_s1[143], input0_s0[143]}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_1130, sbox_inst_35_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_t3_AND_U1 ( .a ({input0_s1[142], input0_s0[142]}), .b ({input0_s1[143], input0_s0[143]}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_1131, sbox_inst_35_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_t4_AND_U1 ( .a ({input0_s1[140], input0_s0[140]}), .b ({input0_s1[141], input0_s0[141]}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_1132, sbox_inst_35_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U12 ( .a ({new_AGEMA_signal_1141, sbox_inst_34_T3}), .b ({new_AGEMA_signal_1493, sbox_inst_34_n17}), .c ({new_AGEMA_signal_1695, sbox_inst_34_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U6 ( .a ({new_AGEMA_signal_1142, sbox_inst_34_T4}), .b ({new_AGEMA_signal_1140, sbox_inst_34_T2}), .c ({new_AGEMA_signal_1491, sbox_inst_34_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U5 ( .a ({new_AGEMA_signal_1139, sbox_inst_34_T1}), .b ({input0_s1[138], input0_s0[138]}), .c ({new_AGEMA_signal_1492, sbox_inst_34_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U4 ( .a ({new_AGEMA_signal_1698, sbox_inst_34_n11}), .b ({input0_s1[137], input0_s0[137]}), .c ({output0_s1[34], output0_s0[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U3 ( .a ({input0_s1[139], input0_s0[139]}), .b ({new_AGEMA_signal_1493, sbox_inst_34_n17}), .c ({new_AGEMA_signal_1698, sbox_inst_34_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U2 ( .a ({input0_s1[136], input0_s0[136]}), .b ({new_AGEMA_signal_1136, sbox_inst_34_T0}), .c ({new_AGEMA_signal_1493, sbox_inst_34_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_t0_AND_U1 ( .a ({input0_s1[137], input0_s0[137]}), .b ({input0_s1[138], input0_s0[138]}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_1136, sbox_inst_34_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_t1_AND_U1 ( .a ({input0_s1[136], input0_s0[136]}), .b ({input0_s1[139], input0_s0[139]}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_1139, sbox_inst_34_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_t2_AND_U1 ( .a ({input0_s1[137], input0_s0[137]}), .b ({input0_s1[139], input0_s0[139]}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_1140, sbox_inst_34_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_t3_AND_U1 ( .a ({input0_s1[138], input0_s0[138]}), .b ({input0_s1[139], input0_s0[139]}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_1141, sbox_inst_34_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_t4_AND_U1 ( .a ({input0_s1[136], input0_s0[136]}), .b ({input0_s1[137], input0_s0[137]}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_1142, sbox_inst_34_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U12 ( .a ({new_AGEMA_signal_1151, sbox_inst_33_T3}), .b ({new_AGEMA_signal_1498, sbox_inst_33_n17}), .c ({new_AGEMA_signal_1700, sbox_inst_33_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U6 ( .a ({new_AGEMA_signal_1152, sbox_inst_33_T4}), .b ({new_AGEMA_signal_1150, sbox_inst_33_T2}), .c ({new_AGEMA_signal_1496, sbox_inst_33_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U5 ( .a ({new_AGEMA_signal_1149, sbox_inst_33_T1}), .b ({input0_s1[134], input0_s0[134]}), .c ({new_AGEMA_signal_1497, sbox_inst_33_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U4 ( .a ({new_AGEMA_signal_1703, sbox_inst_33_n11}), .b ({input0_s1[133], input0_s0[133]}), .c ({output0_s1[33], output0_s0[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U3 ( .a ({input0_s1[135], input0_s0[135]}), .b ({new_AGEMA_signal_1498, sbox_inst_33_n17}), .c ({new_AGEMA_signal_1703, sbox_inst_33_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U2 ( .a ({input0_s1[132], input0_s0[132]}), .b ({new_AGEMA_signal_1146, sbox_inst_33_T0}), .c ({new_AGEMA_signal_1498, sbox_inst_33_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_t0_AND_U1 ( .a ({input0_s1[133], input0_s0[133]}), .b ({input0_s1[134], input0_s0[134]}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_1146, sbox_inst_33_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_t1_AND_U1 ( .a ({input0_s1[132], input0_s0[132]}), .b ({input0_s1[135], input0_s0[135]}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_1149, sbox_inst_33_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_t2_AND_U1 ( .a ({input0_s1[133], input0_s0[133]}), .b ({input0_s1[135], input0_s0[135]}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_1150, sbox_inst_33_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_t3_AND_U1 ( .a ({input0_s1[134], input0_s0[134]}), .b ({input0_s1[135], input0_s0[135]}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_1151, sbox_inst_33_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_t4_AND_U1 ( .a ({input0_s1[132], input0_s0[132]}), .b ({input0_s1[133], input0_s0[133]}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_1152, sbox_inst_33_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U12 ( .a ({new_AGEMA_signal_1161, sbox_inst_32_T3}), .b ({new_AGEMA_signal_1503, sbox_inst_32_n17}), .c ({new_AGEMA_signal_1705, sbox_inst_32_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U6 ( .a ({new_AGEMA_signal_1162, sbox_inst_32_T4}), .b ({new_AGEMA_signal_1160, sbox_inst_32_T2}), .c ({new_AGEMA_signal_1501, sbox_inst_32_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U5 ( .a ({new_AGEMA_signal_1159, sbox_inst_32_T1}), .b ({input0_s1[130], input0_s0[130]}), .c ({new_AGEMA_signal_1502, sbox_inst_32_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U4 ( .a ({new_AGEMA_signal_1708, sbox_inst_32_n11}), .b ({input0_s1[129], input0_s0[129]}), .c ({output0_s1[32], output0_s0[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U3 ( .a ({input0_s1[131], input0_s0[131]}), .b ({new_AGEMA_signal_1503, sbox_inst_32_n17}), .c ({new_AGEMA_signal_1708, sbox_inst_32_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U2 ( .a ({input0_s1[128], input0_s0[128]}), .b ({new_AGEMA_signal_1156, sbox_inst_32_T0}), .c ({new_AGEMA_signal_1503, sbox_inst_32_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_t0_AND_U1 ( .a ({input0_s1[129], input0_s0[129]}), .b ({input0_s1[130], input0_s0[130]}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_1156, sbox_inst_32_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_t1_AND_U1 ( .a ({input0_s1[128], input0_s0[128]}), .b ({input0_s1[131], input0_s0[131]}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_1159, sbox_inst_32_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_t2_AND_U1 ( .a ({input0_s1[129], input0_s0[129]}), .b ({input0_s1[131], input0_s0[131]}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_1160, sbox_inst_32_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_t3_AND_U1 ( .a ({input0_s1[130], input0_s0[130]}), .b ({input0_s1[131], input0_s0[131]}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_1161, sbox_inst_32_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_t4_AND_U1 ( .a ({input0_s1[128], input0_s0[128]}), .b ({input0_s1[129], input0_s0[129]}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_1162, sbox_inst_32_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U12 ( .a ({new_AGEMA_signal_1171, sbox_inst_31_T3}), .b ({new_AGEMA_signal_1508, sbox_inst_31_n17}), .c ({new_AGEMA_signal_1710, sbox_inst_31_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U6 ( .a ({new_AGEMA_signal_1172, sbox_inst_31_T4}), .b ({new_AGEMA_signal_1170, sbox_inst_31_T2}), .c ({new_AGEMA_signal_1506, sbox_inst_31_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U5 ( .a ({new_AGEMA_signal_1169, sbox_inst_31_T1}), .b ({input0_s1[126], input0_s0[126]}), .c ({new_AGEMA_signal_1507, sbox_inst_31_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U4 ( .a ({new_AGEMA_signal_1713, sbox_inst_31_n11}), .b ({input0_s1[125], input0_s0[125]}), .c ({output0_s1[31], output0_s0[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U3 ( .a ({input0_s1[127], input0_s0[127]}), .b ({new_AGEMA_signal_1508, sbox_inst_31_n17}), .c ({new_AGEMA_signal_1713, sbox_inst_31_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U2 ( .a ({input0_s1[124], input0_s0[124]}), .b ({new_AGEMA_signal_1166, sbox_inst_31_T0}), .c ({new_AGEMA_signal_1508, sbox_inst_31_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_t0_AND_U1 ( .a ({input0_s1[125], input0_s0[125]}), .b ({input0_s1[126], input0_s0[126]}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_1166, sbox_inst_31_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_t1_AND_U1 ( .a ({input0_s1[124], input0_s0[124]}), .b ({input0_s1[127], input0_s0[127]}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_1169, sbox_inst_31_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_t2_AND_U1 ( .a ({input0_s1[125], input0_s0[125]}), .b ({input0_s1[127], input0_s0[127]}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_1170, sbox_inst_31_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_t3_AND_U1 ( .a ({input0_s1[126], input0_s0[126]}), .b ({input0_s1[127], input0_s0[127]}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_1171, sbox_inst_31_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_t4_AND_U1 ( .a ({input0_s1[124], input0_s0[124]}), .b ({input0_s1[125], input0_s0[125]}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_1172, sbox_inst_31_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U12 ( .a ({new_AGEMA_signal_1181, sbox_inst_30_T3}), .b ({new_AGEMA_signal_1513, sbox_inst_30_n17}), .c ({new_AGEMA_signal_1715, sbox_inst_30_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U6 ( .a ({new_AGEMA_signal_1182, sbox_inst_30_T4}), .b ({new_AGEMA_signal_1180, sbox_inst_30_T2}), .c ({new_AGEMA_signal_1511, sbox_inst_30_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U5 ( .a ({new_AGEMA_signal_1179, sbox_inst_30_T1}), .b ({input0_s1[122], input0_s0[122]}), .c ({new_AGEMA_signal_1512, sbox_inst_30_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U4 ( .a ({new_AGEMA_signal_1718, sbox_inst_30_n11}), .b ({input0_s1[121], input0_s0[121]}), .c ({output0_s1[30], output0_s0[30]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U3 ( .a ({input0_s1[123], input0_s0[123]}), .b ({new_AGEMA_signal_1513, sbox_inst_30_n17}), .c ({new_AGEMA_signal_1718, sbox_inst_30_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U2 ( .a ({input0_s1[120], input0_s0[120]}), .b ({new_AGEMA_signal_1176, sbox_inst_30_T0}), .c ({new_AGEMA_signal_1513, sbox_inst_30_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_t0_AND_U1 ( .a ({input0_s1[121], input0_s0[121]}), .b ({input0_s1[122], input0_s0[122]}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_1176, sbox_inst_30_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_t1_AND_U1 ( .a ({input0_s1[120], input0_s0[120]}), .b ({input0_s1[123], input0_s0[123]}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_1179, sbox_inst_30_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_t2_AND_U1 ( .a ({input0_s1[121], input0_s0[121]}), .b ({input0_s1[123], input0_s0[123]}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_1180, sbox_inst_30_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_t3_AND_U1 ( .a ({input0_s1[122], input0_s0[122]}), .b ({input0_s1[123], input0_s0[123]}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_1181, sbox_inst_30_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_t4_AND_U1 ( .a ({input0_s1[120], input0_s0[120]}), .b ({input0_s1[121], input0_s0[121]}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_1182, sbox_inst_30_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U12 ( .a ({new_AGEMA_signal_1191, sbox_inst_29_T3}), .b ({new_AGEMA_signal_1518, sbox_inst_29_n17}), .c ({new_AGEMA_signal_1720, sbox_inst_29_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U6 ( .a ({new_AGEMA_signal_1192, sbox_inst_29_T4}), .b ({new_AGEMA_signal_1190, sbox_inst_29_T2}), .c ({new_AGEMA_signal_1516, sbox_inst_29_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U5 ( .a ({new_AGEMA_signal_1189, sbox_inst_29_T1}), .b ({input0_s1[118], input0_s0[118]}), .c ({new_AGEMA_signal_1517, sbox_inst_29_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U4 ( .a ({new_AGEMA_signal_1723, sbox_inst_29_n11}), .b ({input0_s1[117], input0_s0[117]}), .c ({output0_s1[29], output0_s0[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U3 ( .a ({input0_s1[119], input0_s0[119]}), .b ({new_AGEMA_signal_1518, sbox_inst_29_n17}), .c ({new_AGEMA_signal_1723, sbox_inst_29_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U2 ( .a ({input0_s1[116], input0_s0[116]}), .b ({new_AGEMA_signal_1186, sbox_inst_29_T0}), .c ({new_AGEMA_signal_1518, sbox_inst_29_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_t0_AND_U1 ( .a ({input0_s1[117], input0_s0[117]}), .b ({input0_s1[118], input0_s0[118]}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_1186, sbox_inst_29_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_t1_AND_U1 ( .a ({input0_s1[116], input0_s0[116]}), .b ({input0_s1[119], input0_s0[119]}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_1189, sbox_inst_29_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_t2_AND_U1 ( .a ({input0_s1[117], input0_s0[117]}), .b ({input0_s1[119], input0_s0[119]}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_1190, sbox_inst_29_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_t3_AND_U1 ( .a ({input0_s1[118], input0_s0[118]}), .b ({input0_s1[119], input0_s0[119]}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_1191, sbox_inst_29_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_t4_AND_U1 ( .a ({input0_s1[116], input0_s0[116]}), .b ({input0_s1[117], input0_s0[117]}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_1192, sbox_inst_29_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U12 ( .a ({new_AGEMA_signal_1201, sbox_inst_28_T3}), .b ({new_AGEMA_signal_1523, sbox_inst_28_n17}), .c ({new_AGEMA_signal_1725, sbox_inst_28_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U6 ( .a ({new_AGEMA_signal_1202, sbox_inst_28_T4}), .b ({new_AGEMA_signal_1200, sbox_inst_28_T2}), .c ({new_AGEMA_signal_1521, sbox_inst_28_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U5 ( .a ({new_AGEMA_signal_1199, sbox_inst_28_T1}), .b ({input0_s1[114], input0_s0[114]}), .c ({new_AGEMA_signal_1522, sbox_inst_28_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U4 ( .a ({new_AGEMA_signal_1728, sbox_inst_28_n11}), .b ({input0_s1[113], input0_s0[113]}), .c ({output0_s1[28], output0_s0[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U3 ( .a ({input0_s1[115], input0_s0[115]}), .b ({new_AGEMA_signal_1523, sbox_inst_28_n17}), .c ({new_AGEMA_signal_1728, sbox_inst_28_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U2 ( .a ({input0_s1[112], input0_s0[112]}), .b ({new_AGEMA_signal_1196, sbox_inst_28_T0}), .c ({new_AGEMA_signal_1523, sbox_inst_28_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_t0_AND_U1 ( .a ({input0_s1[113], input0_s0[113]}), .b ({input0_s1[114], input0_s0[114]}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_1196, sbox_inst_28_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_t1_AND_U1 ( .a ({input0_s1[112], input0_s0[112]}), .b ({input0_s1[115], input0_s0[115]}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_1199, sbox_inst_28_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_t2_AND_U1 ( .a ({input0_s1[113], input0_s0[113]}), .b ({input0_s1[115], input0_s0[115]}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_1200, sbox_inst_28_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_t3_AND_U1 ( .a ({input0_s1[114], input0_s0[114]}), .b ({input0_s1[115], input0_s0[115]}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_1201, sbox_inst_28_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_t4_AND_U1 ( .a ({input0_s1[112], input0_s0[112]}), .b ({input0_s1[113], input0_s0[113]}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_1202, sbox_inst_28_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U12 ( .a ({new_AGEMA_signal_1211, sbox_inst_27_T3}), .b ({new_AGEMA_signal_1528, sbox_inst_27_n17}), .c ({new_AGEMA_signal_1730, sbox_inst_27_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U6 ( .a ({new_AGEMA_signal_1212, sbox_inst_27_T4}), .b ({new_AGEMA_signal_1210, sbox_inst_27_T2}), .c ({new_AGEMA_signal_1526, sbox_inst_27_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U5 ( .a ({new_AGEMA_signal_1209, sbox_inst_27_T1}), .b ({input0_s1[110], input0_s0[110]}), .c ({new_AGEMA_signal_1527, sbox_inst_27_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U4 ( .a ({new_AGEMA_signal_1733, sbox_inst_27_n11}), .b ({input0_s1[109], input0_s0[109]}), .c ({output0_s1[27], output0_s0[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U3 ( .a ({input0_s1[111], input0_s0[111]}), .b ({new_AGEMA_signal_1528, sbox_inst_27_n17}), .c ({new_AGEMA_signal_1733, sbox_inst_27_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U2 ( .a ({input0_s1[108], input0_s0[108]}), .b ({new_AGEMA_signal_1206, sbox_inst_27_T0}), .c ({new_AGEMA_signal_1528, sbox_inst_27_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_t0_AND_U1 ( .a ({input0_s1[109], input0_s0[109]}), .b ({input0_s1[110], input0_s0[110]}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_1206, sbox_inst_27_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_t1_AND_U1 ( .a ({input0_s1[108], input0_s0[108]}), .b ({input0_s1[111], input0_s0[111]}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_1209, sbox_inst_27_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_t2_AND_U1 ( .a ({input0_s1[109], input0_s0[109]}), .b ({input0_s1[111], input0_s0[111]}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_1210, sbox_inst_27_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_t3_AND_U1 ( .a ({input0_s1[110], input0_s0[110]}), .b ({input0_s1[111], input0_s0[111]}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_1211, sbox_inst_27_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_t4_AND_U1 ( .a ({input0_s1[108], input0_s0[108]}), .b ({input0_s1[109], input0_s0[109]}), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_1212, sbox_inst_27_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U12 ( .a ({new_AGEMA_signal_1221, sbox_inst_26_T3}), .b ({new_AGEMA_signal_1533, sbox_inst_26_n17}), .c ({new_AGEMA_signal_1735, sbox_inst_26_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U6 ( .a ({new_AGEMA_signal_1222, sbox_inst_26_T4}), .b ({new_AGEMA_signal_1220, sbox_inst_26_T2}), .c ({new_AGEMA_signal_1531, sbox_inst_26_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U5 ( .a ({new_AGEMA_signal_1219, sbox_inst_26_T1}), .b ({input0_s1[106], input0_s0[106]}), .c ({new_AGEMA_signal_1532, sbox_inst_26_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U4 ( .a ({new_AGEMA_signal_1738, sbox_inst_26_n11}), .b ({input0_s1[105], input0_s0[105]}), .c ({output0_s1[26], output0_s0[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U3 ( .a ({input0_s1[107], input0_s0[107]}), .b ({new_AGEMA_signal_1533, sbox_inst_26_n17}), .c ({new_AGEMA_signal_1738, sbox_inst_26_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U2 ( .a ({input0_s1[104], input0_s0[104]}), .b ({new_AGEMA_signal_1216, sbox_inst_26_T0}), .c ({new_AGEMA_signal_1533, sbox_inst_26_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_t0_AND_U1 ( .a ({input0_s1[105], input0_s0[105]}), .b ({input0_s1[106], input0_s0[106]}), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_1216, sbox_inst_26_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_t1_AND_U1 ( .a ({input0_s1[104], input0_s0[104]}), .b ({input0_s1[107], input0_s0[107]}), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_1219, sbox_inst_26_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_t2_AND_U1 ( .a ({input0_s1[105], input0_s0[105]}), .b ({input0_s1[107], input0_s0[107]}), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_1220, sbox_inst_26_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_t3_AND_U1 ( .a ({input0_s1[106], input0_s0[106]}), .b ({input0_s1[107], input0_s0[107]}), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_1221, sbox_inst_26_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_t4_AND_U1 ( .a ({input0_s1[104], input0_s0[104]}), .b ({input0_s1[105], input0_s0[105]}), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_1222, sbox_inst_26_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U12 ( .a ({new_AGEMA_signal_1231, sbox_inst_25_T3}), .b ({new_AGEMA_signal_1538, sbox_inst_25_n17}), .c ({new_AGEMA_signal_1740, sbox_inst_25_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U6 ( .a ({new_AGEMA_signal_1232, sbox_inst_25_T4}), .b ({new_AGEMA_signal_1230, sbox_inst_25_T2}), .c ({new_AGEMA_signal_1536, sbox_inst_25_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U5 ( .a ({new_AGEMA_signal_1229, sbox_inst_25_T1}), .b ({input0_s1[102], input0_s0[102]}), .c ({new_AGEMA_signal_1537, sbox_inst_25_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U4 ( .a ({new_AGEMA_signal_1743, sbox_inst_25_n11}), .b ({input0_s1[101], input0_s0[101]}), .c ({output0_s1[25], output0_s0[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U3 ( .a ({input0_s1[103], input0_s0[103]}), .b ({new_AGEMA_signal_1538, sbox_inst_25_n17}), .c ({new_AGEMA_signal_1743, sbox_inst_25_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U2 ( .a ({input0_s1[100], input0_s0[100]}), .b ({new_AGEMA_signal_1226, sbox_inst_25_T0}), .c ({new_AGEMA_signal_1538, sbox_inst_25_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_t0_AND_U1 ( .a ({input0_s1[101], input0_s0[101]}), .b ({input0_s1[102], input0_s0[102]}), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_1226, sbox_inst_25_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_t1_AND_U1 ( .a ({input0_s1[100], input0_s0[100]}), .b ({input0_s1[103], input0_s0[103]}), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_1229, sbox_inst_25_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_t2_AND_U1 ( .a ({input0_s1[101], input0_s0[101]}), .b ({input0_s1[103], input0_s0[103]}), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_1230, sbox_inst_25_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_t3_AND_U1 ( .a ({input0_s1[102], input0_s0[102]}), .b ({input0_s1[103], input0_s0[103]}), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_1231, sbox_inst_25_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_t4_AND_U1 ( .a ({input0_s1[100], input0_s0[100]}), .b ({input0_s1[101], input0_s0[101]}), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_1232, sbox_inst_25_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U12 ( .a ({new_AGEMA_signal_1241, sbox_inst_24_T3}), .b ({new_AGEMA_signal_1543, sbox_inst_24_n17}), .c ({new_AGEMA_signal_1745, sbox_inst_24_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U6 ( .a ({new_AGEMA_signal_1242, sbox_inst_24_T4}), .b ({new_AGEMA_signal_1240, sbox_inst_24_T2}), .c ({new_AGEMA_signal_1541, sbox_inst_24_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U5 ( .a ({new_AGEMA_signal_1239, sbox_inst_24_T1}), .b ({input0_s1[98], input0_s0[98]}), .c ({new_AGEMA_signal_1542, sbox_inst_24_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U4 ( .a ({new_AGEMA_signal_1748, sbox_inst_24_n11}), .b ({input0_s1[97], input0_s0[97]}), .c ({output0_s1[24], output0_s0[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U3 ( .a ({input0_s1[99], input0_s0[99]}), .b ({new_AGEMA_signal_1543, sbox_inst_24_n17}), .c ({new_AGEMA_signal_1748, sbox_inst_24_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U2 ( .a ({input0_s1[96], input0_s0[96]}), .b ({new_AGEMA_signal_1236, sbox_inst_24_T0}), .c ({new_AGEMA_signal_1543, sbox_inst_24_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_t0_AND_U1 ( .a ({input0_s1[97], input0_s0[97]}), .b ({input0_s1[98], input0_s0[98]}), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_1236, sbox_inst_24_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_t1_AND_U1 ( .a ({input0_s1[96], input0_s0[96]}), .b ({input0_s1[99], input0_s0[99]}), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_1239, sbox_inst_24_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_t2_AND_U1 ( .a ({input0_s1[97], input0_s0[97]}), .b ({input0_s1[99], input0_s0[99]}), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_1240, sbox_inst_24_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_t3_AND_U1 ( .a ({input0_s1[98], input0_s0[98]}), .b ({input0_s1[99], input0_s0[99]}), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_1241, sbox_inst_24_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_t4_AND_U1 ( .a ({input0_s1[96], input0_s0[96]}), .b ({input0_s1[97], input0_s0[97]}), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_1242, sbox_inst_24_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U12 ( .a ({new_AGEMA_signal_1251, sbox_inst_23_T3}), .b ({new_AGEMA_signal_1548, sbox_inst_23_n17}), .c ({new_AGEMA_signal_1750, sbox_inst_23_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U6 ( .a ({new_AGEMA_signal_1252, sbox_inst_23_T4}), .b ({new_AGEMA_signal_1250, sbox_inst_23_T2}), .c ({new_AGEMA_signal_1546, sbox_inst_23_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U5 ( .a ({new_AGEMA_signal_1249, sbox_inst_23_T1}), .b ({input0_s1[94], input0_s0[94]}), .c ({new_AGEMA_signal_1547, sbox_inst_23_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U4 ( .a ({new_AGEMA_signal_1753, sbox_inst_23_n11}), .b ({input0_s1[93], input0_s0[93]}), .c ({output0_s1[23], output0_s0[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U3 ( .a ({input0_s1[95], input0_s0[95]}), .b ({new_AGEMA_signal_1548, sbox_inst_23_n17}), .c ({new_AGEMA_signal_1753, sbox_inst_23_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U2 ( .a ({input0_s1[92], input0_s0[92]}), .b ({new_AGEMA_signal_1246, sbox_inst_23_T0}), .c ({new_AGEMA_signal_1548, sbox_inst_23_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_t0_AND_U1 ( .a ({input0_s1[93], input0_s0[93]}), .b ({input0_s1[94], input0_s0[94]}), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_1246, sbox_inst_23_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_t1_AND_U1 ( .a ({input0_s1[92], input0_s0[92]}), .b ({input0_s1[95], input0_s0[95]}), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_1249, sbox_inst_23_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_t2_AND_U1 ( .a ({input0_s1[93], input0_s0[93]}), .b ({input0_s1[95], input0_s0[95]}), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_1250, sbox_inst_23_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_t3_AND_U1 ( .a ({input0_s1[94], input0_s0[94]}), .b ({input0_s1[95], input0_s0[95]}), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_1251, sbox_inst_23_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_t4_AND_U1 ( .a ({input0_s1[92], input0_s0[92]}), .b ({input0_s1[93], input0_s0[93]}), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_1252, sbox_inst_23_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U12 ( .a ({new_AGEMA_signal_1261, sbox_inst_22_T3}), .b ({new_AGEMA_signal_1553, sbox_inst_22_n17}), .c ({new_AGEMA_signal_1755, sbox_inst_22_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U6 ( .a ({new_AGEMA_signal_1262, sbox_inst_22_T4}), .b ({new_AGEMA_signal_1260, sbox_inst_22_T2}), .c ({new_AGEMA_signal_1551, sbox_inst_22_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U5 ( .a ({new_AGEMA_signal_1259, sbox_inst_22_T1}), .b ({input0_s1[90], input0_s0[90]}), .c ({new_AGEMA_signal_1552, sbox_inst_22_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U4 ( .a ({new_AGEMA_signal_1758, sbox_inst_22_n11}), .b ({input0_s1[89], input0_s0[89]}), .c ({output0_s1[22], output0_s0[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U3 ( .a ({input0_s1[91], input0_s0[91]}), .b ({new_AGEMA_signal_1553, sbox_inst_22_n17}), .c ({new_AGEMA_signal_1758, sbox_inst_22_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U2 ( .a ({input0_s1[88], input0_s0[88]}), .b ({new_AGEMA_signal_1256, sbox_inst_22_T0}), .c ({new_AGEMA_signal_1553, sbox_inst_22_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_t0_AND_U1 ( .a ({input0_s1[89], input0_s0[89]}), .b ({input0_s1[90], input0_s0[90]}), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_1256, sbox_inst_22_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_t1_AND_U1 ( .a ({input0_s1[88], input0_s0[88]}), .b ({input0_s1[91], input0_s0[91]}), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_1259, sbox_inst_22_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_t2_AND_U1 ( .a ({input0_s1[89], input0_s0[89]}), .b ({input0_s1[91], input0_s0[91]}), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_1260, sbox_inst_22_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_t3_AND_U1 ( .a ({input0_s1[90], input0_s0[90]}), .b ({input0_s1[91], input0_s0[91]}), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_1261, sbox_inst_22_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_t4_AND_U1 ( .a ({input0_s1[88], input0_s0[88]}), .b ({input0_s1[89], input0_s0[89]}), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_1262, sbox_inst_22_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U12 ( .a ({new_AGEMA_signal_1271, sbox_inst_21_T3}), .b ({new_AGEMA_signal_1558, sbox_inst_21_n17}), .c ({new_AGEMA_signal_1760, sbox_inst_21_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U6 ( .a ({new_AGEMA_signal_1272, sbox_inst_21_T4}), .b ({new_AGEMA_signal_1270, sbox_inst_21_T2}), .c ({new_AGEMA_signal_1556, sbox_inst_21_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U5 ( .a ({new_AGEMA_signal_1269, sbox_inst_21_T1}), .b ({input0_s1[86], input0_s0[86]}), .c ({new_AGEMA_signal_1557, sbox_inst_21_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U4 ( .a ({new_AGEMA_signal_1763, sbox_inst_21_n11}), .b ({input0_s1[85], input0_s0[85]}), .c ({output0_s1[21], output0_s0[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U3 ( .a ({input0_s1[87], input0_s0[87]}), .b ({new_AGEMA_signal_1558, sbox_inst_21_n17}), .c ({new_AGEMA_signal_1763, sbox_inst_21_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U2 ( .a ({input0_s1[84], input0_s0[84]}), .b ({new_AGEMA_signal_1266, sbox_inst_21_T0}), .c ({new_AGEMA_signal_1558, sbox_inst_21_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_t0_AND_U1 ( .a ({input0_s1[85], input0_s0[85]}), .b ({input0_s1[86], input0_s0[86]}), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_1266, sbox_inst_21_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_t1_AND_U1 ( .a ({input0_s1[84], input0_s0[84]}), .b ({input0_s1[87], input0_s0[87]}), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_1269, sbox_inst_21_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_t2_AND_U1 ( .a ({input0_s1[85], input0_s0[85]}), .b ({input0_s1[87], input0_s0[87]}), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_1270, sbox_inst_21_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_t3_AND_U1 ( .a ({input0_s1[86], input0_s0[86]}), .b ({input0_s1[87], input0_s0[87]}), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_1271, sbox_inst_21_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_t4_AND_U1 ( .a ({input0_s1[84], input0_s0[84]}), .b ({input0_s1[85], input0_s0[85]}), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_1272, sbox_inst_21_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U12 ( .a ({new_AGEMA_signal_1281, sbox_inst_20_T3}), .b ({new_AGEMA_signal_1563, sbox_inst_20_n17}), .c ({new_AGEMA_signal_1765, sbox_inst_20_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U6 ( .a ({new_AGEMA_signal_1282, sbox_inst_20_T4}), .b ({new_AGEMA_signal_1280, sbox_inst_20_T2}), .c ({new_AGEMA_signal_1561, sbox_inst_20_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U5 ( .a ({new_AGEMA_signal_1279, sbox_inst_20_T1}), .b ({input0_s1[82], input0_s0[82]}), .c ({new_AGEMA_signal_1562, sbox_inst_20_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U4 ( .a ({new_AGEMA_signal_1768, sbox_inst_20_n11}), .b ({input0_s1[81], input0_s0[81]}), .c ({output0_s1[20], output0_s0[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U3 ( .a ({input0_s1[83], input0_s0[83]}), .b ({new_AGEMA_signal_1563, sbox_inst_20_n17}), .c ({new_AGEMA_signal_1768, sbox_inst_20_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U2 ( .a ({input0_s1[80], input0_s0[80]}), .b ({new_AGEMA_signal_1276, sbox_inst_20_T0}), .c ({new_AGEMA_signal_1563, sbox_inst_20_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_t0_AND_U1 ( .a ({input0_s1[81], input0_s0[81]}), .b ({input0_s1[82], input0_s0[82]}), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_1276, sbox_inst_20_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_t1_AND_U1 ( .a ({input0_s1[80], input0_s0[80]}), .b ({input0_s1[83], input0_s0[83]}), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_1279, sbox_inst_20_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_t2_AND_U1 ( .a ({input0_s1[81], input0_s0[81]}), .b ({input0_s1[83], input0_s0[83]}), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_1280, sbox_inst_20_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_t3_AND_U1 ( .a ({input0_s1[82], input0_s0[82]}), .b ({input0_s1[83], input0_s0[83]}), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_1281, sbox_inst_20_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_t4_AND_U1 ( .a ({input0_s1[80], input0_s0[80]}), .b ({input0_s1[81], input0_s0[81]}), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_1282, sbox_inst_20_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U12 ( .a ({new_AGEMA_signal_1291, sbox_inst_19_T3}), .b ({new_AGEMA_signal_1568, sbox_inst_19_n17}), .c ({new_AGEMA_signal_1770, sbox_inst_19_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U6 ( .a ({new_AGEMA_signal_1292, sbox_inst_19_T4}), .b ({new_AGEMA_signal_1290, sbox_inst_19_T2}), .c ({new_AGEMA_signal_1566, sbox_inst_19_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U5 ( .a ({new_AGEMA_signal_1289, sbox_inst_19_T1}), .b ({input0_s1[78], input0_s0[78]}), .c ({new_AGEMA_signal_1567, sbox_inst_19_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U4 ( .a ({new_AGEMA_signal_1773, sbox_inst_19_n11}), .b ({input0_s1[77], input0_s0[77]}), .c ({output0_s1[19], output0_s0[19]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U3 ( .a ({input0_s1[79], input0_s0[79]}), .b ({new_AGEMA_signal_1568, sbox_inst_19_n17}), .c ({new_AGEMA_signal_1773, sbox_inst_19_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U2 ( .a ({input0_s1[76], input0_s0[76]}), .b ({new_AGEMA_signal_1286, sbox_inst_19_T0}), .c ({new_AGEMA_signal_1568, sbox_inst_19_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_t0_AND_U1 ( .a ({input0_s1[77], input0_s0[77]}), .b ({input0_s1[78], input0_s0[78]}), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_1286, sbox_inst_19_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_t1_AND_U1 ( .a ({input0_s1[76], input0_s0[76]}), .b ({input0_s1[79], input0_s0[79]}), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_1289, sbox_inst_19_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_t2_AND_U1 ( .a ({input0_s1[77], input0_s0[77]}), .b ({input0_s1[79], input0_s0[79]}), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_1290, sbox_inst_19_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_t3_AND_U1 ( .a ({input0_s1[78], input0_s0[78]}), .b ({input0_s1[79], input0_s0[79]}), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_1291, sbox_inst_19_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_t4_AND_U1 ( .a ({input0_s1[76], input0_s0[76]}), .b ({input0_s1[77], input0_s0[77]}), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_1292, sbox_inst_19_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U12 ( .a ({new_AGEMA_signal_1301, sbox_inst_18_T3}), .b ({new_AGEMA_signal_1573, sbox_inst_18_n17}), .c ({new_AGEMA_signal_1775, sbox_inst_18_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U6 ( .a ({new_AGEMA_signal_1302, sbox_inst_18_T4}), .b ({new_AGEMA_signal_1300, sbox_inst_18_T2}), .c ({new_AGEMA_signal_1571, sbox_inst_18_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U5 ( .a ({new_AGEMA_signal_1299, sbox_inst_18_T1}), .b ({input0_s1[74], input0_s0[74]}), .c ({new_AGEMA_signal_1572, sbox_inst_18_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U4 ( .a ({new_AGEMA_signal_1778, sbox_inst_18_n11}), .b ({input0_s1[73], input0_s0[73]}), .c ({output0_s1[18], output0_s0[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U3 ( .a ({input0_s1[75], input0_s0[75]}), .b ({new_AGEMA_signal_1573, sbox_inst_18_n17}), .c ({new_AGEMA_signal_1778, sbox_inst_18_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U2 ( .a ({input0_s1[72], input0_s0[72]}), .b ({new_AGEMA_signal_1296, sbox_inst_18_T0}), .c ({new_AGEMA_signal_1573, sbox_inst_18_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_t0_AND_U1 ( .a ({input0_s1[73], input0_s0[73]}), .b ({input0_s1[74], input0_s0[74]}), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_1296, sbox_inst_18_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_t1_AND_U1 ( .a ({input0_s1[72], input0_s0[72]}), .b ({input0_s1[75], input0_s0[75]}), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_1299, sbox_inst_18_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_t2_AND_U1 ( .a ({input0_s1[73], input0_s0[73]}), .b ({input0_s1[75], input0_s0[75]}), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_1300, sbox_inst_18_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_t3_AND_U1 ( .a ({input0_s1[74], input0_s0[74]}), .b ({input0_s1[75], input0_s0[75]}), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_1301, sbox_inst_18_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_t4_AND_U1 ( .a ({input0_s1[72], input0_s0[72]}), .b ({input0_s1[73], input0_s0[73]}), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_1302, sbox_inst_18_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U12 ( .a ({new_AGEMA_signal_1311, sbox_inst_17_T3}), .b ({new_AGEMA_signal_1578, sbox_inst_17_n17}), .c ({new_AGEMA_signal_1780, sbox_inst_17_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U6 ( .a ({new_AGEMA_signal_1312, sbox_inst_17_T4}), .b ({new_AGEMA_signal_1310, sbox_inst_17_T2}), .c ({new_AGEMA_signal_1576, sbox_inst_17_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U5 ( .a ({new_AGEMA_signal_1309, sbox_inst_17_T1}), .b ({input0_s1[70], input0_s0[70]}), .c ({new_AGEMA_signal_1577, sbox_inst_17_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U4 ( .a ({new_AGEMA_signal_1783, sbox_inst_17_n11}), .b ({input0_s1[69], input0_s0[69]}), .c ({output0_s1[17], output0_s0[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U3 ( .a ({input0_s1[71], input0_s0[71]}), .b ({new_AGEMA_signal_1578, sbox_inst_17_n17}), .c ({new_AGEMA_signal_1783, sbox_inst_17_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U2 ( .a ({input0_s1[68], input0_s0[68]}), .b ({new_AGEMA_signal_1306, sbox_inst_17_T0}), .c ({new_AGEMA_signal_1578, sbox_inst_17_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_t0_AND_U1 ( .a ({input0_s1[69], input0_s0[69]}), .b ({input0_s1[70], input0_s0[70]}), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_1306, sbox_inst_17_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_t1_AND_U1 ( .a ({input0_s1[68], input0_s0[68]}), .b ({input0_s1[71], input0_s0[71]}), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_1309, sbox_inst_17_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_t2_AND_U1 ( .a ({input0_s1[69], input0_s0[69]}), .b ({input0_s1[71], input0_s0[71]}), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_1310, sbox_inst_17_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_t3_AND_U1 ( .a ({input0_s1[70], input0_s0[70]}), .b ({input0_s1[71], input0_s0[71]}), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_1311, sbox_inst_17_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_t4_AND_U1 ( .a ({input0_s1[68], input0_s0[68]}), .b ({input0_s1[69], input0_s0[69]}), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_1312, sbox_inst_17_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U12 ( .a ({new_AGEMA_signal_1321, sbox_inst_16_T3}), .b ({new_AGEMA_signal_1583, sbox_inst_16_n17}), .c ({new_AGEMA_signal_1785, sbox_inst_16_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U6 ( .a ({new_AGEMA_signal_1322, sbox_inst_16_T4}), .b ({new_AGEMA_signal_1320, sbox_inst_16_T2}), .c ({new_AGEMA_signal_1581, sbox_inst_16_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U5 ( .a ({new_AGEMA_signal_1319, sbox_inst_16_T1}), .b ({input0_s1[66], input0_s0[66]}), .c ({new_AGEMA_signal_1582, sbox_inst_16_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U4 ( .a ({new_AGEMA_signal_1788, sbox_inst_16_n11}), .b ({input0_s1[65], input0_s0[65]}), .c ({output0_s1[16], output0_s0[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U3 ( .a ({input0_s1[67], input0_s0[67]}), .b ({new_AGEMA_signal_1583, sbox_inst_16_n17}), .c ({new_AGEMA_signal_1788, sbox_inst_16_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U2 ( .a ({input0_s1[64], input0_s0[64]}), .b ({new_AGEMA_signal_1316, sbox_inst_16_T0}), .c ({new_AGEMA_signal_1583, sbox_inst_16_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_t0_AND_U1 ( .a ({input0_s1[65], input0_s0[65]}), .b ({input0_s1[66], input0_s0[66]}), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_1316, sbox_inst_16_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_t1_AND_U1 ( .a ({input0_s1[64], input0_s0[64]}), .b ({input0_s1[67], input0_s0[67]}), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_1319, sbox_inst_16_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_t2_AND_U1 ( .a ({input0_s1[65], input0_s0[65]}), .b ({input0_s1[67], input0_s0[67]}), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_1320, sbox_inst_16_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_t3_AND_U1 ( .a ({input0_s1[66], input0_s0[66]}), .b ({input0_s1[67], input0_s0[67]}), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_1321, sbox_inst_16_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_t4_AND_U1 ( .a ({input0_s1[64], input0_s0[64]}), .b ({input0_s1[65], input0_s0[65]}), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_1322, sbox_inst_16_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U12 ( .a ({new_AGEMA_signal_1331, sbox_inst_15_T3}), .b ({new_AGEMA_signal_1588, sbox_inst_15_n17}), .c ({new_AGEMA_signal_1790, sbox_inst_15_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U6 ( .a ({new_AGEMA_signal_1332, sbox_inst_15_T4}), .b ({new_AGEMA_signal_1330, sbox_inst_15_T2}), .c ({new_AGEMA_signal_1586, sbox_inst_15_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U5 ( .a ({new_AGEMA_signal_1329, sbox_inst_15_T1}), .b ({input0_s1[62], input0_s0[62]}), .c ({new_AGEMA_signal_1587, sbox_inst_15_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U4 ( .a ({new_AGEMA_signal_1793, sbox_inst_15_n11}), .b ({input0_s1[61], input0_s0[61]}), .c ({output0_s1[15], output0_s0[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U3 ( .a ({input0_s1[63], input0_s0[63]}), .b ({new_AGEMA_signal_1588, sbox_inst_15_n17}), .c ({new_AGEMA_signal_1793, sbox_inst_15_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U2 ( .a ({input0_s1[60], input0_s0[60]}), .b ({new_AGEMA_signal_1326, sbox_inst_15_T0}), .c ({new_AGEMA_signal_1588, sbox_inst_15_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_t0_AND_U1 ( .a ({input0_s1[61], input0_s0[61]}), .b ({input0_s1[62], input0_s0[62]}), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_1326, sbox_inst_15_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_t1_AND_U1 ( .a ({input0_s1[60], input0_s0[60]}), .b ({input0_s1[63], input0_s0[63]}), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_1329, sbox_inst_15_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_t2_AND_U1 ( .a ({input0_s1[61], input0_s0[61]}), .b ({input0_s1[63], input0_s0[63]}), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_1330, sbox_inst_15_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_t3_AND_U1 ( .a ({input0_s1[62], input0_s0[62]}), .b ({input0_s1[63], input0_s0[63]}), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_1331, sbox_inst_15_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_t4_AND_U1 ( .a ({input0_s1[60], input0_s0[60]}), .b ({input0_s1[61], input0_s0[61]}), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_1332, sbox_inst_15_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U12 ( .a ({new_AGEMA_signal_1341, sbox_inst_14_T3}), .b ({new_AGEMA_signal_1593, sbox_inst_14_n17}), .c ({new_AGEMA_signal_1795, sbox_inst_14_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U6 ( .a ({new_AGEMA_signal_1342, sbox_inst_14_T4}), .b ({new_AGEMA_signal_1340, sbox_inst_14_T2}), .c ({new_AGEMA_signal_1591, sbox_inst_14_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U5 ( .a ({new_AGEMA_signal_1339, sbox_inst_14_T1}), .b ({input0_s1[58], input0_s0[58]}), .c ({new_AGEMA_signal_1592, sbox_inst_14_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U4 ( .a ({new_AGEMA_signal_1798, sbox_inst_14_n11}), .b ({input0_s1[57], input0_s0[57]}), .c ({output0_s1[14], output0_s0[14]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U3 ( .a ({input0_s1[59], input0_s0[59]}), .b ({new_AGEMA_signal_1593, sbox_inst_14_n17}), .c ({new_AGEMA_signal_1798, sbox_inst_14_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U2 ( .a ({input0_s1[56], input0_s0[56]}), .b ({new_AGEMA_signal_1336, sbox_inst_14_T0}), .c ({new_AGEMA_signal_1593, sbox_inst_14_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_t0_AND_U1 ( .a ({input0_s1[57], input0_s0[57]}), .b ({input0_s1[58], input0_s0[58]}), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_1336, sbox_inst_14_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_t1_AND_U1 ( .a ({input0_s1[56], input0_s0[56]}), .b ({input0_s1[59], input0_s0[59]}), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_1339, sbox_inst_14_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_t2_AND_U1 ( .a ({input0_s1[57], input0_s0[57]}), .b ({input0_s1[59], input0_s0[59]}), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_1340, sbox_inst_14_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_t3_AND_U1 ( .a ({input0_s1[58], input0_s0[58]}), .b ({input0_s1[59], input0_s0[59]}), .clk (clk), .r (Fresh[128]), .c ({new_AGEMA_signal_1341, sbox_inst_14_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_t4_AND_U1 ( .a ({input0_s1[56], input0_s0[56]}), .b ({input0_s1[57], input0_s0[57]}), .clk (clk), .r (Fresh[129]), .c ({new_AGEMA_signal_1342, sbox_inst_14_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U12 ( .a ({new_AGEMA_signal_1351, sbox_inst_13_T3}), .b ({new_AGEMA_signal_1598, sbox_inst_13_n17}), .c ({new_AGEMA_signal_1800, sbox_inst_13_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U6 ( .a ({new_AGEMA_signal_1352, sbox_inst_13_T4}), .b ({new_AGEMA_signal_1350, sbox_inst_13_T2}), .c ({new_AGEMA_signal_1596, sbox_inst_13_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U5 ( .a ({new_AGEMA_signal_1349, sbox_inst_13_T1}), .b ({input0_s1[54], input0_s0[54]}), .c ({new_AGEMA_signal_1597, sbox_inst_13_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U4 ( .a ({new_AGEMA_signal_1803, sbox_inst_13_n11}), .b ({input0_s1[53], input0_s0[53]}), .c ({output0_s1[13], output0_s0[13]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U3 ( .a ({input0_s1[55], input0_s0[55]}), .b ({new_AGEMA_signal_1598, sbox_inst_13_n17}), .c ({new_AGEMA_signal_1803, sbox_inst_13_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U2 ( .a ({input0_s1[52], input0_s0[52]}), .b ({new_AGEMA_signal_1346, sbox_inst_13_T0}), .c ({new_AGEMA_signal_1598, sbox_inst_13_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_t0_AND_U1 ( .a ({input0_s1[53], input0_s0[53]}), .b ({input0_s1[54], input0_s0[54]}), .clk (clk), .r (Fresh[130]), .c ({new_AGEMA_signal_1346, sbox_inst_13_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_t1_AND_U1 ( .a ({input0_s1[52], input0_s0[52]}), .b ({input0_s1[55], input0_s0[55]}), .clk (clk), .r (Fresh[131]), .c ({new_AGEMA_signal_1349, sbox_inst_13_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_t2_AND_U1 ( .a ({input0_s1[53], input0_s0[53]}), .b ({input0_s1[55], input0_s0[55]}), .clk (clk), .r (Fresh[132]), .c ({new_AGEMA_signal_1350, sbox_inst_13_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_t3_AND_U1 ( .a ({input0_s1[54], input0_s0[54]}), .b ({input0_s1[55], input0_s0[55]}), .clk (clk), .r (Fresh[133]), .c ({new_AGEMA_signal_1351, sbox_inst_13_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_t4_AND_U1 ( .a ({input0_s1[52], input0_s0[52]}), .b ({input0_s1[53], input0_s0[53]}), .clk (clk), .r (Fresh[134]), .c ({new_AGEMA_signal_1352, sbox_inst_13_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U12 ( .a ({new_AGEMA_signal_1361, sbox_inst_12_T3}), .b ({new_AGEMA_signal_1603, sbox_inst_12_n17}), .c ({new_AGEMA_signal_1805, sbox_inst_12_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U6 ( .a ({new_AGEMA_signal_1362, sbox_inst_12_T4}), .b ({new_AGEMA_signal_1360, sbox_inst_12_T2}), .c ({new_AGEMA_signal_1601, sbox_inst_12_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U5 ( .a ({new_AGEMA_signal_1359, sbox_inst_12_T1}), .b ({input0_s1[50], input0_s0[50]}), .c ({new_AGEMA_signal_1602, sbox_inst_12_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U4 ( .a ({new_AGEMA_signal_1808, sbox_inst_12_n11}), .b ({input0_s1[49], input0_s0[49]}), .c ({output0_s1[12], output0_s0[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U3 ( .a ({input0_s1[51], input0_s0[51]}), .b ({new_AGEMA_signal_1603, sbox_inst_12_n17}), .c ({new_AGEMA_signal_1808, sbox_inst_12_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U2 ( .a ({input0_s1[48], input0_s0[48]}), .b ({new_AGEMA_signal_1356, sbox_inst_12_T0}), .c ({new_AGEMA_signal_1603, sbox_inst_12_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_t0_AND_U1 ( .a ({input0_s1[49], input0_s0[49]}), .b ({input0_s1[50], input0_s0[50]}), .clk (clk), .r (Fresh[135]), .c ({new_AGEMA_signal_1356, sbox_inst_12_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_t1_AND_U1 ( .a ({input0_s1[48], input0_s0[48]}), .b ({input0_s1[51], input0_s0[51]}), .clk (clk), .r (Fresh[136]), .c ({new_AGEMA_signal_1359, sbox_inst_12_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_t2_AND_U1 ( .a ({input0_s1[49], input0_s0[49]}), .b ({input0_s1[51], input0_s0[51]}), .clk (clk), .r (Fresh[137]), .c ({new_AGEMA_signal_1360, sbox_inst_12_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_t3_AND_U1 ( .a ({input0_s1[50], input0_s0[50]}), .b ({input0_s1[51], input0_s0[51]}), .clk (clk), .r (Fresh[138]), .c ({new_AGEMA_signal_1361, sbox_inst_12_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_t4_AND_U1 ( .a ({input0_s1[48], input0_s0[48]}), .b ({input0_s1[49], input0_s0[49]}), .clk (clk), .r (Fresh[139]), .c ({new_AGEMA_signal_1362, sbox_inst_12_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U12 ( .a ({new_AGEMA_signal_1371, sbox_inst_11_T3}), .b ({new_AGEMA_signal_1608, sbox_inst_11_n17}), .c ({new_AGEMA_signal_1810, sbox_inst_11_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U6 ( .a ({new_AGEMA_signal_1372, sbox_inst_11_T4}), .b ({new_AGEMA_signal_1370, sbox_inst_11_T2}), .c ({new_AGEMA_signal_1606, sbox_inst_11_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U5 ( .a ({new_AGEMA_signal_1369, sbox_inst_11_T1}), .b ({input0_s1[46], input0_s0[46]}), .c ({new_AGEMA_signal_1607, sbox_inst_11_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U4 ( .a ({new_AGEMA_signal_1813, sbox_inst_11_n11}), .b ({input0_s1[45], input0_s0[45]}), .c ({output0_s1[11], output0_s0[11]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U3 ( .a ({input0_s1[47], input0_s0[47]}), .b ({new_AGEMA_signal_1608, sbox_inst_11_n17}), .c ({new_AGEMA_signal_1813, sbox_inst_11_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U2 ( .a ({input0_s1[44], input0_s0[44]}), .b ({new_AGEMA_signal_1366, sbox_inst_11_T0}), .c ({new_AGEMA_signal_1608, sbox_inst_11_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_t0_AND_U1 ( .a ({input0_s1[45], input0_s0[45]}), .b ({input0_s1[46], input0_s0[46]}), .clk (clk), .r (Fresh[140]), .c ({new_AGEMA_signal_1366, sbox_inst_11_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_t1_AND_U1 ( .a ({input0_s1[44], input0_s0[44]}), .b ({input0_s1[47], input0_s0[47]}), .clk (clk), .r (Fresh[141]), .c ({new_AGEMA_signal_1369, sbox_inst_11_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_t2_AND_U1 ( .a ({input0_s1[45], input0_s0[45]}), .b ({input0_s1[47], input0_s0[47]}), .clk (clk), .r (Fresh[142]), .c ({new_AGEMA_signal_1370, sbox_inst_11_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_t3_AND_U1 ( .a ({input0_s1[46], input0_s0[46]}), .b ({input0_s1[47], input0_s0[47]}), .clk (clk), .r (Fresh[143]), .c ({new_AGEMA_signal_1371, sbox_inst_11_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_t4_AND_U1 ( .a ({input0_s1[44], input0_s0[44]}), .b ({input0_s1[45], input0_s0[45]}), .clk (clk), .r (Fresh[144]), .c ({new_AGEMA_signal_1372, sbox_inst_11_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U12 ( .a ({new_AGEMA_signal_1381, sbox_inst_10_T3}), .b ({new_AGEMA_signal_1613, sbox_inst_10_n17}), .c ({new_AGEMA_signal_1815, sbox_inst_10_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U6 ( .a ({new_AGEMA_signal_1382, sbox_inst_10_T4}), .b ({new_AGEMA_signal_1380, sbox_inst_10_T2}), .c ({new_AGEMA_signal_1611, sbox_inst_10_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U5 ( .a ({new_AGEMA_signal_1379, sbox_inst_10_T1}), .b ({input0_s1[42], input0_s0[42]}), .c ({new_AGEMA_signal_1612, sbox_inst_10_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U4 ( .a ({new_AGEMA_signal_1818, sbox_inst_10_n11}), .b ({input0_s1[41], input0_s0[41]}), .c ({output0_s1[10], output0_s0[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U3 ( .a ({input0_s1[43], input0_s0[43]}), .b ({new_AGEMA_signal_1613, sbox_inst_10_n17}), .c ({new_AGEMA_signal_1818, sbox_inst_10_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U2 ( .a ({input0_s1[40], input0_s0[40]}), .b ({new_AGEMA_signal_1376, sbox_inst_10_T0}), .c ({new_AGEMA_signal_1613, sbox_inst_10_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_t0_AND_U1 ( .a ({input0_s1[41], input0_s0[41]}), .b ({input0_s1[42], input0_s0[42]}), .clk (clk), .r (Fresh[145]), .c ({new_AGEMA_signal_1376, sbox_inst_10_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_t1_AND_U1 ( .a ({input0_s1[40], input0_s0[40]}), .b ({input0_s1[43], input0_s0[43]}), .clk (clk), .r (Fresh[146]), .c ({new_AGEMA_signal_1379, sbox_inst_10_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_t2_AND_U1 ( .a ({input0_s1[41], input0_s0[41]}), .b ({input0_s1[43], input0_s0[43]}), .clk (clk), .r (Fresh[147]), .c ({new_AGEMA_signal_1380, sbox_inst_10_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_t3_AND_U1 ( .a ({input0_s1[42], input0_s0[42]}), .b ({input0_s1[43], input0_s0[43]}), .clk (clk), .r (Fresh[148]), .c ({new_AGEMA_signal_1381, sbox_inst_10_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_t4_AND_U1 ( .a ({input0_s1[40], input0_s0[40]}), .b ({input0_s1[41], input0_s0[41]}), .clk (clk), .r (Fresh[149]), .c ({new_AGEMA_signal_1382, sbox_inst_10_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U12 ( .a ({new_AGEMA_signal_1391, sbox_inst_9_T3}), .b ({new_AGEMA_signal_1618, sbox_inst_9_n17}), .c ({new_AGEMA_signal_1820, sbox_inst_9_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U6 ( .a ({new_AGEMA_signal_1392, sbox_inst_9_T4}), .b ({new_AGEMA_signal_1390, sbox_inst_9_T2}), .c ({new_AGEMA_signal_1616, sbox_inst_9_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U5 ( .a ({new_AGEMA_signal_1389, sbox_inst_9_T1}), .b ({input0_s1[38], input0_s0[38]}), .c ({new_AGEMA_signal_1617, sbox_inst_9_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U4 ( .a ({new_AGEMA_signal_1823, sbox_inst_9_n11}), .b ({input0_s1[37], input0_s0[37]}), .c ({output0_s1[9], output0_s0[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U3 ( .a ({input0_s1[39], input0_s0[39]}), .b ({new_AGEMA_signal_1618, sbox_inst_9_n17}), .c ({new_AGEMA_signal_1823, sbox_inst_9_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U2 ( .a ({input0_s1[36], input0_s0[36]}), .b ({new_AGEMA_signal_1386, sbox_inst_9_T0}), .c ({new_AGEMA_signal_1618, sbox_inst_9_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_t0_AND_U1 ( .a ({input0_s1[37], input0_s0[37]}), .b ({input0_s1[38], input0_s0[38]}), .clk (clk), .r (Fresh[150]), .c ({new_AGEMA_signal_1386, sbox_inst_9_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_t1_AND_U1 ( .a ({input0_s1[36], input0_s0[36]}), .b ({input0_s1[39], input0_s0[39]}), .clk (clk), .r (Fresh[151]), .c ({new_AGEMA_signal_1389, sbox_inst_9_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_t2_AND_U1 ( .a ({input0_s1[37], input0_s0[37]}), .b ({input0_s1[39], input0_s0[39]}), .clk (clk), .r (Fresh[152]), .c ({new_AGEMA_signal_1390, sbox_inst_9_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_t3_AND_U1 ( .a ({input0_s1[38], input0_s0[38]}), .b ({input0_s1[39], input0_s0[39]}), .clk (clk), .r (Fresh[153]), .c ({new_AGEMA_signal_1391, sbox_inst_9_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_t4_AND_U1 ( .a ({input0_s1[36], input0_s0[36]}), .b ({input0_s1[37], input0_s0[37]}), .clk (clk), .r (Fresh[154]), .c ({new_AGEMA_signal_1392, sbox_inst_9_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U12 ( .a ({new_AGEMA_signal_1401, sbox_inst_8_T3}), .b ({new_AGEMA_signal_1623, sbox_inst_8_n17}), .c ({new_AGEMA_signal_1825, sbox_inst_8_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U6 ( .a ({new_AGEMA_signal_1402, sbox_inst_8_T4}), .b ({new_AGEMA_signal_1400, sbox_inst_8_T2}), .c ({new_AGEMA_signal_1621, sbox_inst_8_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U5 ( .a ({new_AGEMA_signal_1399, sbox_inst_8_T1}), .b ({input0_s1[34], input0_s0[34]}), .c ({new_AGEMA_signal_1622, sbox_inst_8_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U4 ( .a ({new_AGEMA_signal_1828, sbox_inst_8_n11}), .b ({input0_s1[33], input0_s0[33]}), .c ({output0_s1[8], output0_s0[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U3 ( .a ({input0_s1[35], input0_s0[35]}), .b ({new_AGEMA_signal_1623, sbox_inst_8_n17}), .c ({new_AGEMA_signal_1828, sbox_inst_8_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U2 ( .a ({input0_s1[32], input0_s0[32]}), .b ({new_AGEMA_signal_1396, sbox_inst_8_T0}), .c ({new_AGEMA_signal_1623, sbox_inst_8_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_t0_AND_U1 ( .a ({input0_s1[33], input0_s0[33]}), .b ({input0_s1[34], input0_s0[34]}), .clk (clk), .r (Fresh[155]), .c ({new_AGEMA_signal_1396, sbox_inst_8_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_t1_AND_U1 ( .a ({input0_s1[32], input0_s0[32]}), .b ({input0_s1[35], input0_s0[35]}), .clk (clk), .r (Fresh[156]), .c ({new_AGEMA_signal_1399, sbox_inst_8_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_t2_AND_U1 ( .a ({input0_s1[33], input0_s0[33]}), .b ({input0_s1[35], input0_s0[35]}), .clk (clk), .r (Fresh[157]), .c ({new_AGEMA_signal_1400, sbox_inst_8_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_t3_AND_U1 ( .a ({input0_s1[34], input0_s0[34]}), .b ({input0_s1[35], input0_s0[35]}), .clk (clk), .r (Fresh[158]), .c ({new_AGEMA_signal_1401, sbox_inst_8_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_t4_AND_U1 ( .a ({input0_s1[32], input0_s0[32]}), .b ({input0_s1[33], input0_s0[33]}), .clk (clk), .r (Fresh[159]), .c ({new_AGEMA_signal_1402, sbox_inst_8_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U12 ( .a ({new_AGEMA_signal_1411, sbox_inst_7_T3}), .b ({new_AGEMA_signal_1628, sbox_inst_7_n17}), .c ({new_AGEMA_signal_1830, sbox_inst_7_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U6 ( .a ({new_AGEMA_signal_1412, sbox_inst_7_T4}), .b ({new_AGEMA_signal_1410, sbox_inst_7_T2}), .c ({new_AGEMA_signal_1626, sbox_inst_7_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U5 ( .a ({new_AGEMA_signal_1409, sbox_inst_7_T1}), .b ({input0_s1[30], input0_s0[30]}), .c ({new_AGEMA_signal_1627, sbox_inst_7_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U4 ( .a ({new_AGEMA_signal_1833, sbox_inst_7_n11}), .b ({input0_s1[29], input0_s0[29]}), .c ({output0_s1[7], output0_s0[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U3 ( .a ({input0_s1[31], input0_s0[31]}), .b ({new_AGEMA_signal_1628, sbox_inst_7_n17}), .c ({new_AGEMA_signal_1833, sbox_inst_7_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U2 ( .a ({input0_s1[28], input0_s0[28]}), .b ({new_AGEMA_signal_1406, sbox_inst_7_T0}), .c ({new_AGEMA_signal_1628, sbox_inst_7_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_t0_AND_U1 ( .a ({input0_s1[29], input0_s0[29]}), .b ({input0_s1[30], input0_s0[30]}), .clk (clk), .r (Fresh[160]), .c ({new_AGEMA_signal_1406, sbox_inst_7_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_t1_AND_U1 ( .a ({input0_s1[28], input0_s0[28]}), .b ({input0_s1[31], input0_s0[31]}), .clk (clk), .r (Fresh[161]), .c ({new_AGEMA_signal_1409, sbox_inst_7_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_t2_AND_U1 ( .a ({input0_s1[29], input0_s0[29]}), .b ({input0_s1[31], input0_s0[31]}), .clk (clk), .r (Fresh[162]), .c ({new_AGEMA_signal_1410, sbox_inst_7_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_t3_AND_U1 ( .a ({input0_s1[30], input0_s0[30]}), .b ({input0_s1[31], input0_s0[31]}), .clk (clk), .r (Fresh[163]), .c ({new_AGEMA_signal_1411, sbox_inst_7_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_t4_AND_U1 ( .a ({input0_s1[28], input0_s0[28]}), .b ({input0_s1[29], input0_s0[29]}), .clk (clk), .r (Fresh[164]), .c ({new_AGEMA_signal_1412, sbox_inst_7_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U12 ( .a ({new_AGEMA_signal_1421, sbox_inst_6_T3}), .b ({new_AGEMA_signal_1633, sbox_inst_6_n17}), .c ({new_AGEMA_signal_1835, sbox_inst_6_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U6 ( .a ({new_AGEMA_signal_1422, sbox_inst_6_T4}), .b ({new_AGEMA_signal_1420, sbox_inst_6_T2}), .c ({new_AGEMA_signal_1631, sbox_inst_6_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U5 ( .a ({new_AGEMA_signal_1419, sbox_inst_6_T1}), .b ({input0_s1[26], input0_s0[26]}), .c ({new_AGEMA_signal_1632, sbox_inst_6_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U4 ( .a ({new_AGEMA_signal_1838, sbox_inst_6_n11}), .b ({input0_s1[25], input0_s0[25]}), .c ({output0_s1[6], output0_s0[6]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U3 ( .a ({input0_s1[27], input0_s0[27]}), .b ({new_AGEMA_signal_1633, sbox_inst_6_n17}), .c ({new_AGEMA_signal_1838, sbox_inst_6_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U2 ( .a ({input0_s1[24], input0_s0[24]}), .b ({new_AGEMA_signal_1416, sbox_inst_6_T0}), .c ({new_AGEMA_signal_1633, sbox_inst_6_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_t0_AND_U1 ( .a ({input0_s1[25], input0_s0[25]}), .b ({input0_s1[26], input0_s0[26]}), .clk (clk), .r (Fresh[165]), .c ({new_AGEMA_signal_1416, sbox_inst_6_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_t1_AND_U1 ( .a ({input0_s1[24], input0_s0[24]}), .b ({input0_s1[27], input0_s0[27]}), .clk (clk), .r (Fresh[166]), .c ({new_AGEMA_signal_1419, sbox_inst_6_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_t2_AND_U1 ( .a ({input0_s1[25], input0_s0[25]}), .b ({input0_s1[27], input0_s0[27]}), .clk (clk), .r (Fresh[167]), .c ({new_AGEMA_signal_1420, sbox_inst_6_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_t3_AND_U1 ( .a ({input0_s1[26], input0_s0[26]}), .b ({input0_s1[27], input0_s0[27]}), .clk (clk), .r (Fresh[168]), .c ({new_AGEMA_signal_1421, sbox_inst_6_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_t4_AND_U1 ( .a ({input0_s1[24], input0_s0[24]}), .b ({input0_s1[25], input0_s0[25]}), .clk (clk), .r (Fresh[169]), .c ({new_AGEMA_signal_1422, sbox_inst_6_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U12 ( .a ({new_AGEMA_signal_1431, sbox_inst_5_T3}), .b ({new_AGEMA_signal_1638, sbox_inst_5_n17}), .c ({new_AGEMA_signal_1840, sbox_inst_5_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U6 ( .a ({new_AGEMA_signal_1432, sbox_inst_5_T4}), .b ({new_AGEMA_signal_1430, sbox_inst_5_T2}), .c ({new_AGEMA_signal_1636, sbox_inst_5_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U5 ( .a ({new_AGEMA_signal_1429, sbox_inst_5_T1}), .b ({input0_s1[22], input0_s0[22]}), .c ({new_AGEMA_signal_1637, sbox_inst_5_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U4 ( .a ({new_AGEMA_signal_1843, sbox_inst_5_n11}), .b ({input0_s1[21], input0_s0[21]}), .c ({output0_s1[5], output0_s0[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U3 ( .a ({input0_s1[23], input0_s0[23]}), .b ({new_AGEMA_signal_1638, sbox_inst_5_n17}), .c ({new_AGEMA_signal_1843, sbox_inst_5_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U2 ( .a ({input0_s1[20], input0_s0[20]}), .b ({new_AGEMA_signal_1426, sbox_inst_5_T0}), .c ({new_AGEMA_signal_1638, sbox_inst_5_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_t0_AND_U1 ( .a ({input0_s1[21], input0_s0[21]}), .b ({input0_s1[22], input0_s0[22]}), .clk (clk), .r (Fresh[170]), .c ({new_AGEMA_signal_1426, sbox_inst_5_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_t1_AND_U1 ( .a ({input0_s1[20], input0_s0[20]}), .b ({input0_s1[23], input0_s0[23]}), .clk (clk), .r (Fresh[171]), .c ({new_AGEMA_signal_1429, sbox_inst_5_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_t2_AND_U1 ( .a ({input0_s1[21], input0_s0[21]}), .b ({input0_s1[23], input0_s0[23]}), .clk (clk), .r (Fresh[172]), .c ({new_AGEMA_signal_1430, sbox_inst_5_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_t3_AND_U1 ( .a ({input0_s1[22], input0_s0[22]}), .b ({input0_s1[23], input0_s0[23]}), .clk (clk), .r (Fresh[173]), .c ({new_AGEMA_signal_1431, sbox_inst_5_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_t4_AND_U1 ( .a ({input0_s1[20], input0_s0[20]}), .b ({input0_s1[21], input0_s0[21]}), .clk (clk), .r (Fresh[174]), .c ({new_AGEMA_signal_1432, sbox_inst_5_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U12 ( .a ({new_AGEMA_signal_1441, sbox_inst_4_T3}), .b ({new_AGEMA_signal_1643, sbox_inst_4_n17}), .c ({new_AGEMA_signal_1845, sbox_inst_4_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U6 ( .a ({new_AGEMA_signal_1442, sbox_inst_4_T4}), .b ({new_AGEMA_signal_1440, sbox_inst_4_T2}), .c ({new_AGEMA_signal_1641, sbox_inst_4_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U5 ( .a ({new_AGEMA_signal_1439, sbox_inst_4_T1}), .b ({input0_s1[18], input0_s0[18]}), .c ({new_AGEMA_signal_1642, sbox_inst_4_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U4 ( .a ({new_AGEMA_signal_1848, sbox_inst_4_n11}), .b ({input0_s1[17], input0_s0[17]}), .c ({output0_s1[4], output0_s0[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U3 ( .a ({input0_s1[19], input0_s0[19]}), .b ({new_AGEMA_signal_1643, sbox_inst_4_n17}), .c ({new_AGEMA_signal_1848, sbox_inst_4_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U2 ( .a ({input0_s1[16], input0_s0[16]}), .b ({new_AGEMA_signal_1436, sbox_inst_4_T0}), .c ({new_AGEMA_signal_1643, sbox_inst_4_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_t0_AND_U1 ( .a ({input0_s1[17], input0_s0[17]}), .b ({input0_s1[18], input0_s0[18]}), .clk (clk), .r (Fresh[175]), .c ({new_AGEMA_signal_1436, sbox_inst_4_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_t1_AND_U1 ( .a ({input0_s1[16], input0_s0[16]}), .b ({input0_s1[19], input0_s0[19]}), .clk (clk), .r (Fresh[176]), .c ({new_AGEMA_signal_1439, sbox_inst_4_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_t2_AND_U1 ( .a ({input0_s1[17], input0_s0[17]}), .b ({input0_s1[19], input0_s0[19]}), .clk (clk), .r (Fresh[177]), .c ({new_AGEMA_signal_1440, sbox_inst_4_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_t3_AND_U1 ( .a ({input0_s1[18], input0_s0[18]}), .b ({input0_s1[19], input0_s0[19]}), .clk (clk), .r (Fresh[178]), .c ({new_AGEMA_signal_1441, sbox_inst_4_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_t4_AND_U1 ( .a ({input0_s1[16], input0_s0[16]}), .b ({input0_s1[17], input0_s0[17]}), .clk (clk), .r (Fresh[179]), .c ({new_AGEMA_signal_1442, sbox_inst_4_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U12 ( .a ({new_AGEMA_signal_1451, sbox_inst_3_T3}), .b ({new_AGEMA_signal_1648, sbox_inst_3_n17}), .c ({new_AGEMA_signal_1850, sbox_inst_3_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U6 ( .a ({new_AGEMA_signal_1452, sbox_inst_3_T4}), .b ({new_AGEMA_signal_1450, sbox_inst_3_T2}), .c ({new_AGEMA_signal_1646, sbox_inst_3_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U5 ( .a ({new_AGEMA_signal_1449, sbox_inst_3_T1}), .b ({input0_s1[14], input0_s0[14]}), .c ({new_AGEMA_signal_1647, sbox_inst_3_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U4 ( .a ({new_AGEMA_signal_1853, sbox_inst_3_n11}), .b ({input0_s1[13], input0_s0[13]}), .c ({output0_s1[3], output0_s0[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U3 ( .a ({input0_s1[15], input0_s0[15]}), .b ({new_AGEMA_signal_1648, sbox_inst_3_n17}), .c ({new_AGEMA_signal_1853, sbox_inst_3_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U2 ( .a ({input0_s1[12], input0_s0[12]}), .b ({new_AGEMA_signal_1446, sbox_inst_3_T0}), .c ({new_AGEMA_signal_1648, sbox_inst_3_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_t0_AND_U1 ( .a ({input0_s1[13], input0_s0[13]}), .b ({input0_s1[14], input0_s0[14]}), .clk (clk), .r (Fresh[180]), .c ({new_AGEMA_signal_1446, sbox_inst_3_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_t1_AND_U1 ( .a ({input0_s1[12], input0_s0[12]}), .b ({input0_s1[15], input0_s0[15]}), .clk (clk), .r (Fresh[181]), .c ({new_AGEMA_signal_1449, sbox_inst_3_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_t2_AND_U1 ( .a ({input0_s1[13], input0_s0[13]}), .b ({input0_s1[15], input0_s0[15]}), .clk (clk), .r (Fresh[182]), .c ({new_AGEMA_signal_1450, sbox_inst_3_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_t3_AND_U1 ( .a ({input0_s1[14], input0_s0[14]}), .b ({input0_s1[15], input0_s0[15]}), .clk (clk), .r (Fresh[183]), .c ({new_AGEMA_signal_1451, sbox_inst_3_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_t4_AND_U1 ( .a ({input0_s1[12], input0_s0[12]}), .b ({input0_s1[13], input0_s0[13]}), .clk (clk), .r (Fresh[184]), .c ({new_AGEMA_signal_1452, sbox_inst_3_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U12 ( .a ({new_AGEMA_signal_1461, sbox_inst_2_T3}), .b ({new_AGEMA_signal_1653, sbox_inst_2_n17}), .c ({new_AGEMA_signal_1855, sbox_inst_2_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U6 ( .a ({new_AGEMA_signal_1462, sbox_inst_2_T4}), .b ({new_AGEMA_signal_1460, sbox_inst_2_T2}), .c ({new_AGEMA_signal_1651, sbox_inst_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U5 ( .a ({new_AGEMA_signal_1459, sbox_inst_2_T1}), .b ({input0_s1[10], input0_s0[10]}), .c ({new_AGEMA_signal_1652, sbox_inst_2_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U4 ( .a ({new_AGEMA_signal_1858, sbox_inst_2_n11}), .b ({input0_s1[9], input0_s0[9]}), .c ({output0_s1[2], output0_s0[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U3 ( .a ({input0_s1[11], input0_s0[11]}), .b ({new_AGEMA_signal_1653, sbox_inst_2_n17}), .c ({new_AGEMA_signal_1858, sbox_inst_2_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U2 ( .a ({input0_s1[8], input0_s0[8]}), .b ({new_AGEMA_signal_1456, sbox_inst_2_T0}), .c ({new_AGEMA_signal_1653, sbox_inst_2_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_t0_AND_U1 ( .a ({input0_s1[9], input0_s0[9]}), .b ({input0_s1[10], input0_s0[10]}), .clk (clk), .r (Fresh[185]), .c ({new_AGEMA_signal_1456, sbox_inst_2_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_t1_AND_U1 ( .a ({input0_s1[8], input0_s0[8]}), .b ({input0_s1[11], input0_s0[11]}), .clk (clk), .r (Fresh[186]), .c ({new_AGEMA_signal_1459, sbox_inst_2_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_t2_AND_U1 ( .a ({input0_s1[9], input0_s0[9]}), .b ({input0_s1[11], input0_s0[11]}), .clk (clk), .r (Fresh[187]), .c ({new_AGEMA_signal_1460, sbox_inst_2_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_t3_AND_U1 ( .a ({input0_s1[10], input0_s0[10]}), .b ({input0_s1[11], input0_s0[11]}), .clk (clk), .r (Fresh[188]), .c ({new_AGEMA_signal_1461, sbox_inst_2_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_t4_AND_U1 ( .a ({input0_s1[8], input0_s0[8]}), .b ({input0_s1[9], input0_s0[9]}), .clk (clk), .r (Fresh[189]), .c ({new_AGEMA_signal_1462, sbox_inst_2_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U12 ( .a ({new_AGEMA_signal_1661, sbox_inst_1_T3}), .b ({new_AGEMA_signal_1861, sbox_inst_1_n17}), .c ({new_AGEMA_signal_2024, sbox_inst_1_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U6 ( .a ({new_AGEMA_signal_1662, sbox_inst_1_T4}), .b ({new_AGEMA_signal_1660, sbox_inst_1_T2}), .c ({new_AGEMA_signal_1859, sbox_inst_1_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U5 ( .a ({new_AGEMA_signal_1659, sbox_inst_1_T1}), .b ({new_AGEMA_signal_1084, input_array_6}), .c ({new_AGEMA_signal_1860, sbox_inst_1_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U4 ( .a ({new_AGEMA_signal_2027, sbox_inst_1_n11}), .b ({new_AGEMA_signal_1082, input_array_5}), .c ({output0_s1[1], output0_s0[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U3 ( .a ({input0_s1[7], input0_s0[7]}), .b ({new_AGEMA_signal_1861, sbox_inst_1_n17}), .c ({new_AGEMA_signal_2027, sbox_inst_1_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U2 ( .a ({new_AGEMA_signal_1086, input_array_4}), .b ({new_AGEMA_signal_1657, sbox_inst_1_T0}), .c ({new_AGEMA_signal_1861, sbox_inst_1_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_t0_AND_U1 ( .a ({new_AGEMA_signal_1082, input_array_5}), .b ({new_AGEMA_signal_1084, input_array_6}), .clk (clk), .r (Fresh[190]), .c ({new_AGEMA_signal_1657, sbox_inst_1_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_t1_AND_U1 ( .a ({new_AGEMA_signal_1086, input_array_4}), .b ({input0_s1[7], input0_s0[7]}), .clk (clk), .r (Fresh[191]), .c ({new_AGEMA_signal_1659, sbox_inst_1_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_t2_AND_U1 ( .a ({new_AGEMA_signal_1082, input_array_5}), .b ({input0_s1[7], input0_s0[7]}), .clk (clk), .r (Fresh[192]), .c ({new_AGEMA_signal_1660, sbox_inst_1_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_t3_AND_U1 ( .a ({new_AGEMA_signal_1084, input_array_6}), .b ({input0_s1[7], input0_s0[7]}), .clk (clk), .r (Fresh[193]), .c ({new_AGEMA_signal_1661, sbox_inst_1_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_t4_AND_U1 ( .a ({new_AGEMA_signal_1086, input_array_4}), .b ({new_AGEMA_signal_1082, input_array_5}), .clk (clk), .r (Fresh[194]), .c ({new_AGEMA_signal_1662, sbox_inst_1_T4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U12 ( .a ({new_AGEMA_signal_1667, sbox_inst_0_T3}), .b ({new_AGEMA_signal_1866, sbox_inst_0_n17}), .c ({new_AGEMA_signal_2029, sbox_inst_0_n19}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U6 ( .a ({new_AGEMA_signal_1668, sbox_inst_0_T4}), .b ({new_AGEMA_signal_1666, sbox_inst_0_T2}), .c ({new_AGEMA_signal_1864, sbox_inst_0_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U5 ( .a ({new_AGEMA_signal_1665, sbox_inst_0_T1}), .b ({new_AGEMA_signal_1090, input_array_2}), .c ({new_AGEMA_signal_1865, sbox_inst_0_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U4 ( .a ({new_AGEMA_signal_2032, sbox_inst_0_n11}), .b ({new_AGEMA_signal_1076, input_array_1}), .c ({output0_s1[0], output0_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U3 ( .a ({new_AGEMA_signal_1088, input_array_3}), .b ({new_AGEMA_signal_1866, sbox_inst_0_n17}), .c ({new_AGEMA_signal_2032, sbox_inst_0_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U2 ( .a ({new_AGEMA_signal_1092, input_array_0}), .b ({new_AGEMA_signal_1664, sbox_inst_0_T0}), .c ({new_AGEMA_signal_1866, sbox_inst_0_n17}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_t0_AND_U1 ( .a ({new_AGEMA_signal_1076, input_array_1}), .b ({new_AGEMA_signal_1090, input_array_2}), .clk (clk), .r (Fresh[195]), .c ({new_AGEMA_signal_1664, sbox_inst_0_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_t1_AND_U1 ( .a ({new_AGEMA_signal_1092, input_array_0}), .b ({new_AGEMA_signal_1088, input_array_3}), .clk (clk), .r (Fresh[196]), .c ({new_AGEMA_signal_1665, sbox_inst_0_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_t2_AND_U1 ( .a ({new_AGEMA_signal_1076, input_array_1}), .b ({new_AGEMA_signal_1088, input_array_3}), .clk (clk), .r (Fresh[197]), .c ({new_AGEMA_signal_1666, sbox_inst_0_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_t3_AND_U1 ( .a ({new_AGEMA_signal_1090, input_array_2}), .b ({new_AGEMA_signal_1088, input_array_3}), .clk (clk), .r (Fresh[198]), .c ({new_AGEMA_signal_1667, sbox_inst_0_T3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_t4_AND_U1 ( .a ({new_AGEMA_signal_1092, input_array_0}), .b ({new_AGEMA_signal_1076, input_array_1}), .clk (clk), .r (Fresh[199]), .c ({new_AGEMA_signal_1668, sbox_inst_0_T4}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U15 ( .a ({new_AGEMA_signal_1466, sbox_inst_39_T2}), .b ({new_AGEMA_signal_2033, sbox_inst_39_n20}), .c ({output0_s1[79], output0_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U14 ( .a ({new_AGEMA_signal_1870, sbox_inst_39_n19}), .b ({new_AGEMA_signal_1869, sbox_inst_39_n18}), .c ({new_AGEMA_signal_2033, sbox_inst_39_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U13 ( .a ({new_AGEMA_signal_1465, sbox_inst_39_T1}), .b ({new_AGEMA_signal_1672, sbox_inst_39_T5}), .c ({new_AGEMA_signal_1869, sbox_inst_39_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U11 ( .a ({new_AGEMA_signal_1078, input_array[157]}), .b ({new_AGEMA_signal_1871, sbox_inst_39_n16}), .c ({output0_s1[119], output0_s0[119]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U10 ( .a ({new_AGEMA_signal_1670, sbox_inst_39_n15}), .b ({new_AGEMA_signal_1672, sbox_inst_39_T5}), .c ({new_AGEMA_signal_1871, sbox_inst_39_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U9 ( .a ({new_AGEMA_signal_1670, sbox_inst_39_n15}), .b ({new_AGEMA_signal_2035, sbox_inst_39_n14}), .c ({output0_s1[159], output0_s0[159]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U8 ( .a ({new_AGEMA_signal_1669, sbox_inst_39_n13}), .b ({new_AGEMA_signal_1872, sbox_inst_39_n12}), .c ({new_AGEMA_signal_2035, sbox_inst_39_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_U7 ( .a ({new_AGEMA_signal_1673, sbox_inst_39_T6}), .b ({new_AGEMA_signal_1094, input_array[159]}), .c ({new_AGEMA_signal_1872, sbox_inst_39_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_t5_AND_U1 ( .a ({new_AGEMA_signal_1078, input_array[157]}), .b ({new_AGEMA_signal_1467, sbox_inst_39_T3}), .clk (clk), .r (Fresh[200]), .c ({new_AGEMA_signal_1672, sbox_inst_39_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_39_t6_AND_U1 ( .a ({new_AGEMA_signal_1463, sbox_inst_39_L0}), .b ({new_AGEMA_signal_1465, sbox_inst_39_T1}), .clk (clk), .r (Fresh[201]), .c ({new_AGEMA_signal_1673, sbox_inst_39_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U15 ( .a ({new_AGEMA_signal_1473, sbox_inst_38_T2}), .b ({new_AGEMA_signal_2037, sbox_inst_38_n20}), .c ({output0_s1[78], output0_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U14 ( .a ({new_AGEMA_signal_1875, sbox_inst_38_n19}), .b ({new_AGEMA_signal_1874, sbox_inst_38_n18}), .c ({new_AGEMA_signal_2037, sbox_inst_38_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U13 ( .a ({new_AGEMA_signal_1472, sbox_inst_38_T1}), .b ({new_AGEMA_signal_1677, sbox_inst_38_T5}), .c ({new_AGEMA_signal_1874, sbox_inst_38_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U11 ( .a ({new_AGEMA_signal_1080, input_array[153]}), .b ({new_AGEMA_signal_1876, sbox_inst_38_n16}), .c ({output0_s1[118], output0_s0[118]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U10 ( .a ({new_AGEMA_signal_1675, sbox_inst_38_n15}), .b ({new_AGEMA_signal_1677, sbox_inst_38_T5}), .c ({new_AGEMA_signal_1876, sbox_inst_38_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U9 ( .a ({new_AGEMA_signal_1675, sbox_inst_38_n15}), .b ({new_AGEMA_signal_2039, sbox_inst_38_n14}), .c ({output0_s1[158], output0_s0[158]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U8 ( .a ({new_AGEMA_signal_1674, sbox_inst_38_n13}), .b ({new_AGEMA_signal_1877, sbox_inst_38_n12}), .c ({new_AGEMA_signal_2039, sbox_inst_38_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_U7 ( .a ({new_AGEMA_signal_1678, sbox_inst_38_T6}), .b ({new_AGEMA_signal_1100, input_array[155]}), .c ({new_AGEMA_signal_1877, sbox_inst_38_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_t5_AND_U1 ( .a ({new_AGEMA_signal_1080, input_array[153]}), .b ({new_AGEMA_signal_1474, sbox_inst_38_T3}), .clk (clk), .r (Fresh[202]), .c ({new_AGEMA_signal_1677, sbox_inst_38_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_38_t6_AND_U1 ( .a ({new_AGEMA_signal_1469, sbox_inst_38_L0}), .b ({new_AGEMA_signal_1472, sbox_inst_38_T1}), .clk (clk), .r (Fresh[203]), .c ({new_AGEMA_signal_1678, sbox_inst_38_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U15 ( .a ({new_AGEMA_signal_1110, sbox_inst_37_T2}), .b ({new_AGEMA_signal_1879, sbox_inst_37_n20}), .c ({output0_s1[77], output0_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U14 ( .a ({new_AGEMA_signal_1680, sbox_inst_37_n19}), .b ({new_AGEMA_signal_1679, sbox_inst_37_n18}), .c ({new_AGEMA_signal_1879, sbox_inst_37_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U13 ( .a ({new_AGEMA_signal_1109, sbox_inst_37_T1}), .b ({new_AGEMA_signal_1479, sbox_inst_37_T5}), .c ({new_AGEMA_signal_1679, sbox_inst_37_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U11 ( .a ({input0_s1[149], input0_s0[149]}), .b ({new_AGEMA_signal_1681, sbox_inst_37_n16}), .c ({output0_s1[117], output0_s0[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U10 ( .a ({new_AGEMA_signal_1477, sbox_inst_37_n15}), .b ({new_AGEMA_signal_1479, sbox_inst_37_T5}), .c ({new_AGEMA_signal_1681, sbox_inst_37_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U9 ( .a ({new_AGEMA_signal_1477, sbox_inst_37_n15}), .b ({new_AGEMA_signal_1881, sbox_inst_37_n14}), .c ({output0_s1[157], output0_s0[157]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U8 ( .a ({new_AGEMA_signal_1476, sbox_inst_37_n13}), .b ({new_AGEMA_signal_1682, sbox_inst_37_n12}), .c ({new_AGEMA_signal_1881, sbox_inst_37_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_U7 ( .a ({new_AGEMA_signal_1480, sbox_inst_37_T6}), .b ({input0_s1[151], input0_s0[151]}), .c ({new_AGEMA_signal_1682, sbox_inst_37_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_t5_AND_U1 ( .a ({input0_s1[149], input0_s0[149]}), .b ({new_AGEMA_signal_1111, sbox_inst_37_T3}), .clk (clk), .r (Fresh[204]), .c ({new_AGEMA_signal_1479, sbox_inst_37_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_37_t6_AND_U1 ( .a ({new_AGEMA_signal_1105, sbox_inst_37_L0}), .b ({new_AGEMA_signal_1109, sbox_inst_37_T1}), .clk (clk), .r (Fresh[205]), .c ({new_AGEMA_signal_1480, sbox_inst_37_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U15 ( .a ({new_AGEMA_signal_1120, sbox_inst_36_T2}), .b ({new_AGEMA_signal_1883, sbox_inst_36_n20}), .c ({output0_s1[76], output0_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U14 ( .a ({new_AGEMA_signal_1685, sbox_inst_36_n19}), .b ({new_AGEMA_signal_1684, sbox_inst_36_n18}), .c ({new_AGEMA_signal_1883, sbox_inst_36_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U13 ( .a ({new_AGEMA_signal_1119, sbox_inst_36_T1}), .b ({new_AGEMA_signal_1484, sbox_inst_36_T5}), .c ({new_AGEMA_signal_1684, sbox_inst_36_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U11 ( .a ({input0_s1[145], input0_s0[145]}), .b ({new_AGEMA_signal_1686, sbox_inst_36_n16}), .c ({output0_s1[116], output0_s0[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U10 ( .a ({new_AGEMA_signal_1482, sbox_inst_36_n15}), .b ({new_AGEMA_signal_1484, sbox_inst_36_T5}), .c ({new_AGEMA_signal_1686, sbox_inst_36_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U9 ( .a ({new_AGEMA_signal_1482, sbox_inst_36_n15}), .b ({new_AGEMA_signal_1885, sbox_inst_36_n14}), .c ({output0_s1[156], output0_s0[156]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U8 ( .a ({new_AGEMA_signal_1481, sbox_inst_36_n13}), .b ({new_AGEMA_signal_1687, sbox_inst_36_n12}), .c ({new_AGEMA_signal_1885, sbox_inst_36_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_U7 ( .a ({new_AGEMA_signal_1485, sbox_inst_36_T6}), .b ({input0_s1[147], input0_s0[147]}), .c ({new_AGEMA_signal_1687, sbox_inst_36_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_t5_AND_U1 ( .a ({input0_s1[145], input0_s0[145]}), .b ({new_AGEMA_signal_1121, sbox_inst_36_T3}), .clk (clk), .r (Fresh[206]), .c ({new_AGEMA_signal_1484, sbox_inst_36_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_36_t6_AND_U1 ( .a ({new_AGEMA_signal_1115, sbox_inst_36_L0}), .b ({new_AGEMA_signal_1119, sbox_inst_36_T1}), .clk (clk), .r (Fresh[207]), .c ({new_AGEMA_signal_1485, sbox_inst_36_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U15 ( .a ({new_AGEMA_signal_1130, sbox_inst_35_T2}), .b ({new_AGEMA_signal_1887, sbox_inst_35_n20}), .c ({output0_s1[75], output0_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U14 ( .a ({new_AGEMA_signal_1690, sbox_inst_35_n19}), .b ({new_AGEMA_signal_1689, sbox_inst_35_n18}), .c ({new_AGEMA_signal_1887, sbox_inst_35_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U13 ( .a ({new_AGEMA_signal_1129, sbox_inst_35_T1}), .b ({new_AGEMA_signal_1489, sbox_inst_35_T5}), .c ({new_AGEMA_signal_1689, sbox_inst_35_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U11 ( .a ({input0_s1[141], input0_s0[141]}), .b ({new_AGEMA_signal_1691, sbox_inst_35_n16}), .c ({output0_s1[115], output0_s0[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U10 ( .a ({new_AGEMA_signal_1487, sbox_inst_35_n15}), .b ({new_AGEMA_signal_1489, sbox_inst_35_T5}), .c ({new_AGEMA_signal_1691, sbox_inst_35_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U9 ( .a ({new_AGEMA_signal_1487, sbox_inst_35_n15}), .b ({new_AGEMA_signal_1889, sbox_inst_35_n14}), .c ({output0_s1[155], output0_s0[155]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U8 ( .a ({new_AGEMA_signal_1486, sbox_inst_35_n13}), .b ({new_AGEMA_signal_1692, sbox_inst_35_n12}), .c ({new_AGEMA_signal_1889, sbox_inst_35_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_U7 ( .a ({new_AGEMA_signal_1490, sbox_inst_35_T6}), .b ({input0_s1[143], input0_s0[143]}), .c ({new_AGEMA_signal_1692, sbox_inst_35_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_t5_AND_U1 ( .a ({input0_s1[141], input0_s0[141]}), .b ({new_AGEMA_signal_1131, sbox_inst_35_T3}), .clk (clk), .r (Fresh[208]), .c ({new_AGEMA_signal_1489, sbox_inst_35_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_35_t6_AND_U1 ( .a ({new_AGEMA_signal_1125, sbox_inst_35_L0}), .b ({new_AGEMA_signal_1129, sbox_inst_35_T1}), .clk (clk), .r (Fresh[209]), .c ({new_AGEMA_signal_1490, sbox_inst_35_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U15 ( .a ({new_AGEMA_signal_1140, sbox_inst_34_T2}), .b ({new_AGEMA_signal_1891, sbox_inst_34_n20}), .c ({output0_s1[74], output0_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U14 ( .a ({new_AGEMA_signal_1695, sbox_inst_34_n19}), .b ({new_AGEMA_signal_1694, sbox_inst_34_n18}), .c ({new_AGEMA_signal_1891, sbox_inst_34_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U13 ( .a ({new_AGEMA_signal_1139, sbox_inst_34_T1}), .b ({new_AGEMA_signal_1494, sbox_inst_34_T5}), .c ({new_AGEMA_signal_1694, sbox_inst_34_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U11 ( .a ({input0_s1[137], input0_s0[137]}), .b ({new_AGEMA_signal_1696, sbox_inst_34_n16}), .c ({output0_s1[114], output0_s0[114]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U10 ( .a ({new_AGEMA_signal_1492, sbox_inst_34_n15}), .b ({new_AGEMA_signal_1494, sbox_inst_34_T5}), .c ({new_AGEMA_signal_1696, sbox_inst_34_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U9 ( .a ({new_AGEMA_signal_1492, sbox_inst_34_n15}), .b ({new_AGEMA_signal_1893, sbox_inst_34_n14}), .c ({output0_s1[154], output0_s0[154]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U8 ( .a ({new_AGEMA_signal_1491, sbox_inst_34_n13}), .b ({new_AGEMA_signal_1697, sbox_inst_34_n12}), .c ({new_AGEMA_signal_1893, sbox_inst_34_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_U7 ( .a ({new_AGEMA_signal_1495, sbox_inst_34_T6}), .b ({input0_s1[139], input0_s0[139]}), .c ({new_AGEMA_signal_1697, sbox_inst_34_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_t5_AND_U1 ( .a ({input0_s1[137], input0_s0[137]}), .b ({new_AGEMA_signal_1141, sbox_inst_34_T3}), .clk (clk), .r (Fresh[210]), .c ({new_AGEMA_signal_1494, sbox_inst_34_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_34_t6_AND_U1 ( .a ({new_AGEMA_signal_1135, sbox_inst_34_L0}), .b ({new_AGEMA_signal_1139, sbox_inst_34_T1}), .clk (clk), .r (Fresh[211]), .c ({new_AGEMA_signal_1495, sbox_inst_34_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U15 ( .a ({new_AGEMA_signal_1150, sbox_inst_33_T2}), .b ({new_AGEMA_signal_1895, sbox_inst_33_n20}), .c ({output0_s1[73], output0_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U14 ( .a ({new_AGEMA_signal_1700, sbox_inst_33_n19}), .b ({new_AGEMA_signal_1699, sbox_inst_33_n18}), .c ({new_AGEMA_signal_1895, sbox_inst_33_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U13 ( .a ({new_AGEMA_signal_1149, sbox_inst_33_T1}), .b ({new_AGEMA_signal_1499, sbox_inst_33_T5}), .c ({new_AGEMA_signal_1699, sbox_inst_33_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U11 ( .a ({input0_s1[133], input0_s0[133]}), .b ({new_AGEMA_signal_1701, sbox_inst_33_n16}), .c ({output0_s1[113], output0_s0[113]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U10 ( .a ({new_AGEMA_signal_1497, sbox_inst_33_n15}), .b ({new_AGEMA_signal_1499, sbox_inst_33_T5}), .c ({new_AGEMA_signal_1701, sbox_inst_33_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U9 ( .a ({new_AGEMA_signal_1497, sbox_inst_33_n15}), .b ({new_AGEMA_signal_1897, sbox_inst_33_n14}), .c ({output0_s1[153], output0_s0[153]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U8 ( .a ({new_AGEMA_signal_1496, sbox_inst_33_n13}), .b ({new_AGEMA_signal_1702, sbox_inst_33_n12}), .c ({new_AGEMA_signal_1897, sbox_inst_33_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_U7 ( .a ({new_AGEMA_signal_1500, sbox_inst_33_T6}), .b ({input0_s1[135], input0_s0[135]}), .c ({new_AGEMA_signal_1702, sbox_inst_33_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_t5_AND_U1 ( .a ({input0_s1[133], input0_s0[133]}), .b ({new_AGEMA_signal_1151, sbox_inst_33_T3}), .clk (clk), .r (Fresh[212]), .c ({new_AGEMA_signal_1499, sbox_inst_33_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_33_t6_AND_U1 ( .a ({new_AGEMA_signal_1145, sbox_inst_33_L0}), .b ({new_AGEMA_signal_1149, sbox_inst_33_T1}), .clk (clk), .r (Fresh[213]), .c ({new_AGEMA_signal_1500, sbox_inst_33_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U15 ( .a ({new_AGEMA_signal_1160, sbox_inst_32_T2}), .b ({new_AGEMA_signal_1899, sbox_inst_32_n20}), .c ({output0_s1[72], output0_s0[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U14 ( .a ({new_AGEMA_signal_1705, sbox_inst_32_n19}), .b ({new_AGEMA_signal_1704, sbox_inst_32_n18}), .c ({new_AGEMA_signal_1899, sbox_inst_32_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U13 ( .a ({new_AGEMA_signal_1159, sbox_inst_32_T1}), .b ({new_AGEMA_signal_1504, sbox_inst_32_T5}), .c ({new_AGEMA_signal_1704, sbox_inst_32_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U11 ( .a ({input0_s1[129], input0_s0[129]}), .b ({new_AGEMA_signal_1706, sbox_inst_32_n16}), .c ({output0_s1[112], output0_s0[112]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U10 ( .a ({new_AGEMA_signal_1502, sbox_inst_32_n15}), .b ({new_AGEMA_signal_1504, sbox_inst_32_T5}), .c ({new_AGEMA_signal_1706, sbox_inst_32_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U9 ( .a ({new_AGEMA_signal_1502, sbox_inst_32_n15}), .b ({new_AGEMA_signal_1901, sbox_inst_32_n14}), .c ({output0_s1[152], output0_s0[152]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U8 ( .a ({new_AGEMA_signal_1501, sbox_inst_32_n13}), .b ({new_AGEMA_signal_1707, sbox_inst_32_n12}), .c ({new_AGEMA_signal_1901, sbox_inst_32_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_U7 ( .a ({new_AGEMA_signal_1505, sbox_inst_32_T6}), .b ({input0_s1[131], input0_s0[131]}), .c ({new_AGEMA_signal_1707, sbox_inst_32_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_t5_AND_U1 ( .a ({input0_s1[129], input0_s0[129]}), .b ({new_AGEMA_signal_1161, sbox_inst_32_T3}), .clk (clk), .r (Fresh[214]), .c ({new_AGEMA_signal_1504, sbox_inst_32_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_32_t6_AND_U1 ( .a ({new_AGEMA_signal_1155, sbox_inst_32_L0}), .b ({new_AGEMA_signal_1159, sbox_inst_32_T1}), .clk (clk), .r (Fresh[215]), .c ({new_AGEMA_signal_1505, sbox_inst_32_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U15 ( .a ({new_AGEMA_signal_1170, sbox_inst_31_T2}), .b ({new_AGEMA_signal_1903, sbox_inst_31_n20}), .c ({output0_s1[71], output0_s0[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U14 ( .a ({new_AGEMA_signal_1710, sbox_inst_31_n19}), .b ({new_AGEMA_signal_1709, sbox_inst_31_n18}), .c ({new_AGEMA_signal_1903, sbox_inst_31_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U13 ( .a ({new_AGEMA_signal_1169, sbox_inst_31_T1}), .b ({new_AGEMA_signal_1509, sbox_inst_31_T5}), .c ({new_AGEMA_signal_1709, sbox_inst_31_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U11 ( .a ({input0_s1[125], input0_s0[125]}), .b ({new_AGEMA_signal_1711, sbox_inst_31_n16}), .c ({output0_s1[111], output0_s0[111]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U10 ( .a ({new_AGEMA_signal_1507, sbox_inst_31_n15}), .b ({new_AGEMA_signal_1509, sbox_inst_31_T5}), .c ({new_AGEMA_signal_1711, sbox_inst_31_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U9 ( .a ({new_AGEMA_signal_1507, sbox_inst_31_n15}), .b ({new_AGEMA_signal_1905, sbox_inst_31_n14}), .c ({output0_s1[151], output0_s0[151]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U8 ( .a ({new_AGEMA_signal_1506, sbox_inst_31_n13}), .b ({new_AGEMA_signal_1712, sbox_inst_31_n12}), .c ({new_AGEMA_signal_1905, sbox_inst_31_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_U7 ( .a ({new_AGEMA_signal_1510, sbox_inst_31_T6}), .b ({input0_s1[127], input0_s0[127]}), .c ({new_AGEMA_signal_1712, sbox_inst_31_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_t5_AND_U1 ( .a ({input0_s1[125], input0_s0[125]}), .b ({new_AGEMA_signal_1171, sbox_inst_31_T3}), .clk (clk), .r (Fresh[216]), .c ({new_AGEMA_signal_1509, sbox_inst_31_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_31_t6_AND_U1 ( .a ({new_AGEMA_signal_1165, sbox_inst_31_L0}), .b ({new_AGEMA_signal_1169, sbox_inst_31_T1}), .clk (clk), .r (Fresh[217]), .c ({new_AGEMA_signal_1510, sbox_inst_31_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U15 ( .a ({new_AGEMA_signal_1180, sbox_inst_30_T2}), .b ({new_AGEMA_signal_1907, sbox_inst_30_n20}), .c ({output0_s1[70], output0_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U14 ( .a ({new_AGEMA_signal_1715, sbox_inst_30_n19}), .b ({new_AGEMA_signal_1714, sbox_inst_30_n18}), .c ({new_AGEMA_signal_1907, sbox_inst_30_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U13 ( .a ({new_AGEMA_signal_1179, sbox_inst_30_T1}), .b ({new_AGEMA_signal_1514, sbox_inst_30_T5}), .c ({new_AGEMA_signal_1714, sbox_inst_30_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U11 ( .a ({input0_s1[121], input0_s0[121]}), .b ({new_AGEMA_signal_1716, sbox_inst_30_n16}), .c ({output0_s1[110], output0_s0[110]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U10 ( .a ({new_AGEMA_signal_1512, sbox_inst_30_n15}), .b ({new_AGEMA_signal_1514, sbox_inst_30_T5}), .c ({new_AGEMA_signal_1716, sbox_inst_30_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U9 ( .a ({new_AGEMA_signal_1512, sbox_inst_30_n15}), .b ({new_AGEMA_signal_1909, sbox_inst_30_n14}), .c ({output0_s1[150], output0_s0[150]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U8 ( .a ({new_AGEMA_signal_1511, sbox_inst_30_n13}), .b ({new_AGEMA_signal_1717, sbox_inst_30_n12}), .c ({new_AGEMA_signal_1909, sbox_inst_30_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_U7 ( .a ({new_AGEMA_signal_1515, sbox_inst_30_T6}), .b ({input0_s1[123], input0_s0[123]}), .c ({new_AGEMA_signal_1717, sbox_inst_30_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_t5_AND_U1 ( .a ({input0_s1[121], input0_s0[121]}), .b ({new_AGEMA_signal_1181, sbox_inst_30_T3}), .clk (clk), .r (Fresh[218]), .c ({new_AGEMA_signal_1514, sbox_inst_30_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_30_t6_AND_U1 ( .a ({new_AGEMA_signal_1175, sbox_inst_30_L0}), .b ({new_AGEMA_signal_1179, sbox_inst_30_T1}), .clk (clk), .r (Fresh[219]), .c ({new_AGEMA_signal_1515, sbox_inst_30_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U15 ( .a ({new_AGEMA_signal_1190, sbox_inst_29_T2}), .b ({new_AGEMA_signal_1911, sbox_inst_29_n20}), .c ({output0_s1[69], output0_s0[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U14 ( .a ({new_AGEMA_signal_1720, sbox_inst_29_n19}), .b ({new_AGEMA_signal_1719, sbox_inst_29_n18}), .c ({new_AGEMA_signal_1911, sbox_inst_29_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U13 ( .a ({new_AGEMA_signal_1189, sbox_inst_29_T1}), .b ({new_AGEMA_signal_1519, sbox_inst_29_T5}), .c ({new_AGEMA_signal_1719, sbox_inst_29_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U11 ( .a ({input0_s1[117], input0_s0[117]}), .b ({new_AGEMA_signal_1721, sbox_inst_29_n16}), .c ({output0_s1[109], output0_s0[109]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U10 ( .a ({new_AGEMA_signal_1517, sbox_inst_29_n15}), .b ({new_AGEMA_signal_1519, sbox_inst_29_T5}), .c ({new_AGEMA_signal_1721, sbox_inst_29_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U9 ( .a ({new_AGEMA_signal_1517, sbox_inst_29_n15}), .b ({new_AGEMA_signal_1913, sbox_inst_29_n14}), .c ({output0_s1[149], output0_s0[149]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U8 ( .a ({new_AGEMA_signal_1516, sbox_inst_29_n13}), .b ({new_AGEMA_signal_1722, sbox_inst_29_n12}), .c ({new_AGEMA_signal_1913, sbox_inst_29_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_U7 ( .a ({new_AGEMA_signal_1520, sbox_inst_29_T6}), .b ({input0_s1[119], input0_s0[119]}), .c ({new_AGEMA_signal_1722, sbox_inst_29_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_t5_AND_U1 ( .a ({input0_s1[117], input0_s0[117]}), .b ({new_AGEMA_signal_1191, sbox_inst_29_T3}), .clk (clk), .r (Fresh[220]), .c ({new_AGEMA_signal_1519, sbox_inst_29_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_29_t6_AND_U1 ( .a ({new_AGEMA_signal_1185, sbox_inst_29_L0}), .b ({new_AGEMA_signal_1189, sbox_inst_29_T1}), .clk (clk), .r (Fresh[221]), .c ({new_AGEMA_signal_1520, sbox_inst_29_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U15 ( .a ({new_AGEMA_signal_1200, sbox_inst_28_T2}), .b ({new_AGEMA_signal_1915, sbox_inst_28_n20}), .c ({output0_s1[68], output0_s0[68]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U14 ( .a ({new_AGEMA_signal_1725, sbox_inst_28_n19}), .b ({new_AGEMA_signal_1724, sbox_inst_28_n18}), .c ({new_AGEMA_signal_1915, sbox_inst_28_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U13 ( .a ({new_AGEMA_signal_1199, sbox_inst_28_T1}), .b ({new_AGEMA_signal_1524, sbox_inst_28_T5}), .c ({new_AGEMA_signal_1724, sbox_inst_28_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U11 ( .a ({input0_s1[113], input0_s0[113]}), .b ({new_AGEMA_signal_1726, sbox_inst_28_n16}), .c ({output0_s1[108], output0_s0[108]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U10 ( .a ({new_AGEMA_signal_1522, sbox_inst_28_n15}), .b ({new_AGEMA_signal_1524, sbox_inst_28_T5}), .c ({new_AGEMA_signal_1726, sbox_inst_28_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U9 ( .a ({new_AGEMA_signal_1522, sbox_inst_28_n15}), .b ({new_AGEMA_signal_1917, sbox_inst_28_n14}), .c ({output0_s1[148], output0_s0[148]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U8 ( .a ({new_AGEMA_signal_1521, sbox_inst_28_n13}), .b ({new_AGEMA_signal_1727, sbox_inst_28_n12}), .c ({new_AGEMA_signal_1917, sbox_inst_28_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_U7 ( .a ({new_AGEMA_signal_1525, sbox_inst_28_T6}), .b ({input0_s1[115], input0_s0[115]}), .c ({new_AGEMA_signal_1727, sbox_inst_28_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_t5_AND_U1 ( .a ({input0_s1[113], input0_s0[113]}), .b ({new_AGEMA_signal_1201, sbox_inst_28_T3}), .clk (clk), .r (Fresh[222]), .c ({new_AGEMA_signal_1524, sbox_inst_28_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_28_t6_AND_U1 ( .a ({new_AGEMA_signal_1195, sbox_inst_28_L0}), .b ({new_AGEMA_signal_1199, sbox_inst_28_T1}), .clk (clk), .r (Fresh[223]), .c ({new_AGEMA_signal_1525, sbox_inst_28_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U15 ( .a ({new_AGEMA_signal_1210, sbox_inst_27_T2}), .b ({new_AGEMA_signal_1919, sbox_inst_27_n20}), .c ({output0_s1[67], output0_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U14 ( .a ({new_AGEMA_signal_1730, sbox_inst_27_n19}), .b ({new_AGEMA_signal_1729, sbox_inst_27_n18}), .c ({new_AGEMA_signal_1919, sbox_inst_27_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U13 ( .a ({new_AGEMA_signal_1209, sbox_inst_27_T1}), .b ({new_AGEMA_signal_1529, sbox_inst_27_T5}), .c ({new_AGEMA_signal_1729, sbox_inst_27_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U11 ( .a ({input0_s1[109], input0_s0[109]}), .b ({new_AGEMA_signal_1731, sbox_inst_27_n16}), .c ({output0_s1[107], output0_s0[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U10 ( .a ({new_AGEMA_signal_1527, sbox_inst_27_n15}), .b ({new_AGEMA_signal_1529, sbox_inst_27_T5}), .c ({new_AGEMA_signal_1731, sbox_inst_27_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U9 ( .a ({new_AGEMA_signal_1527, sbox_inst_27_n15}), .b ({new_AGEMA_signal_1921, sbox_inst_27_n14}), .c ({output0_s1[147], output0_s0[147]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U8 ( .a ({new_AGEMA_signal_1526, sbox_inst_27_n13}), .b ({new_AGEMA_signal_1732, sbox_inst_27_n12}), .c ({new_AGEMA_signal_1921, sbox_inst_27_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_U7 ( .a ({new_AGEMA_signal_1530, sbox_inst_27_T6}), .b ({input0_s1[111], input0_s0[111]}), .c ({new_AGEMA_signal_1732, sbox_inst_27_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_t5_AND_U1 ( .a ({input0_s1[109], input0_s0[109]}), .b ({new_AGEMA_signal_1211, sbox_inst_27_T3}), .clk (clk), .r (Fresh[224]), .c ({new_AGEMA_signal_1529, sbox_inst_27_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_27_t6_AND_U1 ( .a ({new_AGEMA_signal_1205, sbox_inst_27_L0}), .b ({new_AGEMA_signal_1209, sbox_inst_27_T1}), .clk (clk), .r (Fresh[225]), .c ({new_AGEMA_signal_1530, sbox_inst_27_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U15 ( .a ({new_AGEMA_signal_1220, sbox_inst_26_T2}), .b ({new_AGEMA_signal_1923, sbox_inst_26_n20}), .c ({output0_s1[66], output0_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U14 ( .a ({new_AGEMA_signal_1735, sbox_inst_26_n19}), .b ({new_AGEMA_signal_1734, sbox_inst_26_n18}), .c ({new_AGEMA_signal_1923, sbox_inst_26_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U13 ( .a ({new_AGEMA_signal_1219, sbox_inst_26_T1}), .b ({new_AGEMA_signal_1534, sbox_inst_26_T5}), .c ({new_AGEMA_signal_1734, sbox_inst_26_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U11 ( .a ({input0_s1[105], input0_s0[105]}), .b ({new_AGEMA_signal_1736, sbox_inst_26_n16}), .c ({output0_s1[106], output0_s0[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U10 ( .a ({new_AGEMA_signal_1532, sbox_inst_26_n15}), .b ({new_AGEMA_signal_1534, sbox_inst_26_T5}), .c ({new_AGEMA_signal_1736, sbox_inst_26_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U9 ( .a ({new_AGEMA_signal_1532, sbox_inst_26_n15}), .b ({new_AGEMA_signal_1925, sbox_inst_26_n14}), .c ({output0_s1[146], output0_s0[146]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U8 ( .a ({new_AGEMA_signal_1531, sbox_inst_26_n13}), .b ({new_AGEMA_signal_1737, sbox_inst_26_n12}), .c ({new_AGEMA_signal_1925, sbox_inst_26_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_U7 ( .a ({new_AGEMA_signal_1535, sbox_inst_26_T6}), .b ({input0_s1[107], input0_s0[107]}), .c ({new_AGEMA_signal_1737, sbox_inst_26_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_t5_AND_U1 ( .a ({input0_s1[105], input0_s0[105]}), .b ({new_AGEMA_signal_1221, sbox_inst_26_T3}), .clk (clk), .r (Fresh[226]), .c ({new_AGEMA_signal_1534, sbox_inst_26_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_26_t6_AND_U1 ( .a ({new_AGEMA_signal_1215, sbox_inst_26_L0}), .b ({new_AGEMA_signal_1219, sbox_inst_26_T1}), .clk (clk), .r (Fresh[227]), .c ({new_AGEMA_signal_1535, sbox_inst_26_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U15 ( .a ({new_AGEMA_signal_1230, sbox_inst_25_T2}), .b ({new_AGEMA_signal_1927, sbox_inst_25_n20}), .c ({output0_s1[65], output0_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U14 ( .a ({new_AGEMA_signal_1740, sbox_inst_25_n19}), .b ({new_AGEMA_signal_1739, sbox_inst_25_n18}), .c ({new_AGEMA_signal_1927, sbox_inst_25_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U13 ( .a ({new_AGEMA_signal_1229, sbox_inst_25_T1}), .b ({new_AGEMA_signal_1539, sbox_inst_25_T5}), .c ({new_AGEMA_signal_1739, sbox_inst_25_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U11 ( .a ({input0_s1[101], input0_s0[101]}), .b ({new_AGEMA_signal_1741, sbox_inst_25_n16}), .c ({output0_s1[105], output0_s0[105]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U10 ( .a ({new_AGEMA_signal_1537, sbox_inst_25_n15}), .b ({new_AGEMA_signal_1539, sbox_inst_25_T5}), .c ({new_AGEMA_signal_1741, sbox_inst_25_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U9 ( .a ({new_AGEMA_signal_1537, sbox_inst_25_n15}), .b ({new_AGEMA_signal_1929, sbox_inst_25_n14}), .c ({output0_s1[145], output0_s0[145]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U8 ( .a ({new_AGEMA_signal_1536, sbox_inst_25_n13}), .b ({new_AGEMA_signal_1742, sbox_inst_25_n12}), .c ({new_AGEMA_signal_1929, sbox_inst_25_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_U7 ( .a ({new_AGEMA_signal_1540, sbox_inst_25_T6}), .b ({input0_s1[103], input0_s0[103]}), .c ({new_AGEMA_signal_1742, sbox_inst_25_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_t5_AND_U1 ( .a ({input0_s1[101], input0_s0[101]}), .b ({new_AGEMA_signal_1231, sbox_inst_25_T3}), .clk (clk), .r (Fresh[228]), .c ({new_AGEMA_signal_1539, sbox_inst_25_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_25_t6_AND_U1 ( .a ({new_AGEMA_signal_1225, sbox_inst_25_L0}), .b ({new_AGEMA_signal_1229, sbox_inst_25_T1}), .clk (clk), .r (Fresh[229]), .c ({new_AGEMA_signal_1540, sbox_inst_25_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U15 ( .a ({new_AGEMA_signal_1240, sbox_inst_24_T2}), .b ({new_AGEMA_signal_1931, sbox_inst_24_n20}), .c ({output0_s1[64], output0_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U14 ( .a ({new_AGEMA_signal_1745, sbox_inst_24_n19}), .b ({new_AGEMA_signal_1744, sbox_inst_24_n18}), .c ({new_AGEMA_signal_1931, sbox_inst_24_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U13 ( .a ({new_AGEMA_signal_1239, sbox_inst_24_T1}), .b ({new_AGEMA_signal_1544, sbox_inst_24_T5}), .c ({new_AGEMA_signal_1744, sbox_inst_24_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U11 ( .a ({input0_s1[97], input0_s0[97]}), .b ({new_AGEMA_signal_1746, sbox_inst_24_n16}), .c ({output0_s1[104], output0_s0[104]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U10 ( .a ({new_AGEMA_signal_1542, sbox_inst_24_n15}), .b ({new_AGEMA_signal_1544, sbox_inst_24_T5}), .c ({new_AGEMA_signal_1746, sbox_inst_24_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U9 ( .a ({new_AGEMA_signal_1542, sbox_inst_24_n15}), .b ({new_AGEMA_signal_1933, sbox_inst_24_n14}), .c ({output0_s1[144], output0_s0[144]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U8 ( .a ({new_AGEMA_signal_1541, sbox_inst_24_n13}), .b ({new_AGEMA_signal_1747, sbox_inst_24_n12}), .c ({new_AGEMA_signal_1933, sbox_inst_24_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_U7 ( .a ({new_AGEMA_signal_1545, sbox_inst_24_T6}), .b ({input0_s1[99], input0_s0[99]}), .c ({new_AGEMA_signal_1747, sbox_inst_24_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_t5_AND_U1 ( .a ({input0_s1[97], input0_s0[97]}), .b ({new_AGEMA_signal_1241, sbox_inst_24_T3}), .clk (clk), .r (Fresh[230]), .c ({new_AGEMA_signal_1544, sbox_inst_24_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_24_t6_AND_U1 ( .a ({new_AGEMA_signal_1235, sbox_inst_24_L0}), .b ({new_AGEMA_signal_1239, sbox_inst_24_T1}), .clk (clk), .r (Fresh[231]), .c ({new_AGEMA_signal_1545, sbox_inst_24_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U15 ( .a ({new_AGEMA_signal_1250, sbox_inst_23_T2}), .b ({new_AGEMA_signal_1935, sbox_inst_23_n20}), .c ({output0_s1[63], output0_s0[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U14 ( .a ({new_AGEMA_signal_1750, sbox_inst_23_n19}), .b ({new_AGEMA_signal_1749, sbox_inst_23_n18}), .c ({new_AGEMA_signal_1935, sbox_inst_23_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U13 ( .a ({new_AGEMA_signal_1249, sbox_inst_23_T1}), .b ({new_AGEMA_signal_1549, sbox_inst_23_T5}), .c ({new_AGEMA_signal_1749, sbox_inst_23_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U11 ( .a ({input0_s1[93], input0_s0[93]}), .b ({new_AGEMA_signal_1751, sbox_inst_23_n16}), .c ({output0_s1[103], output0_s0[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U10 ( .a ({new_AGEMA_signal_1547, sbox_inst_23_n15}), .b ({new_AGEMA_signal_1549, sbox_inst_23_T5}), .c ({new_AGEMA_signal_1751, sbox_inst_23_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U9 ( .a ({new_AGEMA_signal_1547, sbox_inst_23_n15}), .b ({new_AGEMA_signal_1937, sbox_inst_23_n14}), .c ({output0_s1[143], output0_s0[143]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U8 ( .a ({new_AGEMA_signal_1546, sbox_inst_23_n13}), .b ({new_AGEMA_signal_1752, sbox_inst_23_n12}), .c ({new_AGEMA_signal_1937, sbox_inst_23_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_U7 ( .a ({new_AGEMA_signal_1550, sbox_inst_23_T6}), .b ({input0_s1[95], input0_s0[95]}), .c ({new_AGEMA_signal_1752, sbox_inst_23_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_t5_AND_U1 ( .a ({input0_s1[93], input0_s0[93]}), .b ({new_AGEMA_signal_1251, sbox_inst_23_T3}), .clk (clk), .r (Fresh[232]), .c ({new_AGEMA_signal_1549, sbox_inst_23_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_23_t6_AND_U1 ( .a ({new_AGEMA_signal_1245, sbox_inst_23_L0}), .b ({new_AGEMA_signal_1249, sbox_inst_23_T1}), .clk (clk), .r (Fresh[233]), .c ({new_AGEMA_signal_1550, sbox_inst_23_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U15 ( .a ({new_AGEMA_signal_1260, sbox_inst_22_T2}), .b ({new_AGEMA_signal_1939, sbox_inst_22_n20}), .c ({output0_s1[62], output0_s0[62]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U14 ( .a ({new_AGEMA_signal_1755, sbox_inst_22_n19}), .b ({new_AGEMA_signal_1754, sbox_inst_22_n18}), .c ({new_AGEMA_signal_1939, sbox_inst_22_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U13 ( .a ({new_AGEMA_signal_1259, sbox_inst_22_T1}), .b ({new_AGEMA_signal_1554, sbox_inst_22_T5}), .c ({new_AGEMA_signal_1754, sbox_inst_22_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U11 ( .a ({input0_s1[89], input0_s0[89]}), .b ({new_AGEMA_signal_1756, sbox_inst_22_n16}), .c ({output0_s1[102], output0_s0[102]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U10 ( .a ({new_AGEMA_signal_1552, sbox_inst_22_n15}), .b ({new_AGEMA_signal_1554, sbox_inst_22_T5}), .c ({new_AGEMA_signal_1756, sbox_inst_22_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U9 ( .a ({new_AGEMA_signal_1552, sbox_inst_22_n15}), .b ({new_AGEMA_signal_1941, sbox_inst_22_n14}), .c ({output0_s1[142], output0_s0[142]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U8 ( .a ({new_AGEMA_signal_1551, sbox_inst_22_n13}), .b ({new_AGEMA_signal_1757, sbox_inst_22_n12}), .c ({new_AGEMA_signal_1941, sbox_inst_22_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_U7 ( .a ({new_AGEMA_signal_1555, sbox_inst_22_T6}), .b ({input0_s1[91], input0_s0[91]}), .c ({new_AGEMA_signal_1757, sbox_inst_22_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_t5_AND_U1 ( .a ({input0_s1[89], input0_s0[89]}), .b ({new_AGEMA_signal_1261, sbox_inst_22_T3}), .clk (clk), .r (Fresh[234]), .c ({new_AGEMA_signal_1554, sbox_inst_22_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_22_t6_AND_U1 ( .a ({new_AGEMA_signal_1255, sbox_inst_22_L0}), .b ({new_AGEMA_signal_1259, sbox_inst_22_T1}), .clk (clk), .r (Fresh[235]), .c ({new_AGEMA_signal_1555, sbox_inst_22_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U15 ( .a ({new_AGEMA_signal_1270, sbox_inst_21_T2}), .b ({new_AGEMA_signal_1943, sbox_inst_21_n20}), .c ({output0_s1[61], output0_s0[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U14 ( .a ({new_AGEMA_signal_1760, sbox_inst_21_n19}), .b ({new_AGEMA_signal_1759, sbox_inst_21_n18}), .c ({new_AGEMA_signal_1943, sbox_inst_21_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U13 ( .a ({new_AGEMA_signal_1269, sbox_inst_21_T1}), .b ({new_AGEMA_signal_1559, sbox_inst_21_T5}), .c ({new_AGEMA_signal_1759, sbox_inst_21_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U11 ( .a ({input0_s1[85], input0_s0[85]}), .b ({new_AGEMA_signal_1761, sbox_inst_21_n16}), .c ({output0_s1[101], output0_s0[101]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U10 ( .a ({new_AGEMA_signal_1557, sbox_inst_21_n15}), .b ({new_AGEMA_signal_1559, sbox_inst_21_T5}), .c ({new_AGEMA_signal_1761, sbox_inst_21_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U9 ( .a ({new_AGEMA_signal_1557, sbox_inst_21_n15}), .b ({new_AGEMA_signal_1945, sbox_inst_21_n14}), .c ({output0_s1[141], output0_s0[141]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U8 ( .a ({new_AGEMA_signal_1556, sbox_inst_21_n13}), .b ({new_AGEMA_signal_1762, sbox_inst_21_n12}), .c ({new_AGEMA_signal_1945, sbox_inst_21_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_U7 ( .a ({new_AGEMA_signal_1560, sbox_inst_21_T6}), .b ({input0_s1[87], input0_s0[87]}), .c ({new_AGEMA_signal_1762, sbox_inst_21_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_t5_AND_U1 ( .a ({input0_s1[85], input0_s0[85]}), .b ({new_AGEMA_signal_1271, sbox_inst_21_T3}), .clk (clk), .r (Fresh[236]), .c ({new_AGEMA_signal_1559, sbox_inst_21_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_21_t6_AND_U1 ( .a ({new_AGEMA_signal_1265, sbox_inst_21_L0}), .b ({new_AGEMA_signal_1269, sbox_inst_21_T1}), .clk (clk), .r (Fresh[237]), .c ({new_AGEMA_signal_1560, sbox_inst_21_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U15 ( .a ({new_AGEMA_signal_1280, sbox_inst_20_T2}), .b ({new_AGEMA_signal_1947, sbox_inst_20_n20}), .c ({output0_s1[60], output0_s0[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U14 ( .a ({new_AGEMA_signal_1765, sbox_inst_20_n19}), .b ({new_AGEMA_signal_1764, sbox_inst_20_n18}), .c ({new_AGEMA_signal_1947, sbox_inst_20_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U13 ( .a ({new_AGEMA_signal_1279, sbox_inst_20_T1}), .b ({new_AGEMA_signal_1564, sbox_inst_20_T5}), .c ({new_AGEMA_signal_1764, sbox_inst_20_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U11 ( .a ({input0_s1[81], input0_s0[81]}), .b ({new_AGEMA_signal_1766, sbox_inst_20_n16}), .c ({output0_s1[100], output0_s0[100]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U10 ( .a ({new_AGEMA_signal_1562, sbox_inst_20_n15}), .b ({new_AGEMA_signal_1564, sbox_inst_20_T5}), .c ({new_AGEMA_signal_1766, sbox_inst_20_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U9 ( .a ({new_AGEMA_signal_1562, sbox_inst_20_n15}), .b ({new_AGEMA_signal_1949, sbox_inst_20_n14}), .c ({output0_s1[140], output0_s0[140]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U8 ( .a ({new_AGEMA_signal_1561, sbox_inst_20_n13}), .b ({new_AGEMA_signal_1767, sbox_inst_20_n12}), .c ({new_AGEMA_signal_1949, sbox_inst_20_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_U7 ( .a ({new_AGEMA_signal_1565, sbox_inst_20_T6}), .b ({input0_s1[83], input0_s0[83]}), .c ({new_AGEMA_signal_1767, sbox_inst_20_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_t5_AND_U1 ( .a ({input0_s1[81], input0_s0[81]}), .b ({new_AGEMA_signal_1281, sbox_inst_20_T3}), .clk (clk), .r (Fresh[238]), .c ({new_AGEMA_signal_1564, sbox_inst_20_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_20_t6_AND_U1 ( .a ({new_AGEMA_signal_1275, sbox_inst_20_L0}), .b ({new_AGEMA_signal_1279, sbox_inst_20_T1}), .clk (clk), .r (Fresh[239]), .c ({new_AGEMA_signal_1565, sbox_inst_20_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U15 ( .a ({new_AGEMA_signal_1290, sbox_inst_19_T2}), .b ({new_AGEMA_signal_1951, sbox_inst_19_n20}), .c ({output0_s1[59], output0_s0[59]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U14 ( .a ({new_AGEMA_signal_1770, sbox_inst_19_n19}), .b ({new_AGEMA_signal_1769, sbox_inst_19_n18}), .c ({new_AGEMA_signal_1951, sbox_inst_19_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U13 ( .a ({new_AGEMA_signal_1289, sbox_inst_19_T1}), .b ({new_AGEMA_signal_1569, sbox_inst_19_T5}), .c ({new_AGEMA_signal_1769, sbox_inst_19_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U11 ( .a ({input0_s1[77], input0_s0[77]}), .b ({new_AGEMA_signal_1771, sbox_inst_19_n16}), .c ({output0_s1[99], output0_s0[99]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U10 ( .a ({new_AGEMA_signal_1567, sbox_inst_19_n15}), .b ({new_AGEMA_signal_1569, sbox_inst_19_T5}), .c ({new_AGEMA_signal_1771, sbox_inst_19_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U9 ( .a ({new_AGEMA_signal_1567, sbox_inst_19_n15}), .b ({new_AGEMA_signal_1953, sbox_inst_19_n14}), .c ({output0_s1[139], output0_s0[139]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U8 ( .a ({new_AGEMA_signal_1566, sbox_inst_19_n13}), .b ({new_AGEMA_signal_1772, sbox_inst_19_n12}), .c ({new_AGEMA_signal_1953, sbox_inst_19_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_U7 ( .a ({new_AGEMA_signal_1570, sbox_inst_19_T6}), .b ({input0_s1[79], input0_s0[79]}), .c ({new_AGEMA_signal_1772, sbox_inst_19_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_t5_AND_U1 ( .a ({input0_s1[77], input0_s0[77]}), .b ({new_AGEMA_signal_1291, sbox_inst_19_T3}), .clk (clk), .r (Fresh[240]), .c ({new_AGEMA_signal_1569, sbox_inst_19_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_19_t6_AND_U1 ( .a ({new_AGEMA_signal_1285, sbox_inst_19_L0}), .b ({new_AGEMA_signal_1289, sbox_inst_19_T1}), .clk (clk), .r (Fresh[241]), .c ({new_AGEMA_signal_1570, sbox_inst_19_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U15 ( .a ({new_AGEMA_signal_1300, sbox_inst_18_T2}), .b ({new_AGEMA_signal_1955, sbox_inst_18_n20}), .c ({output0_s1[58], output0_s0[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U14 ( .a ({new_AGEMA_signal_1775, sbox_inst_18_n19}), .b ({new_AGEMA_signal_1774, sbox_inst_18_n18}), .c ({new_AGEMA_signal_1955, sbox_inst_18_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U13 ( .a ({new_AGEMA_signal_1299, sbox_inst_18_T1}), .b ({new_AGEMA_signal_1574, sbox_inst_18_T5}), .c ({new_AGEMA_signal_1774, sbox_inst_18_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U11 ( .a ({input0_s1[73], input0_s0[73]}), .b ({new_AGEMA_signal_1776, sbox_inst_18_n16}), .c ({output0_s1[98], output0_s0[98]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U10 ( .a ({new_AGEMA_signal_1572, sbox_inst_18_n15}), .b ({new_AGEMA_signal_1574, sbox_inst_18_T5}), .c ({new_AGEMA_signal_1776, sbox_inst_18_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U9 ( .a ({new_AGEMA_signal_1572, sbox_inst_18_n15}), .b ({new_AGEMA_signal_1957, sbox_inst_18_n14}), .c ({output0_s1[138], output0_s0[138]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U8 ( .a ({new_AGEMA_signal_1571, sbox_inst_18_n13}), .b ({new_AGEMA_signal_1777, sbox_inst_18_n12}), .c ({new_AGEMA_signal_1957, sbox_inst_18_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_U7 ( .a ({new_AGEMA_signal_1575, sbox_inst_18_T6}), .b ({input0_s1[75], input0_s0[75]}), .c ({new_AGEMA_signal_1777, sbox_inst_18_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_t5_AND_U1 ( .a ({input0_s1[73], input0_s0[73]}), .b ({new_AGEMA_signal_1301, sbox_inst_18_T3}), .clk (clk), .r (Fresh[242]), .c ({new_AGEMA_signal_1574, sbox_inst_18_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_18_t6_AND_U1 ( .a ({new_AGEMA_signal_1295, sbox_inst_18_L0}), .b ({new_AGEMA_signal_1299, sbox_inst_18_T1}), .clk (clk), .r (Fresh[243]), .c ({new_AGEMA_signal_1575, sbox_inst_18_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U15 ( .a ({new_AGEMA_signal_1310, sbox_inst_17_T2}), .b ({new_AGEMA_signal_1959, sbox_inst_17_n20}), .c ({output0_s1[57], output0_s0[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U14 ( .a ({new_AGEMA_signal_1780, sbox_inst_17_n19}), .b ({new_AGEMA_signal_1779, sbox_inst_17_n18}), .c ({new_AGEMA_signal_1959, sbox_inst_17_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U13 ( .a ({new_AGEMA_signal_1309, sbox_inst_17_T1}), .b ({new_AGEMA_signal_1579, sbox_inst_17_T5}), .c ({new_AGEMA_signal_1779, sbox_inst_17_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U11 ( .a ({input0_s1[69], input0_s0[69]}), .b ({new_AGEMA_signal_1781, sbox_inst_17_n16}), .c ({output0_s1[97], output0_s0[97]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U10 ( .a ({new_AGEMA_signal_1577, sbox_inst_17_n15}), .b ({new_AGEMA_signal_1579, sbox_inst_17_T5}), .c ({new_AGEMA_signal_1781, sbox_inst_17_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U9 ( .a ({new_AGEMA_signal_1577, sbox_inst_17_n15}), .b ({new_AGEMA_signal_1961, sbox_inst_17_n14}), .c ({output0_s1[137], output0_s0[137]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U8 ( .a ({new_AGEMA_signal_1576, sbox_inst_17_n13}), .b ({new_AGEMA_signal_1782, sbox_inst_17_n12}), .c ({new_AGEMA_signal_1961, sbox_inst_17_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_U7 ( .a ({new_AGEMA_signal_1580, sbox_inst_17_T6}), .b ({input0_s1[71], input0_s0[71]}), .c ({new_AGEMA_signal_1782, sbox_inst_17_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_t5_AND_U1 ( .a ({input0_s1[69], input0_s0[69]}), .b ({new_AGEMA_signal_1311, sbox_inst_17_T3}), .clk (clk), .r (Fresh[244]), .c ({new_AGEMA_signal_1579, sbox_inst_17_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_17_t6_AND_U1 ( .a ({new_AGEMA_signal_1305, sbox_inst_17_L0}), .b ({new_AGEMA_signal_1309, sbox_inst_17_T1}), .clk (clk), .r (Fresh[245]), .c ({new_AGEMA_signal_1580, sbox_inst_17_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U15 ( .a ({new_AGEMA_signal_1320, sbox_inst_16_T2}), .b ({new_AGEMA_signal_1963, sbox_inst_16_n20}), .c ({output0_s1[56], output0_s0[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U14 ( .a ({new_AGEMA_signal_1785, sbox_inst_16_n19}), .b ({new_AGEMA_signal_1784, sbox_inst_16_n18}), .c ({new_AGEMA_signal_1963, sbox_inst_16_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U13 ( .a ({new_AGEMA_signal_1319, sbox_inst_16_T1}), .b ({new_AGEMA_signal_1584, sbox_inst_16_T5}), .c ({new_AGEMA_signal_1784, sbox_inst_16_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U11 ( .a ({input0_s1[65], input0_s0[65]}), .b ({new_AGEMA_signal_1786, sbox_inst_16_n16}), .c ({output0_s1[96], output0_s0[96]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U10 ( .a ({new_AGEMA_signal_1582, sbox_inst_16_n15}), .b ({new_AGEMA_signal_1584, sbox_inst_16_T5}), .c ({new_AGEMA_signal_1786, sbox_inst_16_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U9 ( .a ({new_AGEMA_signal_1582, sbox_inst_16_n15}), .b ({new_AGEMA_signal_1965, sbox_inst_16_n14}), .c ({output0_s1[136], output0_s0[136]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U8 ( .a ({new_AGEMA_signal_1581, sbox_inst_16_n13}), .b ({new_AGEMA_signal_1787, sbox_inst_16_n12}), .c ({new_AGEMA_signal_1965, sbox_inst_16_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_U7 ( .a ({new_AGEMA_signal_1585, sbox_inst_16_T6}), .b ({input0_s1[67], input0_s0[67]}), .c ({new_AGEMA_signal_1787, sbox_inst_16_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_t5_AND_U1 ( .a ({input0_s1[65], input0_s0[65]}), .b ({new_AGEMA_signal_1321, sbox_inst_16_T3}), .clk (clk), .r (Fresh[246]), .c ({new_AGEMA_signal_1584, sbox_inst_16_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_16_t6_AND_U1 ( .a ({new_AGEMA_signal_1315, sbox_inst_16_L0}), .b ({new_AGEMA_signal_1319, sbox_inst_16_T1}), .clk (clk), .r (Fresh[247]), .c ({new_AGEMA_signal_1585, sbox_inst_16_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U15 ( .a ({new_AGEMA_signal_1330, sbox_inst_15_T2}), .b ({new_AGEMA_signal_1967, sbox_inst_15_n20}), .c ({output0_s1[55], output0_s0[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U14 ( .a ({new_AGEMA_signal_1790, sbox_inst_15_n19}), .b ({new_AGEMA_signal_1789, sbox_inst_15_n18}), .c ({new_AGEMA_signal_1967, sbox_inst_15_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U13 ( .a ({new_AGEMA_signal_1329, sbox_inst_15_T1}), .b ({new_AGEMA_signal_1589, sbox_inst_15_T5}), .c ({new_AGEMA_signal_1789, sbox_inst_15_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U11 ( .a ({input0_s1[61], input0_s0[61]}), .b ({new_AGEMA_signal_1791, sbox_inst_15_n16}), .c ({output0_s1[95], output0_s0[95]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U10 ( .a ({new_AGEMA_signal_1587, sbox_inst_15_n15}), .b ({new_AGEMA_signal_1589, sbox_inst_15_T5}), .c ({new_AGEMA_signal_1791, sbox_inst_15_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U9 ( .a ({new_AGEMA_signal_1587, sbox_inst_15_n15}), .b ({new_AGEMA_signal_1969, sbox_inst_15_n14}), .c ({output0_s1[135], output0_s0[135]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U8 ( .a ({new_AGEMA_signal_1586, sbox_inst_15_n13}), .b ({new_AGEMA_signal_1792, sbox_inst_15_n12}), .c ({new_AGEMA_signal_1969, sbox_inst_15_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_U7 ( .a ({new_AGEMA_signal_1590, sbox_inst_15_T6}), .b ({input0_s1[63], input0_s0[63]}), .c ({new_AGEMA_signal_1792, sbox_inst_15_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_t5_AND_U1 ( .a ({input0_s1[61], input0_s0[61]}), .b ({new_AGEMA_signal_1331, sbox_inst_15_T3}), .clk (clk), .r (Fresh[248]), .c ({new_AGEMA_signal_1589, sbox_inst_15_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_15_t6_AND_U1 ( .a ({new_AGEMA_signal_1325, sbox_inst_15_L0}), .b ({new_AGEMA_signal_1329, sbox_inst_15_T1}), .clk (clk), .r (Fresh[249]), .c ({new_AGEMA_signal_1590, sbox_inst_15_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U15 ( .a ({new_AGEMA_signal_1340, sbox_inst_14_T2}), .b ({new_AGEMA_signal_1971, sbox_inst_14_n20}), .c ({output0_s1[54], output0_s0[54]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U14 ( .a ({new_AGEMA_signal_1795, sbox_inst_14_n19}), .b ({new_AGEMA_signal_1794, sbox_inst_14_n18}), .c ({new_AGEMA_signal_1971, sbox_inst_14_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U13 ( .a ({new_AGEMA_signal_1339, sbox_inst_14_T1}), .b ({new_AGEMA_signal_1594, sbox_inst_14_T5}), .c ({new_AGEMA_signal_1794, sbox_inst_14_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U11 ( .a ({input0_s1[57], input0_s0[57]}), .b ({new_AGEMA_signal_1796, sbox_inst_14_n16}), .c ({output0_s1[94], output0_s0[94]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U10 ( .a ({new_AGEMA_signal_1592, sbox_inst_14_n15}), .b ({new_AGEMA_signal_1594, sbox_inst_14_T5}), .c ({new_AGEMA_signal_1796, sbox_inst_14_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U9 ( .a ({new_AGEMA_signal_1592, sbox_inst_14_n15}), .b ({new_AGEMA_signal_1973, sbox_inst_14_n14}), .c ({output0_s1[134], output0_s0[134]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U8 ( .a ({new_AGEMA_signal_1591, sbox_inst_14_n13}), .b ({new_AGEMA_signal_1797, sbox_inst_14_n12}), .c ({new_AGEMA_signal_1973, sbox_inst_14_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_U7 ( .a ({new_AGEMA_signal_1595, sbox_inst_14_T6}), .b ({input0_s1[59], input0_s0[59]}), .c ({new_AGEMA_signal_1797, sbox_inst_14_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_t5_AND_U1 ( .a ({input0_s1[57], input0_s0[57]}), .b ({new_AGEMA_signal_1341, sbox_inst_14_T3}), .clk (clk), .r (Fresh[250]), .c ({new_AGEMA_signal_1594, sbox_inst_14_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_14_t6_AND_U1 ( .a ({new_AGEMA_signal_1335, sbox_inst_14_L0}), .b ({new_AGEMA_signal_1339, sbox_inst_14_T1}), .clk (clk), .r (Fresh[251]), .c ({new_AGEMA_signal_1595, sbox_inst_14_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U15 ( .a ({new_AGEMA_signal_1350, sbox_inst_13_T2}), .b ({new_AGEMA_signal_1975, sbox_inst_13_n20}), .c ({output0_s1[53], output0_s0[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U14 ( .a ({new_AGEMA_signal_1800, sbox_inst_13_n19}), .b ({new_AGEMA_signal_1799, sbox_inst_13_n18}), .c ({new_AGEMA_signal_1975, sbox_inst_13_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U13 ( .a ({new_AGEMA_signal_1349, sbox_inst_13_T1}), .b ({new_AGEMA_signal_1599, sbox_inst_13_T5}), .c ({new_AGEMA_signal_1799, sbox_inst_13_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U11 ( .a ({input0_s1[53], input0_s0[53]}), .b ({new_AGEMA_signal_1801, sbox_inst_13_n16}), .c ({output0_s1[93], output0_s0[93]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U10 ( .a ({new_AGEMA_signal_1597, sbox_inst_13_n15}), .b ({new_AGEMA_signal_1599, sbox_inst_13_T5}), .c ({new_AGEMA_signal_1801, sbox_inst_13_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U9 ( .a ({new_AGEMA_signal_1597, sbox_inst_13_n15}), .b ({new_AGEMA_signal_1977, sbox_inst_13_n14}), .c ({output0_s1[133], output0_s0[133]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U8 ( .a ({new_AGEMA_signal_1596, sbox_inst_13_n13}), .b ({new_AGEMA_signal_1802, sbox_inst_13_n12}), .c ({new_AGEMA_signal_1977, sbox_inst_13_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_U7 ( .a ({new_AGEMA_signal_1600, sbox_inst_13_T6}), .b ({input0_s1[55], input0_s0[55]}), .c ({new_AGEMA_signal_1802, sbox_inst_13_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_t5_AND_U1 ( .a ({input0_s1[53], input0_s0[53]}), .b ({new_AGEMA_signal_1351, sbox_inst_13_T3}), .clk (clk), .r (Fresh[252]), .c ({new_AGEMA_signal_1599, sbox_inst_13_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_13_t6_AND_U1 ( .a ({new_AGEMA_signal_1345, sbox_inst_13_L0}), .b ({new_AGEMA_signal_1349, sbox_inst_13_T1}), .clk (clk), .r (Fresh[253]), .c ({new_AGEMA_signal_1600, sbox_inst_13_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U15 ( .a ({new_AGEMA_signal_1360, sbox_inst_12_T2}), .b ({new_AGEMA_signal_1979, sbox_inst_12_n20}), .c ({output0_s1[52], output0_s0[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U14 ( .a ({new_AGEMA_signal_1805, sbox_inst_12_n19}), .b ({new_AGEMA_signal_1804, sbox_inst_12_n18}), .c ({new_AGEMA_signal_1979, sbox_inst_12_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U13 ( .a ({new_AGEMA_signal_1359, sbox_inst_12_T1}), .b ({new_AGEMA_signal_1604, sbox_inst_12_T5}), .c ({new_AGEMA_signal_1804, sbox_inst_12_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U11 ( .a ({input0_s1[49], input0_s0[49]}), .b ({new_AGEMA_signal_1806, sbox_inst_12_n16}), .c ({output0_s1[92], output0_s0[92]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U10 ( .a ({new_AGEMA_signal_1602, sbox_inst_12_n15}), .b ({new_AGEMA_signal_1604, sbox_inst_12_T5}), .c ({new_AGEMA_signal_1806, sbox_inst_12_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U9 ( .a ({new_AGEMA_signal_1602, sbox_inst_12_n15}), .b ({new_AGEMA_signal_1981, sbox_inst_12_n14}), .c ({output0_s1[132], output0_s0[132]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U8 ( .a ({new_AGEMA_signal_1601, sbox_inst_12_n13}), .b ({new_AGEMA_signal_1807, sbox_inst_12_n12}), .c ({new_AGEMA_signal_1981, sbox_inst_12_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_U7 ( .a ({new_AGEMA_signal_1605, sbox_inst_12_T6}), .b ({input0_s1[51], input0_s0[51]}), .c ({new_AGEMA_signal_1807, sbox_inst_12_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_t5_AND_U1 ( .a ({input0_s1[49], input0_s0[49]}), .b ({new_AGEMA_signal_1361, sbox_inst_12_T3}), .clk (clk), .r (Fresh[254]), .c ({new_AGEMA_signal_1604, sbox_inst_12_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_12_t6_AND_U1 ( .a ({new_AGEMA_signal_1355, sbox_inst_12_L0}), .b ({new_AGEMA_signal_1359, sbox_inst_12_T1}), .clk (clk), .r (Fresh[255]), .c ({new_AGEMA_signal_1605, sbox_inst_12_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U15 ( .a ({new_AGEMA_signal_1370, sbox_inst_11_T2}), .b ({new_AGEMA_signal_1983, sbox_inst_11_n20}), .c ({output0_s1[51], output0_s0[51]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U14 ( .a ({new_AGEMA_signal_1810, sbox_inst_11_n19}), .b ({new_AGEMA_signal_1809, sbox_inst_11_n18}), .c ({new_AGEMA_signal_1983, sbox_inst_11_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U13 ( .a ({new_AGEMA_signal_1369, sbox_inst_11_T1}), .b ({new_AGEMA_signal_1609, sbox_inst_11_T5}), .c ({new_AGEMA_signal_1809, sbox_inst_11_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U11 ( .a ({input0_s1[45], input0_s0[45]}), .b ({new_AGEMA_signal_1811, sbox_inst_11_n16}), .c ({output0_s1[91], output0_s0[91]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U10 ( .a ({new_AGEMA_signal_1607, sbox_inst_11_n15}), .b ({new_AGEMA_signal_1609, sbox_inst_11_T5}), .c ({new_AGEMA_signal_1811, sbox_inst_11_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U9 ( .a ({new_AGEMA_signal_1607, sbox_inst_11_n15}), .b ({new_AGEMA_signal_1985, sbox_inst_11_n14}), .c ({output0_s1[131], output0_s0[131]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U8 ( .a ({new_AGEMA_signal_1606, sbox_inst_11_n13}), .b ({new_AGEMA_signal_1812, sbox_inst_11_n12}), .c ({new_AGEMA_signal_1985, sbox_inst_11_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_U7 ( .a ({new_AGEMA_signal_1610, sbox_inst_11_T6}), .b ({input0_s1[47], input0_s0[47]}), .c ({new_AGEMA_signal_1812, sbox_inst_11_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_t5_AND_U1 ( .a ({input0_s1[45], input0_s0[45]}), .b ({new_AGEMA_signal_1371, sbox_inst_11_T3}), .clk (clk), .r (Fresh[256]), .c ({new_AGEMA_signal_1609, sbox_inst_11_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_11_t6_AND_U1 ( .a ({new_AGEMA_signal_1365, sbox_inst_11_L0}), .b ({new_AGEMA_signal_1369, sbox_inst_11_T1}), .clk (clk), .r (Fresh[257]), .c ({new_AGEMA_signal_1610, sbox_inst_11_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U15 ( .a ({new_AGEMA_signal_1380, sbox_inst_10_T2}), .b ({new_AGEMA_signal_1987, sbox_inst_10_n20}), .c ({output0_s1[50], output0_s0[50]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U14 ( .a ({new_AGEMA_signal_1815, sbox_inst_10_n19}), .b ({new_AGEMA_signal_1814, sbox_inst_10_n18}), .c ({new_AGEMA_signal_1987, sbox_inst_10_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U13 ( .a ({new_AGEMA_signal_1379, sbox_inst_10_T1}), .b ({new_AGEMA_signal_1614, sbox_inst_10_T5}), .c ({new_AGEMA_signal_1814, sbox_inst_10_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U11 ( .a ({input0_s1[41], input0_s0[41]}), .b ({new_AGEMA_signal_1816, sbox_inst_10_n16}), .c ({output0_s1[90], output0_s0[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U10 ( .a ({new_AGEMA_signal_1612, sbox_inst_10_n15}), .b ({new_AGEMA_signal_1614, sbox_inst_10_T5}), .c ({new_AGEMA_signal_1816, sbox_inst_10_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U9 ( .a ({new_AGEMA_signal_1612, sbox_inst_10_n15}), .b ({new_AGEMA_signal_1989, sbox_inst_10_n14}), .c ({output0_s1[130], output0_s0[130]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U8 ( .a ({new_AGEMA_signal_1611, sbox_inst_10_n13}), .b ({new_AGEMA_signal_1817, sbox_inst_10_n12}), .c ({new_AGEMA_signal_1989, sbox_inst_10_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_U7 ( .a ({new_AGEMA_signal_1615, sbox_inst_10_T6}), .b ({input0_s1[43], input0_s0[43]}), .c ({new_AGEMA_signal_1817, sbox_inst_10_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_t5_AND_U1 ( .a ({input0_s1[41], input0_s0[41]}), .b ({new_AGEMA_signal_1381, sbox_inst_10_T3}), .clk (clk), .r (Fresh[258]), .c ({new_AGEMA_signal_1614, sbox_inst_10_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_10_t6_AND_U1 ( .a ({new_AGEMA_signal_1375, sbox_inst_10_L0}), .b ({new_AGEMA_signal_1379, sbox_inst_10_T1}), .clk (clk), .r (Fresh[259]), .c ({new_AGEMA_signal_1615, sbox_inst_10_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U15 ( .a ({new_AGEMA_signal_1390, sbox_inst_9_T2}), .b ({new_AGEMA_signal_1991, sbox_inst_9_n20}), .c ({output0_s1[49], output0_s0[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U14 ( .a ({new_AGEMA_signal_1820, sbox_inst_9_n19}), .b ({new_AGEMA_signal_1819, sbox_inst_9_n18}), .c ({new_AGEMA_signal_1991, sbox_inst_9_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U13 ( .a ({new_AGEMA_signal_1389, sbox_inst_9_T1}), .b ({new_AGEMA_signal_1619, sbox_inst_9_T5}), .c ({new_AGEMA_signal_1819, sbox_inst_9_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U11 ( .a ({input0_s1[37], input0_s0[37]}), .b ({new_AGEMA_signal_1821, sbox_inst_9_n16}), .c ({output0_s1[89], output0_s0[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U10 ( .a ({new_AGEMA_signal_1617, sbox_inst_9_n15}), .b ({new_AGEMA_signal_1619, sbox_inst_9_T5}), .c ({new_AGEMA_signal_1821, sbox_inst_9_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U9 ( .a ({new_AGEMA_signal_1617, sbox_inst_9_n15}), .b ({new_AGEMA_signal_1993, sbox_inst_9_n14}), .c ({output0_s1[129], output0_s0[129]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U8 ( .a ({new_AGEMA_signal_1616, sbox_inst_9_n13}), .b ({new_AGEMA_signal_1822, sbox_inst_9_n12}), .c ({new_AGEMA_signal_1993, sbox_inst_9_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_U7 ( .a ({new_AGEMA_signal_1620, sbox_inst_9_T6}), .b ({input0_s1[39], input0_s0[39]}), .c ({new_AGEMA_signal_1822, sbox_inst_9_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_t5_AND_U1 ( .a ({input0_s1[37], input0_s0[37]}), .b ({new_AGEMA_signal_1391, sbox_inst_9_T3}), .clk (clk), .r (Fresh[260]), .c ({new_AGEMA_signal_1619, sbox_inst_9_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_9_t6_AND_U1 ( .a ({new_AGEMA_signal_1385, sbox_inst_9_L0}), .b ({new_AGEMA_signal_1389, sbox_inst_9_T1}), .clk (clk), .r (Fresh[261]), .c ({new_AGEMA_signal_1620, sbox_inst_9_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U15 ( .a ({new_AGEMA_signal_1400, sbox_inst_8_T2}), .b ({new_AGEMA_signal_1995, sbox_inst_8_n20}), .c ({output0_s1[48], output0_s0[48]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U14 ( .a ({new_AGEMA_signal_1825, sbox_inst_8_n19}), .b ({new_AGEMA_signal_1824, sbox_inst_8_n18}), .c ({new_AGEMA_signal_1995, sbox_inst_8_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U13 ( .a ({new_AGEMA_signal_1399, sbox_inst_8_T1}), .b ({new_AGEMA_signal_1624, sbox_inst_8_T5}), .c ({new_AGEMA_signal_1824, sbox_inst_8_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U11 ( .a ({input0_s1[33], input0_s0[33]}), .b ({new_AGEMA_signal_1826, sbox_inst_8_n16}), .c ({output0_s1[88], output0_s0[88]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U10 ( .a ({new_AGEMA_signal_1622, sbox_inst_8_n15}), .b ({new_AGEMA_signal_1624, sbox_inst_8_T5}), .c ({new_AGEMA_signal_1826, sbox_inst_8_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U9 ( .a ({new_AGEMA_signal_1622, sbox_inst_8_n15}), .b ({new_AGEMA_signal_1997, sbox_inst_8_n14}), .c ({output0_s1[128], output0_s0[128]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U8 ( .a ({new_AGEMA_signal_1621, sbox_inst_8_n13}), .b ({new_AGEMA_signal_1827, sbox_inst_8_n12}), .c ({new_AGEMA_signal_1997, sbox_inst_8_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_U7 ( .a ({new_AGEMA_signal_1625, sbox_inst_8_T6}), .b ({input0_s1[35], input0_s0[35]}), .c ({new_AGEMA_signal_1827, sbox_inst_8_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_t5_AND_U1 ( .a ({input0_s1[33], input0_s0[33]}), .b ({new_AGEMA_signal_1401, sbox_inst_8_T3}), .clk (clk), .r (Fresh[262]), .c ({new_AGEMA_signal_1624, sbox_inst_8_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_8_t6_AND_U1 ( .a ({new_AGEMA_signal_1395, sbox_inst_8_L0}), .b ({new_AGEMA_signal_1399, sbox_inst_8_T1}), .clk (clk), .r (Fresh[263]), .c ({new_AGEMA_signal_1625, sbox_inst_8_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U15 ( .a ({new_AGEMA_signal_1410, sbox_inst_7_T2}), .b ({new_AGEMA_signal_1999, sbox_inst_7_n20}), .c ({output0_s1[47], output0_s0[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U14 ( .a ({new_AGEMA_signal_1830, sbox_inst_7_n19}), .b ({new_AGEMA_signal_1829, sbox_inst_7_n18}), .c ({new_AGEMA_signal_1999, sbox_inst_7_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U13 ( .a ({new_AGEMA_signal_1409, sbox_inst_7_T1}), .b ({new_AGEMA_signal_1629, sbox_inst_7_T5}), .c ({new_AGEMA_signal_1829, sbox_inst_7_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U11 ( .a ({input0_s1[29], input0_s0[29]}), .b ({new_AGEMA_signal_1831, sbox_inst_7_n16}), .c ({output0_s1[87], output0_s0[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U10 ( .a ({new_AGEMA_signal_1627, sbox_inst_7_n15}), .b ({new_AGEMA_signal_1629, sbox_inst_7_T5}), .c ({new_AGEMA_signal_1831, sbox_inst_7_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U9 ( .a ({new_AGEMA_signal_1627, sbox_inst_7_n15}), .b ({new_AGEMA_signal_2001, sbox_inst_7_n14}), .c ({output0_s1[127], output0_s0[127]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U8 ( .a ({new_AGEMA_signal_1626, sbox_inst_7_n13}), .b ({new_AGEMA_signal_1832, sbox_inst_7_n12}), .c ({new_AGEMA_signal_2001, sbox_inst_7_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_U7 ( .a ({new_AGEMA_signal_1630, sbox_inst_7_T6}), .b ({input0_s1[31], input0_s0[31]}), .c ({new_AGEMA_signal_1832, sbox_inst_7_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_t5_AND_U1 ( .a ({input0_s1[29], input0_s0[29]}), .b ({new_AGEMA_signal_1411, sbox_inst_7_T3}), .clk (clk), .r (Fresh[264]), .c ({new_AGEMA_signal_1629, sbox_inst_7_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_7_t6_AND_U1 ( .a ({new_AGEMA_signal_1405, sbox_inst_7_L0}), .b ({new_AGEMA_signal_1409, sbox_inst_7_T1}), .clk (clk), .r (Fresh[265]), .c ({new_AGEMA_signal_1630, sbox_inst_7_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U15 ( .a ({new_AGEMA_signal_1420, sbox_inst_6_T2}), .b ({new_AGEMA_signal_2003, sbox_inst_6_n20}), .c ({output0_s1[46], output0_s0[46]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U14 ( .a ({new_AGEMA_signal_1835, sbox_inst_6_n19}), .b ({new_AGEMA_signal_1834, sbox_inst_6_n18}), .c ({new_AGEMA_signal_2003, sbox_inst_6_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U13 ( .a ({new_AGEMA_signal_1419, sbox_inst_6_T1}), .b ({new_AGEMA_signal_1634, sbox_inst_6_T5}), .c ({new_AGEMA_signal_1834, sbox_inst_6_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U11 ( .a ({input0_s1[25], input0_s0[25]}), .b ({new_AGEMA_signal_1836, sbox_inst_6_n16}), .c ({output0_s1[86], output0_s0[86]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U10 ( .a ({new_AGEMA_signal_1632, sbox_inst_6_n15}), .b ({new_AGEMA_signal_1634, sbox_inst_6_T5}), .c ({new_AGEMA_signal_1836, sbox_inst_6_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U9 ( .a ({new_AGEMA_signal_1632, sbox_inst_6_n15}), .b ({new_AGEMA_signal_2005, sbox_inst_6_n14}), .c ({output0_s1[126], output0_s0[126]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U8 ( .a ({new_AGEMA_signal_1631, sbox_inst_6_n13}), .b ({new_AGEMA_signal_1837, sbox_inst_6_n12}), .c ({new_AGEMA_signal_2005, sbox_inst_6_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_U7 ( .a ({new_AGEMA_signal_1635, sbox_inst_6_T6}), .b ({input0_s1[27], input0_s0[27]}), .c ({new_AGEMA_signal_1837, sbox_inst_6_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_t5_AND_U1 ( .a ({input0_s1[25], input0_s0[25]}), .b ({new_AGEMA_signal_1421, sbox_inst_6_T3}), .clk (clk), .r (Fresh[266]), .c ({new_AGEMA_signal_1634, sbox_inst_6_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_6_t6_AND_U1 ( .a ({new_AGEMA_signal_1415, sbox_inst_6_L0}), .b ({new_AGEMA_signal_1419, sbox_inst_6_T1}), .clk (clk), .r (Fresh[267]), .c ({new_AGEMA_signal_1635, sbox_inst_6_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U15 ( .a ({new_AGEMA_signal_1430, sbox_inst_5_T2}), .b ({new_AGEMA_signal_2007, sbox_inst_5_n20}), .c ({output0_s1[45], output0_s0[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U14 ( .a ({new_AGEMA_signal_1840, sbox_inst_5_n19}), .b ({new_AGEMA_signal_1839, sbox_inst_5_n18}), .c ({new_AGEMA_signal_2007, sbox_inst_5_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U13 ( .a ({new_AGEMA_signal_1429, sbox_inst_5_T1}), .b ({new_AGEMA_signal_1639, sbox_inst_5_T5}), .c ({new_AGEMA_signal_1839, sbox_inst_5_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U11 ( .a ({input0_s1[21], input0_s0[21]}), .b ({new_AGEMA_signal_1841, sbox_inst_5_n16}), .c ({output0_s1[85], output0_s0[85]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U10 ( .a ({new_AGEMA_signal_1637, sbox_inst_5_n15}), .b ({new_AGEMA_signal_1639, sbox_inst_5_T5}), .c ({new_AGEMA_signal_1841, sbox_inst_5_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U9 ( .a ({new_AGEMA_signal_1637, sbox_inst_5_n15}), .b ({new_AGEMA_signal_2009, sbox_inst_5_n14}), .c ({output0_s1[125], output0_s0[125]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U8 ( .a ({new_AGEMA_signal_1636, sbox_inst_5_n13}), .b ({new_AGEMA_signal_1842, sbox_inst_5_n12}), .c ({new_AGEMA_signal_2009, sbox_inst_5_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_U7 ( .a ({new_AGEMA_signal_1640, sbox_inst_5_T6}), .b ({input0_s1[23], input0_s0[23]}), .c ({new_AGEMA_signal_1842, sbox_inst_5_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_t5_AND_U1 ( .a ({input0_s1[21], input0_s0[21]}), .b ({new_AGEMA_signal_1431, sbox_inst_5_T3}), .clk (clk), .r (Fresh[268]), .c ({new_AGEMA_signal_1639, sbox_inst_5_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_5_t6_AND_U1 ( .a ({new_AGEMA_signal_1425, sbox_inst_5_L0}), .b ({new_AGEMA_signal_1429, sbox_inst_5_T1}), .clk (clk), .r (Fresh[269]), .c ({new_AGEMA_signal_1640, sbox_inst_5_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U15 ( .a ({new_AGEMA_signal_1440, sbox_inst_4_T2}), .b ({new_AGEMA_signal_2011, sbox_inst_4_n20}), .c ({output0_s1[44], output0_s0[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U14 ( .a ({new_AGEMA_signal_1845, sbox_inst_4_n19}), .b ({new_AGEMA_signal_1844, sbox_inst_4_n18}), .c ({new_AGEMA_signal_2011, sbox_inst_4_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U13 ( .a ({new_AGEMA_signal_1439, sbox_inst_4_T1}), .b ({new_AGEMA_signal_1644, sbox_inst_4_T5}), .c ({new_AGEMA_signal_1844, sbox_inst_4_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U11 ( .a ({input0_s1[17], input0_s0[17]}), .b ({new_AGEMA_signal_1846, sbox_inst_4_n16}), .c ({output0_s1[84], output0_s0[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U10 ( .a ({new_AGEMA_signal_1642, sbox_inst_4_n15}), .b ({new_AGEMA_signal_1644, sbox_inst_4_T5}), .c ({new_AGEMA_signal_1846, sbox_inst_4_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U9 ( .a ({new_AGEMA_signal_1642, sbox_inst_4_n15}), .b ({new_AGEMA_signal_2013, sbox_inst_4_n14}), .c ({output0_s1[124], output0_s0[124]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U8 ( .a ({new_AGEMA_signal_1641, sbox_inst_4_n13}), .b ({new_AGEMA_signal_1847, sbox_inst_4_n12}), .c ({new_AGEMA_signal_2013, sbox_inst_4_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_U7 ( .a ({new_AGEMA_signal_1645, sbox_inst_4_T6}), .b ({input0_s1[19], input0_s0[19]}), .c ({new_AGEMA_signal_1847, sbox_inst_4_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_t5_AND_U1 ( .a ({input0_s1[17], input0_s0[17]}), .b ({new_AGEMA_signal_1441, sbox_inst_4_T3}), .clk (clk), .r (Fresh[270]), .c ({new_AGEMA_signal_1644, sbox_inst_4_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_4_t6_AND_U1 ( .a ({new_AGEMA_signal_1435, sbox_inst_4_L0}), .b ({new_AGEMA_signal_1439, sbox_inst_4_T1}), .clk (clk), .r (Fresh[271]), .c ({new_AGEMA_signal_1645, sbox_inst_4_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U15 ( .a ({new_AGEMA_signal_1450, sbox_inst_3_T2}), .b ({new_AGEMA_signal_2015, sbox_inst_3_n20}), .c ({output0_s1[43], output0_s0[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U14 ( .a ({new_AGEMA_signal_1850, sbox_inst_3_n19}), .b ({new_AGEMA_signal_1849, sbox_inst_3_n18}), .c ({new_AGEMA_signal_2015, sbox_inst_3_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U13 ( .a ({new_AGEMA_signal_1449, sbox_inst_3_T1}), .b ({new_AGEMA_signal_1649, sbox_inst_3_T5}), .c ({new_AGEMA_signal_1849, sbox_inst_3_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U11 ( .a ({input0_s1[13], input0_s0[13]}), .b ({new_AGEMA_signal_1851, sbox_inst_3_n16}), .c ({output0_s1[83], output0_s0[83]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U10 ( .a ({new_AGEMA_signal_1647, sbox_inst_3_n15}), .b ({new_AGEMA_signal_1649, sbox_inst_3_T5}), .c ({new_AGEMA_signal_1851, sbox_inst_3_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U9 ( .a ({new_AGEMA_signal_1647, sbox_inst_3_n15}), .b ({new_AGEMA_signal_2017, sbox_inst_3_n14}), .c ({output0_s1[123], output0_s0[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U8 ( .a ({new_AGEMA_signal_1646, sbox_inst_3_n13}), .b ({new_AGEMA_signal_1852, sbox_inst_3_n12}), .c ({new_AGEMA_signal_2017, sbox_inst_3_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_U7 ( .a ({new_AGEMA_signal_1650, sbox_inst_3_T6}), .b ({input0_s1[15], input0_s0[15]}), .c ({new_AGEMA_signal_1852, sbox_inst_3_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_t5_AND_U1 ( .a ({input0_s1[13], input0_s0[13]}), .b ({new_AGEMA_signal_1451, sbox_inst_3_T3}), .clk (clk), .r (Fresh[272]), .c ({new_AGEMA_signal_1649, sbox_inst_3_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_3_t6_AND_U1 ( .a ({new_AGEMA_signal_1445, sbox_inst_3_L0}), .b ({new_AGEMA_signal_1449, sbox_inst_3_T1}), .clk (clk), .r (Fresh[273]), .c ({new_AGEMA_signal_1650, sbox_inst_3_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U15 ( .a ({new_AGEMA_signal_1460, sbox_inst_2_T2}), .b ({new_AGEMA_signal_2019, sbox_inst_2_n20}), .c ({output0_s1[42], output0_s0[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U14 ( .a ({new_AGEMA_signal_1855, sbox_inst_2_n19}), .b ({new_AGEMA_signal_1854, sbox_inst_2_n18}), .c ({new_AGEMA_signal_2019, sbox_inst_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U13 ( .a ({new_AGEMA_signal_1459, sbox_inst_2_T1}), .b ({new_AGEMA_signal_1654, sbox_inst_2_T5}), .c ({new_AGEMA_signal_1854, sbox_inst_2_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U11 ( .a ({input0_s1[9], input0_s0[9]}), .b ({new_AGEMA_signal_1856, sbox_inst_2_n16}), .c ({output0_s1[82], output0_s0[82]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U10 ( .a ({new_AGEMA_signal_1652, sbox_inst_2_n15}), .b ({new_AGEMA_signal_1654, sbox_inst_2_T5}), .c ({new_AGEMA_signal_1856, sbox_inst_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U9 ( .a ({new_AGEMA_signal_1652, sbox_inst_2_n15}), .b ({new_AGEMA_signal_2021, sbox_inst_2_n14}), .c ({output0_s1[122], output0_s0[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U8 ( .a ({new_AGEMA_signal_1651, sbox_inst_2_n13}), .b ({new_AGEMA_signal_1857, sbox_inst_2_n12}), .c ({new_AGEMA_signal_2021, sbox_inst_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_U7 ( .a ({new_AGEMA_signal_1655, sbox_inst_2_T6}), .b ({input0_s1[11], input0_s0[11]}), .c ({new_AGEMA_signal_1857, sbox_inst_2_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_t5_AND_U1 ( .a ({input0_s1[9], input0_s0[9]}), .b ({new_AGEMA_signal_1461, sbox_inst_2_T3}), .clk (clk), .r (Fresh[274]), .c ({new_AGEMA_signal_1654, sbox_inst_2_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_2_t6_AND_U1 ( .a ({new_AGEMA_signal_1455, sbox_inst_2_L0}), .b ({new_AGEMA_signal_1459, sbox_inst_2_T1}), .clk (clk), .r (Fresh[275]), .c ({new_AGEMA_signal_1655, sbox_inst_2_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U15 ( .a ({new_AGEMA_signal_1660, sbox_inst_1_T2}), .b ({new_AGEMA_signal_2113, sbox_inst_1_n20}), .c ({output0_s1[41], output0_s0[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U14 ( .a ({new_AGEMA_signal_2024, sbox_inst_1_n19}), .b ({new_AGEMA_signal_2023, sbox_inst_1_n18}), .c ({new_AGEMA_signal_2113, sbox_inst_1_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U13 ( .a ({new_AGEMA_signal_1659, sbox_inst_1_T1}), .b ({new_AGEMA_signal_1862, sbox_inst_1_T5}), .c ({new_AGEMA_signal_2023, sbox_inst_1_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U11 ( .a ({new_AGEMA_signal_1082, input_array_5}), .b ({new_AGEMA_signal_2025, sbox_inst_1_n16}), .c ({output0_s1[81], output0_s0[81]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U10 ( .a ({new_AGEMA_signal_1860, sbox_inst_1_n15}), .b ({new_AGEMA_signal_1862, sbox_inst_1_T5}), .c ({new_AGEMA_signal_2025, sbox_inst_1_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U9 ( .a ({new_AGEMA_signal_1860, sbox_inst_1_n15}), .b ({new_AGEMA_signal_2115, sbox_inst_1_n14}), .c ({output0_s1[121], output0_s0[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U8 ( .a ({new_AGEMA_signal_1859, sbox_inst_1_n13}), .b ({new_AGEMA_signal_2026, sbox_inst_1_n12}), .c ({new_AGEMA_signal_2115, sbox_inst_1_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_U7 ( .a ({new_AGEMA_signal_1863, sbox_inst_1_T6}), .b ({input0_s1[7], input0_s0[7]}), .c ({new_AGEMA_signal_2026, sbox_inst_1_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_t5_AND_U1 ( .a ({new_AGEMA_signal_1082, input_array_5}), .b ({new_AGEMA_signal_1661, sbox_inst_1_T3}), .clk (clk), .r (Fresh[276]), .c ({new_AGEMA_signal_1862, sbox_inst_1_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_1_t6_AND_U1 ( .a ({new_AGEMA_signal_1656, sbox_inst_1_L0}), .b ({new_AGEMA_signal_1659, sbox_inst_1_T1}), .clk (clk), .r (Fresh[277]), .c ({new_AGEMA_signal_1863, sbox_inst_1_T6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U15 ( .a ({new_AGEMA_signal_1666, sbox_inst_0_T2}), .b ({new_AGEMA_signal_2117, sbox_inst_0_n20}), .c ({output0_s1[40], output0_s0[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U14 ( .a ({new_AGEMA_signal_2029, sbox_inst_0_n19}), .b ({new_AGEMA_signal_2028, sbox_inst_0_n18}), .c ({new_AGEMA_signal_2117, sbox_inst_0_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U13 ( .a ({new_AGEMA_signal_1665, sbox_inst_0_T1}), .b ({new_AGEMA_signal_1867, sbox_inst_0_T5}), .c ({new_AGEMA_signal_2028, sbox_inst_0_n18}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U11 ( .a ({new_AGEMA_signal_1076, input_array_1}), .b ({new_AGEMA_signal_2030, sbox_inst_0_n16}), .c ({output0_s1[80], output0_s0[80]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U10 ( .a ({new_AGEMA_signal_1865, sbox_inst_0_n15}), .b ({new_AGEMA_signal_1867, sbox_inst_0_T5}), .c ({new_AGEMA_signal_2030, sbox_inst_0_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U9 ( .a ({new_AGEMA_signal_1865, sbox_inst_0_n15}), .b ({new_AGEMA_signal_2119, sbox_inst_0_n14}), .c ({output0_s1[120], output0_s0[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U8 ( .a ({new_AGEMA_signal_1864, sbox_inst_0_n13}), .b ({new_AGEMA_signal_2031, sbox_inst_0_n12}), .c ({new_AGEMA_signal_2119, sbox_inst_0_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_U7 ( .a ({new_AGEMA_signal_1868, sbox_inst_0_T6}), .b ({new_AGEMA_signal_1088, input_array_3}), .c ({new_AGEMA_signal_2031, sbox_inst_0_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_t5_AND_U1 ( .a ({new_AGEMA_signal_1076, input_array_1}), .b ({new_AGEMA_signal_1667, sbox_inst_0_T3}), .clk (clk), .r (Fresh[278]), .c ({new_AGEMA_signal_1867, sbox_inst_0_T5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) sbox_inst_0_t6_AND_U1 ( .a ({new_AGEMA_signal_1663, sbox_inst_0_L0}), .b ({new_AGEMA_signal_1665, sbox_inst_0_T1}), .clk (clk), .r (Fresh[279]), .c ({new_AGEMA_signal_1868, sbox_inst_0_T6}) ) ;
endmodule
