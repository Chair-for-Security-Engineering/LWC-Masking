/* modified netlist. Source: module Photon_256 in file /mnt/c/Users/Amir/Desktop/Papers_in_progress/LWC_Masking/PHOTON-Beetle_first_order/agema_netlist_input/Photon_256.v */
/* clock gating is added to the circuit, the latency increased 6 time(s)  */

module Photon_256_HPC2_ClockGating_d1 (w0_s0, w1_s0, temp_s0, k, p256_sel, clk, w0_s1, w1_s1, temp_s1, Fresh, y0_s0, y1_s0, temp_next_s0, temp_next_s1, y0_s1, y1_s1);
    input [127:0] w0_s0 ;
    input [127:0] w1_s0 ;
    input [127:0] temp_s0 ;
    input [3:0] k ;
    input p256_sel ;
    input clk ;
    input [127:0] w0_s1 ;
    input [127:0] w1_s1 ;
    input [127:0] temp_s1 ;
    input [1119:0] Fresh ;
    output [127:0] y0_s0 ;
    output [127:0] y1_s0 ;
    output [127:0] temp_next_s0 ;
    output [127:0] temp_next_s1 ;
    output [127:0] y0_s1 ;
    output [127:0] y1_s1 ;
    
    wire add_sub1_0_n8 ;
    wire add_sub1_0_n7 ;
    wire add_sub1_0_n6 ;
    wire add_sub1_0_n5 ;
    wire add_sub1_0_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_0_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t0 ;
    wire add_sub1_1_n8 ;
    wire add_sub1_1_n7 ;
    wire add_sub1_1_n6 ;
    wire add_sub1_1_n5 ;
    wire add_sub1_1_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_1_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t0 ;
    wire add_sub1_2_n8 ;
    wire add_sub1_2_n7 ;
    wire add_sub1_2_n6 ;
    wire add_sub1_2_n5 ;
    wire add_sub1_2_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_2_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t0 ;
    wire add_sub1_3_n8 ;
    wire add_sub1_3_n7 ;
    wire add_sub1_3_n6 ;
    wire add_sub1_3_n5 ;
    wire add_sub1_3_addc_rom_ic_out_0_ ;
    wire add_sub1_3_addc_rom_ic_out_1_ ;
    wire add_sub1_3_addc_rom_ic_out_2_ ;
    wire add_sub1_3_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_3_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t0 ;
    wire mcs1_mcs_mat1_0_n128 ;
    wire mcs1_mcs_mat1_0_n127 ;
    wire mcs1_mcs_mat1_0_n126 ;
    wire mcs1_mcs_mat1_0_n125 ;
    wire mcs1_mcs_mat1_0_n124 ;
    wire mcs1_mcs_mat1_0_n123 ;
    wire mcs1_mcs_mat1_0_n122 ;
    wire mcs1_mcs_mat1_0_n121 ;
    wire mcs1_mcs_mat1_0_n120 ;
    wire mcs1_mcs_mat1_0_n119 ;
    wire mcs1_mcs_mat1_0_n118 ;
    wire mcs1_mcs_mat1_0_n117 ;
    wire mcs1_mcs_mat1_0_n116 ;
    wire mcs1_mcs_mat1_0_n115 ;
    wire mcs1_mcs_mat1_0_n114 ;
    wire mcs1_mcs_mat1_0_n113 ;
    wire mcs1_mcs_mat1_0_n112 ;
    wire mcs1_mcs_mat1_0_n111 ;
    wire mcs1_mcs_mat1_0_n110 ;
    wire mcs1_mcs_mat1_0_n109 ;
    wire mcs1_mcs_mat1_0_n108 ;
    wire mcs1_mcs_mat1_0_n107 ;
    wire mcs1_mcs_mat1_0_n106 ;
    wire mcs1_mcs_mat1_0_n105 ;
    wire mcs1_mcs_mat1_0_n104 ;
    wire mcs1_mcs_mat1_0_n103 ;
    wire mcs1_mcs_mat1_0_n102 ;
    wire mcs1_mcs_mat1_0_n101 ;
    wire mcs1_mcs_mat1_0_n100 ;
    wire mcs1_mcs_mat1_0_n99 ;
    wire mcs1_mcs_mat1_0_n98 ;
    wire mcs1_mcs_mat1_0_n97 ;
    wire mcs1_mcs_mat1_0_n96 ;
    wire mcs1_mcs_mat1_0_n95 ;
    wire mcs1_mcs_mat1_0_n94 ;
    wire mcs1_mcs_mat1_0_n93 ;
    wire mcs1_mcs_mat1_0_n92 ;
    wire mcs1_mcs_mat1_0_n91 ;
    wire mcs1_mcs_mat1_0_n90 ;
    wire mcs1_mcs_mat1_0_n89 ;
    wire mcs1_mcs_mat1_0_n88 ;
    wire mcs1_mcs_mat1_0_n87 ;
    wire mcs1_mcs_mat1_0_n86 ;
    wire mcs1_mcs_mat1_0_n85 ;
    wire mcs1_mcs_mat1_0_n84 ;
    wire mcs1_mcs_mat1_0_n83 ;
    wire mcs1_mcs_mat1_0_n82 ;
    wire mcs1_mcs_mat1_0_n81 ;
    wire mcs1_mcs_mat1_0_n80 ;
    wire mcs1_mcs_mat1_0_n79 ;
    wire mcs1_mcs_mat1_0_n78 ;
    wire mcs1_mcs_mat1_0_n77 ;
    wire mcs1_mcs_mat1_0_n76 ;
    wire mcs1_mcs_mat1_0_n75 ;
    wire mcs1_mcs_mat1_0_n74 ;
    wire mcs1_mcs_mat1_0_n73 ;
    wire mcs1_mcs_mat1_0_n72 ;
    wire mcs1_mcs_mat1_0_n71 ;
    wire mcs1_mcs_mat1_0_n70 ;
    wire mcs1_mcs_mat1_0_n69 ;
    wire mcs1_mcs_mat1_0_n68 ;
    wire mcs1_mcs_mat1_0_n67 ;
    wire mcs1_mcs_mat1_0_n66 ;
    wire mcs1_mcs_mat1_0_n65 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_1_n128 ;
    wire mcs1_mcs_mat1_1_n127 ;
    wire mcs1_mcs_mat1_1_n126 ;
    wire mcs1_mcs_mat1_1_n125 ;
    wire mcs1_mcs_mat1_1_n124 ;
    wire mcs1_mcs_mat1_1_n123 ;
    wire mcs1_mcs_mat1_1_n122 ;
    wire mcs1_mcs_mat1_1_n121 ;
    wire mcs1_mcs_mat1_1_n120 ;
    wire mcs1_mcs_mat1_1_n119 ;
    wire mcs1_mcs_mat1_1_n118 ;
    wire mcs1_mcs_mat1_1_n117 ;
    wire mcs1_mcs_mat1_1_n116 ;
    wire mcs1_mcs_mat1_1_n115 ;
    wire mcs1_mcs_mat1_1_n114 ;
    wire mcs1_mcs_mat1_1_n113 ;
    wire mcs1_mcs_mat1_1_n112 ;
    wire mcs1_mcs_mat1_1_n111 ;
    wire mcs1_mcs_mat1_1_n110 ;
    wire mcs1_mcs_mat1_1_n109 ;
    wire mcs1_mcs_mat1_1_n108 ;
    wire mcs1_mcs_mat1_1_n107 ;
    wire mcs1_mcs_mat1_1_n106 ;
    wire mcs1_mcs_mat1_1_n105 ;
    wire mcs1_mcs_mat1_1_n104 ;
    wire mcs1_mcs_mat1_1_n103 ;
    wire mcs1_mcs_mat1_1_n102 ;
    wire mcs1_mcs_mat1_1_n101 ;
    wire mcs1_mcs_mat1_1_n100 ;
    wire mcs1_mcs_mat1_1_n99 ;
    wire mcs1_mcs_mat1_1_n98 ;
    wire mcs1_mcs_mat1_1_n97 ;
    wire mcs1_mcs_mat1_1_n96 ;
    wire mcs1_mcs_mat1_1_n95 ;
    wire mcs1_mcs_mat1_1_n94 ;
    wire mcs1_mcs_mat1_1_n93 ;
    wire mcs1_mcs_mat1_1_n92 ;
    wire mcs1_mcs_mat1_1_n91 ;
    wire mcs1_mcs_mat1_1_n90 ;
    wire mcs1_mcs_mat1_1_n89 ;
    wire mcs1_mcs_mat1_1_n88 ;
    wire mcs1_mcs_mat1_1_n87 ;
    wire mcs1_mcs_mat1_1_n86 ;
    wire mcs1_mcs_mat1_1_n85 ;
    wire mcs1_mcs_mat1_1_n84 ;
    wire mcs1_mcs_mat1_1_n83 ;
    wire mcs1_mcs_mat1_1_n82 ;
    wire mcs1_mcs_mat1_1_n81 ;
    wire mcs1_mcs_mat1_1_n80 ;
    wire mcs1_mcs_mat1_1_n79 ;
    wire mcs1_mcs_mat1_1_n78 ;
    wire mcs1_mcs_mat1_1_n77 ;
    wire mcs1_mcs_mat1_1_n76 ;
    wire mcs1_mcs_mat1_1_n75 ;
    wire mcs1_mcs_mat1_1_n74 ;
    wire mcs1_mcs_mat1_1_n73 ;
    wire mcs1_mcs_mat1_1_n72 ;
    wire mcs1_mcs_mat1_1_n71 ;
    wire mcs1_mcs_mat1_1_n70 ;
    wire mcs1_mcs_mat1_1_n69 ;
    wire mcs1_mcs_mat1_1_n68 ;
    wire mcs1_mcs_mat1_1_n67 ;
    wire mcs1_mcs_mat1_1_n66 ;
    wire mcs1_mcs_mat1_1_n65 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_2_n128 ;
    wire mcs1_mcs_mat1_2_n127 ;
    wire mcs1_mcs_mat1_2_n126 ;
    wire mcs1_mcs_mat1_2_n125 ;
    wire mcs1_mcs_mat1_2_n124 ;
    wire mcs1_mcs_mat1_2_n123 ;
    wire mcs1_mcs_mat1_2_n122 ;
    wire mcs1_mcs_mat1_2_n121 ;
    wire mcs1_mcs_mat1_2_n120 ;
    wire mcs1_mcs_mat1_2_n119 ;
    wire mcs1_mcs_mat1_2_n118 ;
    wire mcs1_mcs_mat1_2_n117 ;
    wire mcs1_mcs_mat1_2_n116 ;
    wire mcs1_mcs_mat1_2_n115 ;
    wire mcs1_mcs_mat1_2_n114 ;
    wire mcs1_mcs_mat1_2_n113 ;
    wire mcs1_mcs_mat1_2_n112 ;
    wire mcs1_mcs_mat1_2_n111 ;
    wire mcs1_mcs_mat1_2_n110 ;
    wire mcs1_mcs_mat1_2_n109 ;
    wire mcs1_mcs_mat1_2_n108 ;
    wire mcs1_mcs_mat1_2_n107 ;
    wire mcs1_mcs_mat1_2_n106 ;
    wire mcs1_mcs_mat1_2_n105 ;
    wire mcs1_mcs_mat1_2_n104 ;
    wire mcs1_mcs_mat1_2_n103 ;
    wire mcs1_mcs_mat1_2_n102 ;
    wire mcs1_mcs_mat1_2_n101 ;
    wire mcs1_mcs_mat1_2_n100 ;
    wire mcs1_mcs_mat1_2_n99 ;
    wire mcs1_mcs_mat1_2_n98 ;
    wire mcs1_mcs_mat1_2_n97 ;
    wire mcs1_mcs_mat1_2_n96 ;
    wire mcs1_mcs_mat1_2_n95 ;
    wire mcs1_mcs_mat1_2_n94 ;
    wire mcs1_mcs_mat1_2_n93 ;
    wire mcs1_mcs_mat1_2_n92 ;
    wire mcs1_mcs_mat1_2_n91 ;
    wire mcs1_mcs_mat1_2_n90 ;
    wire mcs1_mcs_mat1_2_n89 ;
    wire mcs1_mcs_mat1_2_n88 ;
    wire mcs1_mcs_mat1_2_n87 ;
    wire mcs1_mcs_mat1_2_n86 ;
    wire mcs1_mcs_mat1_2_n85 ;
    wire mcs1_mcs_mat1_2_n84 ;
    wire mcs1_mcs_mat1_2_n83 ;
    wire mcs1_mcs_mat1_2_n82 ;
    wire mcs1_mcs_mat1_2_n81 ;
    wire mcs1_mcs_mat1_2_n80 ;
    wire mcs1_mcs_mat1_2_n79 ;
    wire mcs1_mcs_mat1_2_n78 ;
    wire mcs1_mcs_mat1_2_n77 ;
    wire mcs1_mcs_mat1_2_n76 ;
    wire mcs1_mcs_mat1_2_n75 ;
    wire mcs1_mcs_mat1_2_n74 ;
    wire mcs1_mcs_mat1_2_n73 ;
    wire mcs1_mcs_mat1_2_n72 ;
    wire mcs1_mcs_mat1_2_n71 ;
    wire mcs1_mcs_mat1_2_n70 ;
    wire mcs1_mcs_mat1_2_n69 ;
    wire mcs1_mcs_mat1_2_n68 ;
    wire mcs1_mcs_mat1_2_n67 ;
    wire mcs1_mcs_mat1_2_n66 ;
    wire mcs1_mcs_mat1_2_n65 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_3_n128 ;
    wire mcs1_mcs_mat1_3_n127 ;
    wire mcs1_mcs_mat1_3_n126 ;
    wire mcs1_mcs_mat1_3_n125 ;
    wire mcs1_mcs_mat1_3_n124 ;
    wire mcs1_mcs_mat1_3_n123 ;
    wire mcs1_mcs_mat1_3_n122 ;
    wire mcs1_mcs_mat1_3_n121 ;
    wire mcs1_mcs_mat1_3_n120 ;
    wire mcs1_mcs_mat1_3_n119 ;
    wire mcs1_mcs_mat1_3_n118 ;
    wire mcs1_mcs_mat1_3_n117 ;
    wire mcs1_mcs_mat1_3_n116 ;
    wire mcs1_mcs_mat1_3_n115 ;
    wire mcs1_mcs_mat1_3_n114 ;
    wire mcs1_mcs_mat1_3_n113 ;
    wire mcs1_mcs_mat1_3_n112 ;
    wire mcs1_mcs_mat1_3_n111 ;
    wire mcs1_mcs_mat1_3_n110 ;
    wire mcs1_mcs_mat1_3_n109 ;
    wire mcs1_mcs_mat1_3_n108 ;
    wire mcs1_mcs_mat1_3_n107 ;
    wire mcs1_mcs_mat1_3_n106 ;
    wire mcs1_mcs_mat1_3_n105 ;
    wire mcs1_mcs_mat1_3_n104 ;
    wire mcs1_mcs_mat1_3_n103 ;
    wire mcs1_mcs_mat1_3_n102 ;
    wire mcs1_mcs_mat1_3_n101 ;
    wire mcs1_mcs_mat1_3_n100 ;
    wire mcs1_mcs_mat1_3_n99 ;
    wire mcs1_mcs_mat1_3_n98 ;
    wire mcs1_mcs_mat1_3_n97 ;
    wire mcs1_mcs_mat1_3_n96 ;
    wire mcs1_mcs_mat1_3_n95 ;
    wire mcs1_mcs_mat1_3_n94 ;
    wire mcs1_mcs_mat1_3_n93 ;
    wire mcs1_mcs_mat1_3_n92 ;
    wire mcs1_mcs_mat1_3_n91 ;
    wire mcs1_mcs_mat1_3_n90 ;
    wire mcs1_mcs_mat1_3_n89 ;
    wire mcs1_mcs_mat1_3_n88 ;
    wire mcs1_mcs_mat1_3_n87 ;
    wire mcs1_mcs_mat1_3_n86 ;
    wire mcs1_mcs_mat1_3_n85 ;
    wire mcs1_mcs_mat1_3_n84 ;
    wire mcs1_mcs_mat1_3_n83 ;
    wire mcs1_mcs_mat1_3_n82 ;
    wire mcs1_mcs_mat1_3_n81 ;
    wire mcs1_mcs_mat1_3_n80 ;
    wire mcs1_mcs_mat1_3_n79 ;
    wire mcs1_mcs_mat1_3_n78 ;
    wire mcs1_mcs_mat1_3_n77 ;
    wire mcs1_mcs_mat1_3_n76 ;
    wire mcs1_mcs_mat1_3_n75 ;
    wire mcs1_mcs_mat1_3_n74 ;
    wire mcs1_mcs_mat1_3_n73 ;
    wire mcs1_mcs_mat1_3_n72 ;
    wire mcs1_mcs_mat1_3_n71 ;
    wire mcs1_mcs_mat1_3_n70 ;
    wire mcs1_mcs_mat1_3_n69 ;
    wire mcs1_mcs_mat1_3_n68 ;
    wire mcs1_mcs_mat1_3_n67 ;
    wire mcs1_mcs_mat1_3_n66 ;
    wire mcs1_mcs_mat1_3_n65 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_4_n128 ;
    wire mcs1_mcs_mat1_4_n127 ;
    wire mcs1_mcs_mat1_4_n126 ;
    wire mcs1_mcs_mat1_4_n125 ;
    wire mcs1_mcs_mat1_4_n124 ;
    wire mcs1_mcs_mat1_4_n123 ;
    wire mcs1_mcs_mat1_4_n122 ;
    wire mcs1_mcs_mat1_4_n121 ;
    wire mcs1_mcs_mat1_4_n120 ;
    wire mcs1_mcs_mat1_4_n119 ;
    wire mcs1_mcs_mat1_4_n118 ;
    wire mcs1_mcs_mat1_4_n117 ;
    wire mcs1_mcs_mat1_4_n116 ;
    wire mcs1_mcs_mat1_4_n115 ;
    wire mcs1_mcs_mat1_4_n114 ;
    wire mcs1_mcs_mat1_4_n113 ;
    wire mcs1_mcs_mat1_4_n112 ;
    wire mcs1_mcs_mat1_4_n111 ;
    wire mcs1_mcs_mat1_4_n110 ;
    wire mcs1_mcs_mat1_4_n109 ;
    wire mcs1_mcs_mat1_4_n108 ;
    wire mcs1_mcs_mat1_4_n107 ;
    wire mcs1_mcs_mat1_4_n106 ;
    wire mcs1_mcs_mat1_4_n105 ;
    wire mcs1_mcs_mat1_4_n104 ;
    wire mcs1_mcs_mat1_4_n103 ;
    wire mcs1_mcs_mat1_4_n102 ;
    wire mcs1_mcs_mat1_4_n101 ;
    wire mcs1_mcs_mat1_4_n100 ;
    wire mcs1_mcs_mat1_4_n99 ;
    wire mcs1_mcs_mat1_4_n98 ;
    wire mcs1_mcs_mat1_4_n97 ;
    wire mcs1_mcs_mat1_4_n96 ;
    wire mcs1_mcs_mat1_4_n95 ;
    wire mcs1_mcs_mat1_4_n94 ;
    wire mcs1_mcs_mat1_4_n93 ;
    wire mcs1_mcs_mat1_4_n92 ;
    wire mcs1_mcs_mat1_4_n91 ;
    wire mcs1_mcs_mat1_4_n90 ;
    wire mcs1_mcs_mat1_4_n89 ;
    wire mcs1_mcs_mat1_4_n88 ;
    wire mcs1_mcs_mat1_4_n87 ;
    wire mcs1_mcs_mat1_4_n86 ;
    wire mcs1_mcs_mat1_4_n85 ;
    wire mcs1_mcs_mat1_4_n84 ;
    wire mcs1_mcs_mat1_4_n83 ;
    wire mcs1_mcs_mat1_4_n82 ;
    wire mcs1_mcs_mat1_4_n81 ;
    wire mcs1_mcs_mat1_4_n80 ;
    wire mcs1_mcs_mat1_4_n79 ;
    wire mcs1_mcs_mat1_4_n78 ;
    wire mcs1_mcs_mat1_4_n77 ;
    wire mcs1_mcs_mat1_4_n76 ;
    wire mcs1_mcs_mat1_4_n75 ;
    wire mcs1_mcs_mat1_4_n74 ;
    wire mcs1_mcs_mat1_4_n73 ;
    wire mcs1_mcs_mat1_4_n72 ;
    wire mcs1_mcs_mat1_4_n71 ;
    wire mcs1_mcs_mat1_4_n70 ;
    wire mcs1_mcs_mat1_4_n69 ;
    wire mcs1_mcs_mat1_4_n68 ;
    wire mcs1_mcs_mat1_4_n67 ;
    wire mcs1_mcs_mat1_4_n66 ;
    wire mcs1_mcs_mat1_4_n65 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_5_n128 ;
    wire mcs1_mcs_mat1_5_n127 ;
    wire mcs1_mcs_mat1_5_n126 ;
    wire mcs1_mcs_mat1_5_n125 ;
    wire mcs1_mcs_mat1_5_n124 ;
    wire mcs1_mcs_mat1_5_n123 ;
    wire mcs1_mcs_mat1_5_n122 ;
    wire mcs1_mcs_mat1_5_n121 ;
    wire mcs1_mcs_mat1_5_n120 ;
    wire mcs1_mcs_mat1_5_n119 ;
    wire mcs1_mcs_mat1_5_n118 ;
    wire mcs1_mcs_mat1_5_n117 ;
    wire mcs1_mcs_mat1_5_n116 ;
    wire mcs1_mcs_mat1_5_n115 ;
    wire mcs1_mcs_mat1_5_n114 ;
    wire mcs1_mcs_mat1_5_n113 ;
    wire mcs1_mcs_mat1_5_n112 ;
    wire mcs1_mcs_mat1_5_n111 ;
    wire mcs1_mcs_mat1_5_n110 ;
    wire mcs1_mcs_mat1_5_n109 ;
    wire mcs1_mcs_mat1_5_n108 ;
    wire mcs1_mcs_mat1_5_n107 ;
    wire mcs1_mcs_mat1_5_n106 ;
    wire mcs1_mcs_mat1_5_n105 ;
    wire mcs1_mcs_mat1_5_n104 ;
    wire mcs1_mcs_mat1_5_n103 ;
    wire mcs1_mcs_mat1_5_n102 ;
    wire mcs1_mcs_mat1_5_n101 ;
    wire mcs1_mcs_mat1_5_n100 ;
    wire mcs1_mcs_mat1_5_n99 ;
    wire mcs1_mcs_mat1_5_n98 ;
    wire mcs1_mcs_mat1_5_n97 ;
    wire mcs1_mcs_mat1_5_n96 ;
    wire mcs1_mcs_mat1_5_n95 ;
    wire mcs1_mcs_mat1_5_n94 ;
    wire mcs1_mcs_mat1_5_n93 ;
    wire mcs1_mcs_mat1_5_n92 ;
    wire mcs1_mcs_mat1_5_n91 ;
    wire mcs1_mcs_mat1_5_n90 ;
    wire mcs1_mcs_mat1_5_n89 ;
    wire mcs1_mcs_mat1_5_n88 ;
    wire mcs1_mcs_mat1_5_n87 ;
    wire mcs1_mcs_mat1_5_n86 ;
    wire mcs1_mcs_mat1_5_n85 ;
    wire mcs1_mcs_mat1_5_n84 ;
    wire mcs1_mcs_mat1_5_n83 ;
    wire mcs1_mcs_mat1_5_n82 ;
    wire mcs1_mcs_mat1_5_n81 ;
    wire mcs1_mcs_mat1_5_n80 ;
    wire mcs1_mcs_mat1_5_n79 ;
    wire mcs1_mcs_mat1_5_n78 ;
    wire mcs1_mcs_mat1_5_n77 ;
    wire mcs1_mcs_mat1_5_n76 ;
    wire mcs1_mcs_mat1_5_n75 ;
    wire mcs1_mcs_mat1_5_n74 ;
    wire mcs1_mcs_mat1_5_n73 ;
    wire mcs1_mcs_mat1_5_n72 ;
    wire mcs1_mcs_mat1_5_n71 ;
    wire mcs1_mcs_mat1_5_n70 ;
    wire mcs1_mcs_mat1_5_n69 ;
    wire mcs1_mcs_mat1_5_n68 ;
    wire mcs1_mcs_mat1_5_n67 ;
    wire mcs1_mcs_mat1_5_n66 ;
    wire mcs1_mcs_mat1_5_n65 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_6_n128 ;
    wire mcs1_mcs_mat1_6_n127 ;
    wire mcs1_mcs_mat1_6_n126 ;
    wire mcs1_mcs_mat1_6_n125 ;
    wire mcs1_mcs_mat1_6_n124 ;
    wire mcs1_mcs_mat1_6_n123 ;
    wire mcs1_mcs_mat1_6_n122 ;
    wire mcs1_mcs_mat1_6_n121 ;
    wire mcs1_mcs_mat1_6_n120 ;
    wire mcs1_mcs_mat1_6_n119 ;
    wire mcs1_mcs_mat1_6_n118 ;
    wire mcs1_mcs_mat1_6_n117 ;
    wire mcs1_mcs_mat1_6_n116 ;
    wire mcs1_mcs_mat1_6_n115 ;
    wire mcs1_mcs_mat1_6_n114 ;
    wire mcs1_mcs_mat1_6_n113 ;
    wire mcs1_mcs_mat1_6_n112 ;
    wire mcs1_mcs_mat1_6_n111 ;
    wire mcs1_mcs_mat1_6_n110 ;
    wire mcs1_mcs_mat1_6_n109 ;
    wire mcs1_mcs_mat1_6_n108 ;
    wire mcs1_mcs_mat1_6_n107 ;
    wire mcs1_mcs_mat1_6_n106 ;
    wire mcs1_mcs_mat1_6_n105 ;
    wire mcs1_mcs_mat1_6_n104 ;
    wire mcs1_mcs_mat1_6_n103 ;
    wire mcs1_mcs_mat1_6_n102 ;
    wire mcs1_mcs_mat1_6_n101 ;
    wire mcs1_mcs_mat1_6_n100 ;
    wire mcs1_mcs_mat1_6_n99 ;
    wire mcs1_mcs_mat1_6_n98 ;
    wire mcs1_mcs_mat1_6_n97 ;
    wire mcs1_mcs_mat1_6_n96 ;
    wire mcs1_mcs_mat1_6_n95 ;
    wire mcs1_mcs_mat1_6_n94 ;
    wire mcs1_mcs_mat1_6_n93 ;
    wire mcs1_mcs_mat1_6_n92 ;
    wire mcs1_mcs_mat1_6_n91 ;
    wire mcs1_mcs_mat1_6_n90 ;
    wire mcs1_mcs_mat1_6_n89 ;
    wire mcs1_mcs_mat1_6_n88 ;
    wire mcs1_mcs_mat1_6_n87 ;
    wire mcs1_mcs_mat1_6_n86 ;
    wire mcs1_mcs_mat1_6_n85 ;
    wire mcs1_mcs_mat1_6_n84 ;
    wire mcs1_mcs_mat1_6_n83 ;
    wire mcs1_mcs_mat1_6_n82 ;
    wire mcs1_mcs_mat1_6_n81 ;
    wire mcs1_mcs_mat1_6_n80 ;
    wire mcs1_mcs_mat1_6_n79 ;
    wire mcs1_mcs_mat1_6_n78 ;
    wire mcs1_mcs_mat1_6_n77 ;
    wire mcs1_mcs_mat1_6_n76 ;
    wire mcs1_mcs_mat1_6_n75 ;
    wire mcs1_mcs_mat1_6_n74 ;
    wire mcs1_mcs_mat1_6_n73 ;
    wire mcs1_mcs_mat1_6_n72 ;
    wire mcs1_mcs_mat1_6_n71 ;
    wire mcs1_mcs_mat1_6_n70 ;
    wire mcs1_mcs_mat1_6_n69 ;
    wire mcs1_mcs_mat1_6_n68 ;
    wire mcs1_mcs_mat1_6_n67 ;
    wire mcs1_mcs_mat1_6_n66 ;
    wire mcs1_mcs_mat1_6_n65 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_7_n128 ;
    wire mcs1_mcs_mat1_7_n127 ;
    wire mcs1_mcs_mat1_7_n126 ;
    wire mcs1_mcs_mat1_7_n125 ;
    wire mcs1_mcs_mat1_7_n124 ;
    wire mcs1_mcs_mat1_7_n123 ;
    wire mcs1_mcs_mat1_7_n122 ;
    wire mcs1_mcs_mat1_7_n121 ;
    wire mcs1_mcs_mat1_7_n120 ;
    wire mcs1_mcs_mat1_7_n119 ;
    wire mcs1_mcs_mat1_7_n118 ;
    wire mcs1_mcs_mat1_7_n117 ;
    wire mcs1_mcs_mat1_7_n116 ;
    wire mcs1_mcs_mat1_7_n115 ;
    wire mcs1_mcs_mat1_7_n114 ;
    wire mcs1_mcs_mat1_7_n113 ;
    wire mcs1_mcs_mat1_7_n112 ;
    wire mcs1_mcs_mat1_7_n111 ;
    wire mcs1_mcs_mat1_7_n110 ;
    wire mcs1_mcs_mat1_7_n109 ;
    wire mcs1_mcs_mat1_7_n108 ;
    wire mcs1_mcs_mat1_7_n107 ;
    wire mcs1_mcs_mat1_7_n106 ;
    wire mcs1_mcs_mat1_7_n105 ;
    wire mcs1_mcs_mat1_7_n104 ;
    wire mcs1_mcs_mat1_7_n103 ;
    wire mcs1_mcs_mat1_7_n102 ;
    wire mcs1_mcs_mat1_7_n101 ;
    wire mcs1_mcs_mat1_7_n100 ;
    wire mcs1_mcs_mat1_7_n99 ;
    wire mcs1_mcs_mat1_7_n98 ;
    wire mcs1_mcs_mat1_7_n97 ;
    wire mcs1_mcs_mat1_7_n96 ;
    wire mcs1_mcs_mat1_7_n95 ;
    wire mcs1_mcs_mat1_7_n94 ;
    wire mcs1_mcs_mat1_7_n93 ;
    wire mcs1_mcs_mat1_7_n92 ;
    wire mcs1_mcs_mat1_7_n91 ;
    wire mcs1_mcs_mat1_7_n90 ;
    wire mcs1_mcs_mat1_7_n89 ;
    wire mcs1_mcs_mat1_7_n88 ;
    wire mcs1_mcs_mat1_7_n87 ;
    wire mcs1_mcs_mat1_7_n86 ;
    wire mcs1_mcs_mat1_7_n85 ;
    wire mcs1_mcs_mat1_7_n84 ;
    wire mcs1_mcs_mat1_7_n83 ;
    wire mcs1_mcs_mat1_7_n82 ;
    wire mcs1_mcs_mat1_7_n81 ;
    wire mcs1_mcs_mat1_7_n80 ;
    wire mcs1_mcs_mat1_7_n79 ;
    wire mcs1_mcs_mat1_7_n78 ;
    wire mcs1_mcs_mat1_7_n77 ;
    wire mcs1_mcs_mat1_7_n76 ;
    wire mcs1_mcs_mat1_7_n75 ;
    wire mcs1_mcs_mat1_7_n74 ;
    wire mcs1_mcs_mat1_7_n73 ;
    wire mcs1_mcs_mat1_7_n72 ;
    wire mcs1_mcs_mat1_7_n71 ;
    wire mcs1_mcs_mat1_7_n70 ;
    wire mcs1_mcs_mat1_7_n69 ;
    wire mcs1_mcs_mat1_7_n68 ;
    wire mcs1_mcs_mat1_7_n67 ;
    wire mcs1_mcs_mat1_7_n66 ;
    wire mcs1_mcs_mat1_7_n65 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x0x4 ;
    wire [127:0] addc_in ;
    wire [127:0] subc_out ;
    wire [124:1] shiftr_out ;
    wire [255:128] mcs_out ;
    wire [127:0] y0_1 ;
    wire [3:0] add_sub1_0_addc_out ;
    wire [2:0] add_sub1_0_addc_rom_ic_out ;
    wire [3:0] add_sub1_0_addc_rom_rc_out ;
    wire [3:0] add_sub1_1_addc_out ;
    wire [2:0] add_sub1_1_addc_rom_ic_out ;
    wire [3:0] add_sub1_1_addc_rom_rc_out ;
    wire [3:0] add_sub1_2_addc_out ;
    wire [2:0] add_sub1_2_addc_rom_ic_out ;
    wire [3:0] add_sub1_2_addc_rom_rc_out ;
    wire [3:0] add_sub1_3_addc_out ;
    wire [3:0] add_sub1_3_addc_rom_rc_out ;
    wire [127:0] mcs1_mcs_mat1_0_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_1_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_2_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_3_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_4_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_5_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_6_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_7_mcs_out ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10778 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;

    /* cells in depth 0 */
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_0_U1 ( .s (p256_sel), .b ({w0_s1[0], w0_s0[0]}), .a ({w1_s1[0], w1_s0[0]}), .c ({new_AGEMA_signal_5734, addc_in[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_1_U1 ( .s (p256_sel), .b ({w0_s1[1], w0_s0[1]}), .a ({w1_s1[1], w1_s0[1]}), .c ({new_AGEMA_signal_5737, addc_in[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_2_U1 ( .s (p256_sel), .b ({w0_s1[2], w0_s0[2]}), .a ({w1_s1[2], w1_s0[2]}), .c ({new_AGEMA_signal_5740, addc_in[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_3_U1 ( .s (p256_sel), .b ({w0_s1[3], w0_s0[3]}), .a ({w1_s1[3], w1_s0[3]}), .c ({new_AGEMA_signal_5743, addc_in[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_4_U1 ( .s (p256_sel), .b ({w0_s1[4], w0_s0[4]}), .a ({w1_s1[4], w1_s0[4]}), .c ({new_AGEMA_signal_5746, addc_in[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_5_U1 ( .s (p256_sel), .b ({w0_s1[5], w0_s0[5]}), .a ({w1_s1[5], w1_s0[5]}), .c ({new_AGEMA_signal_5749, addc_in[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_6_U1 ( .s (p256_sel), .b ({w0_s1[6], w0_s0[6]}), .a ({w1_s1[6], w1_s0[6]}), .c ({new_AGEMA_signal_5752, addc_in[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_7_U1 ( .s (p256_sel), .b ({w0_s1[7], w0_s0[7]}), .a ({w1_s1[7], w1_s0[7]}), .c ({new_AGEMA_signal_5755, addc_in[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_8_U1 ( .s (p256_sel), .b ({w0_s1[8], w0_s0[8]}), .a ({w1_s1[8], w1_s0[8]}), .c ({new_AGEMA_signal_5758, addc_in[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_9_U1 ( .s (p256_sel), .b ({w0_s1[9], w0_s0[9]}), .a ({w1_s1[9], w1_s0[9]}), .c ({new_AGEMA_signal_5761, addc_in[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_10_U1 ( .s (p256_sel), .b ({w0_s1[10], w0_s0[10]}), .a ({w1_s1[10], w1_s0[10]}), .c ({new_AGEMA_signal_5764, addc_in[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_11_U1 ( .s (p256_sel), .b ({w0_s1[11], w0_s0[11]}), .a ({w1_s1[11], w1_s0[11]}), .c ({new_AGEMA_signal_5767, addc_in[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_12_U1 ( .s (p256_sel), .b ({w0_s1[12], w0_s0[12]}), .a ({w1_s1[12], w1_s0[12]}), .c ({new_AGEMA_signal_5770, addc_in[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_13_U1 ( .s (p256_sel), .b ({w0_s1[13], w0_s0[13]}), .a ({w1_s1[13], w1_s0[13]}), .c ({new_AGEMA_signal_5773, addc_in[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_14_U1 ( .s (p256_sel), .b ({w0_s1[14], w0_s0[14]}), .a ({w1_s1[14], w1_s0[14]}), .c ({new_AGEMA_signal_5776, addc_in[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_15_U1 ( .s (p256_sel), .b ({w0_s1[15], w0_s0[15]}), .a ({w1_s1[15], w1_s0[15]}), .c ({new_AGEMA_signal_5779, addc_in[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_16_U1 ( .s (p256_sel), .b ({w0_s1[16], w0_s0[16]}), .a ({w1_s1[16], w1_s0[16]}), .c ({new_AGEMA_signal_5782, addc_in[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_17_U1 ( .s (p256_sel), .b ({w0_s1[17], w0_s0[17]}), .a ({w1_s1[17], w1_s0[17]}), .c ({new_AGEMA_signal_5785, addc_in[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_18_U1 ( .s (p256_sel), .b ({w0_s1[18], w0_s0[18]}), .a ({w1_s1[18], w1_s0[18]}), .c ({new_AGEMA_signal_5788, addc_in[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_19_U1 ( .s (p256_sel), .b ({w0_s1[19], w0_s0[19]}), .a ({w1_s1[19], w1_s0[19]}), .c ({new_AGEMA_signal_5791, addc_in[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_20_U1 ( .s (p256_sel), .b ({w0_s1[20], w0_s0[20]}), .a ({w1_s1[20], w1_s0[20]}), .c ({new_AGEMA_signal_5794, addc_in[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_21_U1 ( .s (p256_sel), .b ({w0_s1[21], w0_s0[21]}), .a ({w1_s1[21], w1_s0[21]}), .c ({new_AGEMA_signal_5797, addc_in[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_22_U1 ( .s (p256_sel), .b ({w0_s1[22], w0_s0[22]}), .a ({w1_s1[22], w1_s0[22]}), .c ({new_AGEMA_signal_5800, addc_in[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_23_U1 ( .s (p256_sel), .b ({w0_s1[23], w0_s0[23]}), .a ({w1_s1[23], w1_s0[23]}), .c ({new_AGEMA_signal_5803, addc_in[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_24_U1 ( .s (p256_sel), .b ({w0_s1[24], w0_s0[24]}), .a ({w1_s1[24], w1_s0[24]}), .c ({new_AGEMA_signal_5806, addc_in[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_25_U1 ( .s (p256_sel), .b ({w0_s1[25], w0_s0[25]}), .a ({w1_s1[25], w1_s0[25]}), .c ({new_AGEMA_signal_5809, addc_in[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_26_U1 ( .s (p256_sel), .b ({w0_s1[26], w0_s0[26]}), .a ({w1_s1[26], w1_s0[26]}), .c ({new_AGEMA_signal_5812, addc_in[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_27_U1 ( .s (p256_sel), .b ({w0_s1[27], w0_s0[27]}), .a ({w1_s1[27], w1_s0[27]}), .c ({new_AGEMA_signal_5815, addc_in[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_28_U1 ( .s (p256_sel), .b ({w0_s1[28], w0_s0[28]}), .a ({w1_s1[28], w1_s0[28]}), .c ({new_AGEMA_signal_5818, addc_in[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_29_U1 ( .s (p256_sel), .b ({w0_s1[29], w0_s0[29]}), .a ({w1_s1[29], w1_s0[29]}), .c ({new_AGEMA_signal_5821, addc_in[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_30_U1 ( .s (p256_sel), .b ({w0_s1[30], w0_s0[30]}), .a ({w1_s1[30], w1_s0[30]}), .c ({new_AGEMA_signal_5824, addc_in[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_31_U1 ( .s (p256_sel), .b ({w0_s1[31], w0_s0[31]}), .a ({w1_s1[31], w1_s0[31]}), .c ({new_AGEMA_signal_5827, addc_in[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_32_U1 ( .s (p256_sel), .b ({w0_s1[32], w0_s0[32]}), .a ({w1_s1[32], w1_s0[32]}), .c ({new_AGEMA_signal_5830, addc_in[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_33_U1 ( .s (p256_sel), .b ({w0_s1[33], w0_s0[33]}), .a ({w1_s1[33], w1_s0[33]}), .c ({new_AGEMA_signal_5833, addc_in[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_34_U1 ( .s (p256_sel), .b ({w0_s1[34], w0_s0[34]}), .a ({w1_s1[34], w1_s0[34]}), .c ({new_AGEMA_signal_5836, addc_in[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_35_U1 ( .s (p256_sel), .b ({w0_s1[35], w0_s0[35]}), .a ({w1_s1[35], w1_s0[35]}), .c ({new_AGEMA_signal_5839, addc_in[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_36_U1 ( .s (p256_sel), .b ({w0_s1[36], w0_s0[36]}), .a ({w1_s1[36], w1_s0[36]}), .c ({new_AGEMA_signal_5842, addc_in[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_37_U1 ( .s (p256_sel), .b ({w0_s1[37], w0_s0[37]}), .a ({w1_s1[37], w1_s0[37]}), .c ({new_AGEMA_signal_5845, addc_in[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_38_U1 ( .s (p256_sel), .b ({w0_s1[38], w0_s0[38]}), .a ({w1_s1[38], w1_s0[38]}), .c ({new_AGEMA_signal_5848, addc_in[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_39_U1 ( .s (p256_sel), .b ({w0_s1[39], w0_s0[39]}), .a ({w1_s1[39], w1_s0[39]}), .c ({new_AGEMA_signal_5851, addc_in[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_40_U1 ( .s (p256_sel), .b ({w0_s1[40], w0_s0[40]}), .a ({w1_s1[40], w1_s0[40]}), .c ({new_AGEMA_signal_5854, addc_in[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_41_U1 ( .s (p256_sel), .b ({w0_s1[41], w0_s0[41]}), .a ({w1_s1[41], w1_s0[41]}), .c ({new_AGEMA_signal_5857, addc_in[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_42_U1 ( .s (p256_sel), .b ({w0_s1[42], w0_s0[42]}), .a ({w1_s1[42], w1_s0[42]}), .c ({new_AGEMA_signal_5860, addc_in[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_43_U1 ( .s (p256_sel), .b ({w0_s1[43], w0_s0[43]}), .a ({w1_s1[43], w1_s0[43]}), .c ({new_AGEMA_signal_5863, addc_in[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_44_U1 ( .s (p256_sel), .b ({w0_s1[44], w0_s0[44]}), .a ({w1_s1[44], w1_s0[44]}), .c ({new_AGEMA_signal_5866, addc_in[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_45_U1 ( .s (p256_sel), .b ({w0_s1[45], w0_s0[45]}), .a ({w1_s1[45], w1_s0[45]}), .c ({new_AGEMA_signal_5869, addc_in[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_46_U1 ( .s (p256_sel), .b ({w0_s1[46], w0_s0[46]}), .a ({w1_s1[46], w1_s0[46]}), .c ({new_AGEMA_signal_5872, addc_in[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_47_U1 ( .s (p256_sel), .b ({w0_s1[47], w0_s0[47]}), .a ({w1_s1[47], w1_s0[47]}), .c ({new_AGEMA_signal_5875, addc_in[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_48_U1 ( .s (p256_sel), .b ({w0_s1[48], w0_s0[48]}), .a ({w1_s1[48], w1_s0[48]}), .c ({new_AGEMA_signal_5878, addc_in[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_49_U1 ( .s (p256_sel), .b ({w0_s1[49], w0_s0[49]}), .a ({w1_s1[49], w1_s0[49]}), .c ({new_AGEMA_signal_5881, addc_in[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_50_U1 ( .s (p256_sel), .b ({w0_s1[50], w0_s0[50]}), .a ({w1_s1[50], w1_s0[50]}), .c ({new_AGEMA_signal_5884, addc_in[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_51_U1 ( .s (p256_sel), .b ({w0_s1[51], w0_s0[51]}), .a ({w1_s1[51], w1_s0[51]}), .c ({new_AGEMA_signal_5887, addc_in[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_52_U1 ( .s (p256_sel), .b ({w0_s1[52], w0_s0[52]}), .a ({w1_s1[52], w1_s0[52]}), .c ({new_AGEMA_signal_5890, addc_in[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_53_U1 ( .s (p256_sel), .b ({w0_s1[53], w0_s0[53]}), .a ({w1_s1[53], w1_s0[53]}), .c ({new_AGEMA_signal_5893, addc_in[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_54_U1 ( .s (p256_sel), .b ({w0_s1[54], w0_s0[54]}), .a ({w1_s1[54], w1_s0[54]}), .c ({new_AGEMA_signal_5896, addc_in[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_55_U1 ( .s (p256_sel), .b ({w0_s1[55], w0_s0[55]}), .a ({w1_s1[55], w1_s0[55]}), .c ({new_AGEMA_signal_5899, addc_in[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_56_U1 ( .s (p256_sel), .b ({w0_s1[56], w0_s0[56]}), .a ({w1_s1[56], w1_s0[56]}), .c ({new_AGEMA_signal_5902, addc_in[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_57_U1 ( .s (p256_sel), .b ({w0_s1[57], w0_s0[57]}), .a ({w1_s1[57], w1_s0[57]}), .c ({new_AGEMA_signal_5905, addc_in[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_58_U1 ( .s (p256_sel), .b ({w0_s1[58], w0_s0[58]}), .a ({w1_s1[58], w1_s0[58]}), .c ({new_AGEMA_signal_5908, addc_in[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_59_U1 ( .s (p256_sel), .b ({w0_s1[59], w0_s0[59]}), .a ({w1_s1[59], w1_s0[59]}), .c ({new_AGEMA_signal_5911, addc_in[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_60_U1 ( .s (p256_sel), .b ({w0_s1[60], w0_s0[60]}), .a ({w1_s1[60], w1_s0[60]}), .c ({new_AGEMA_signal_5914, addc_in[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_61_U1 ( .s (p256_sel), .b ({w0_s1[61], w0_s0[61]}), .a ({w1_s1[61], w1_s0[61]}), .c ({new_AGEMA_signal_5917, addc_in[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_62_U1 ( .s (p256_sel), .b ({w0_s1[62], w0_s0[62]}), .a ({w1_s1[62], w1_s0[62]}), .c ({new_AGEMA_signal_5920, addc_in[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_63_U1 ( .s (p256_sel), .b ({w0_s1[63], w0_s0[63]}), .a ({w1_s1[63], w1_s0[63]}), .c ({new_AGEMA_signal_5923, addc_in[63]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_64_U1 ( .s (p256_sel), .b ({w0_s1[64], w0_s0[64]}), .a ({w1_s1[64], w1_s0[64]}), .c ({new_AGEMA_signal_5926, addc_in[64]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_65_U1 ( .s (p256_sel), .b ({w0_s1[65], w0_s0[65]}), .a ({w1_s1[65], w1_s0[65]}), .c ({new_AGEMA_signal_5929, addc_in[65]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_66_U1 ( .s (p256_sel), .b ({w0_s1[66], w0_s0[66]}), .a ({w1_s1[66], w1_s0[66]}), .c ({new_AGEMA_signal_5932, addc_in[66]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_67_U1 ( .s (p256_sel), .b ({w0_s1[67], w0_s0[67]}), .a ({w1_s1[67], w1_s0[67]}), .c ({new_AGEMA_signal_5935, addc_in[67]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_68_U1 ( .s (p256_sel), .b ({w0_s1[68], w0_s0[68]}), .a ({w1_s1[68], w1_s0[68]}), .c ({new_AGEMA_signal_5938, addc_in[68]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_69_U1 ( .s (p256_sel), .b ({w0_s1[69], w0_s0[69]}), .a ({w1_s1[69], w1_s0[69]}), .c ({new_AGEMA_signal_5941, addc_in[69]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_70_U1 ( .s (p256_sel), .b ({w0_s1[70], w0_s0[70]}), .a ({w1_s1[70], w1_s0[70]}), .c ({new_AGEMA_signal_5944, addc_in[70]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_71_U1 ( .s (p256_sel), .b ({w0_s1[71], w0_s0[71]}), .a ({w1_s1[71], w1_s0[71]}), .c ({new_AGEMA_signal_5947, addc_in[71]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_72_U1 ( .s (p256_sel), .b ({w0_s1[72], w0_s0[72]}), .a ({w1_s1[72], w1_s0[72]}), .c ({new_AGEMA_signal_5950, addc_in[72]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_73_U1 ( .s (p256_sel), .b ({w0_s1[73], w0_s0[73]}), .a ({w1_s1[73], w1_s0[73]}), .c ({new_AGEMA_signal_5953, addc_in[73]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_74_U1 ( .s (p256_sel), .b ({w0_s1[74], w0_s0[74]}), .a ({w1_s1[74], w1_s0[74]}), .c ({new_AGEMA_signal_5956, addc_in[74]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_75_U1 ( .s (p256_sel), .b ({w0_s1[75], w0_s0[75]}), .a ({w1_s1[75], w1_s0[75]}), .c ({new_AGEMA_signal_5959, addc_in[75]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_76_U1 ( .s (p256_sel), .b ({w0_s1[76], w0_s0[76]}), .a ({w1_s1[76], w1_s0[76]}), .c ({new_AGEMA_signal_5962, addc_in[76]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_77_U1 ( .s (p256_sel), .b ({w0_s1[77], w0_s0[77]}), .a ({w1_s1[77], w1_s0[77]}), .c ({new_AGEMA_signal_5965, addc_in[77]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_78_U1 ( .s (p256_sel), .b ({w0_s1[78], w0_s0[78]}), .a ({w1_s1[78], w1_s0[78]}), .c ({new_AGEMA_signal_5968, addc_in[78]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_79_U1 ( .s (p256_sel), .b ({w0_s1[79], w0_s0[79]}), .a ({w1_s1[79], w1_s0[79]}), .c ({new_AGEMA_signal_5971, addc_in[79]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_80_U1 ( .s (p256_sel), .b ({w0_s1[80], w0_s0[80]}), .a ({w1_s1[80], w1_s0[80]}), .c ({new_AGEMA_signal_5974, addc_in[80]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_81_U1 ( .s (p256_sel), .b ({w0_s1[81], w0_s0[81]}), .a ({w1_s1[81], w1_s0[81]}), .c ({new_AGEMA_signal_5977, addc_in[81]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_82_U1 ( .s (p256_sel), .b ({w0_s1[82], w0_s0[82]}), .a ({w1_s1[82], w1_s0[82]}), .c ({new_AGEMA_signal_5980, addc_in[82]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_83_U1 ( .s (p256_sel), .b ({w0_s1[83], w0_s0[83]}), .a ({w1_s1[83], w1_s0[83]}), .c ({new_AGEMA_signal_5983, addc_in[83]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_84_U1 ( .s (p256_sel), .b ({w0_s1[84], w0_s0[84]}), .a ({w1_s1[84], w1_s0[84]}), .c ({new_AGEMA_signal_5986, addc_in[84]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_85_U1 ( .s (p256_sel), .b ({w0_s1[85], w0_s0[85]}), .a ({w1_s1[85], w1_s0[85]}), .c ({new_AGEMA_signal_5989, addc_in[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_86_U1 ( .s (p256_sel), .b ({w0_s1[86], w0_s0[86]}), .a ({w1_s1[86], w1_s0[86]}), .c ({new_AGEMA_signal_5992, addc_in[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_87_U1 ( .s (p256_sel), .b ({w0_s1[87], w0_s0[87]}), .a ({w1_s1[87], w1_s0[87]}), .c ({new_AGEMA_signal_5995, addc_in[87]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_88_U1 ( .s (p256_sel), .b ({w0_s1[88], w0_s0[88]}), .a ({w1_s1[88], w1_s0[88]}), .c ({new_AGEMA_signal_5998, addc_in[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_89_U1 ( .s (p256_sel), .b ({w0_s1[89], w0_s0[89]}), .a ({w1_s1[89], w1_s0[89]}), .c ({new_AGEMA_signal_6001, addc_in[89]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_90_U1 ( .s (p256_sel), .b ({w0_s1[90], w0_s0[90]}), .a ({w1_s1[90], w1_s0[90]}), .c ({new_AGEMA_signal_6004, addc_in[90]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_91_U1 ( .s (p256_sel), .b ({w0_s1[91], w0_s0[91]}), .a ({w1_s1[91], w1_s0[91]}), .c ({new_AGEMA_signal_6007, addc_in[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_92_U1 ( .s (p256_sel), .b ({w0_s1[92], w0_s0[92]}), .a ({w1_s1[92], w1_s0[92]}), .c ({new_AGEMA_signal_6010, addc_in[92]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_93_U1 ( .s (p256_sel), .b ({w0_s1[93], w0_s0[93]}), .a ({w1_s1[93], w1_s0[93]}), .c ({new_AGEMA_signal_6013, addc_in[93]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_94_U1 ( .s (p256_sel), .b ({w0_s1[94], w0_s0[94]}), .a ({w1_s1[94], w1_s0[94]}), .c ({new_AGEMA_signal_6016, addc_in[94]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_95_U1 ( .s (p256_sel), .b ({w0_s1[95], w0_s0[95]}), .a ({w1_s1[95], w1_s0[95]}), .c ({new_AGEMA_signal_6019, addc_in[95]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_96_U1 ( .s (p256_sel), .b ({w0_s1[96], w0_s0[96]}), .a ({w1_s1[96], w1_s0[96]}), .c ({new_AGEMA_signal_6022, addc_in[96]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_97_U1 ( .s (p256_sel), .b ({w0_s1[97], w0_s0[97]}), .a ({w1_s1[97], w1_s0[97]}), .c ({new_AGEMA_signal_6025, addc_in[97]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_98_U1 ( .s (p256_sel), .b ({w0_s1[98], w0_s0[98]}), .a ({w1_s1[98], w1_s0[98]}), .c ({new_AGEMA_signal_6028, addc_in[98]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_99_U1 ( .s (p256_sel), .b ({w0_s1[99], w0_s0[99]}), .a ({w1_s1[99], w1_s0[99]}), .c ({new_AGEMA_signal_6031, addc_in[99]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_100_U1 ( .s (p256_sel), .b ({w0_s1[100], w0_s0[100]}), .a ({w1_s1[100], w1_s0[100]}), .c ({new_AGEMA_signal_6034, addc_in[100]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_101_U1 ( .s (p256_sel), .b ({w0_s1[101], w0_s0[101]}), .a ({w1_s1[101], w1_s0[101]}), .c ({new_AGEMA_signal_6037, addc_in[101]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_102_U1 ( .s (p256_sel), .b ({w0_s1[102], w0_s0[102]}), .a ({w1_s1[102], w1_s0[102]}), .c ({new_AGEMA_signal_6040, addc_in[102]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_103_U1 ( .s (p256_sel), .b ({w0_s1[103], w0_s0[103]}), .a ({w1_s1[103], w1_s0[103]}), .c ({new_AGEMA_signal_6043, addc_in[103]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_104_U1 ( .s (p256_sel), .b ({w0_s1[104], w0_s0[104]}), .a ({w1_s1[104], w1_s0[104]}), .c ({new_AGEMA_signal_6046, addc_in[104]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_105_U1 ( .s (p256_sel), .b ({w0_s1[105], w0_s0[105]}), .a ({w1_s1[105], w1_s0[105]}), .c ({new_AGEMA_signal_6049, addc_in[105]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_106_U1 ( .s (p256_sel), .b ({w0_s1[106], w0_s0[106]}), .a ({w1_s1[106], w1_s0[106]}), .c ({new_AGEMA_signal_6052, addc_in[106]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_107_U1 ( .s (p256_sel), .b ({w0_s1[107], w0_s0[107]}), .a ({w1_s1[107], w1_s0[107]}), .c ({new_AGEMA_signal_6055, addc_in[107]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_108_U1 ( .s (p256_sel), .b ({w0_s1[108], w0_s0[108]}), .a ({w1_s1[108], w1_s0[108]}), .c ({new_AGEMA_signal_6058, addc_in[108]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_109_U1 ( .s (p256_sel), .b ({w0_s1[109], w0_s0[109]}), .a ({w1_s1[109], w1_s0[109]}), .c ({new_AGEMA_signal_6061, addc_in[109]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_110_U1 ( .s (p256_sel), .b ({w0_s1[110], w0_s0[110]}), .a ({w1_s1[110], w1_s0[110]}), .c ({new_AGEMA_signal_6064, addc_in[110]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_111_U1 ( .s (p256_sel), .b ({w0_s1[111], w0_s0[111]}), .a ({w1_s1[111], w1_s0[111]}), .c ({new_AGEMA_signal_6067, addc_in[111]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_112_U1 ( .s (p256_sel), .b ({w0_s1[112], w0_s0[112]}), .a ({w1_s1[112], w1_s0[112]}), .c ({new_AGEMA_signal_6070, addc_in[112]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_113_U1 ( .s (p256_sel), .b ({w0_s1[113], w0_s0[113]}), .a ({w1_s1[113], w1_s0[113]}), .c ({new_AGEMA_signal_6073, addc_in[113]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_114_U1 ( .s (p256_sel), .b ({w0_s1[114], w0_s0[114]}), .a ({w1_s1[114], w1_s0[114]}), .c ({new_AGEMA_signal_6076, addc_in[114]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_115_U1 ( .s (p256_sel), .b ({w0_s1[115], w0_s0[115]}), .a ({w1_s1[115], w1_s0[115]}), .c ({new_AGEMA_signal_6079, addc_in[115]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_116_U1 ( .s (p256_sel), .b ({w0_s1[116], w0_s0[116]}), .a ({w1_s1[116], w1_s0[116]}), .c ({new_AGEMA_signal_6082, addc_in[116]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_117_U1 ( .s (p256_sel), .b ({w0_s1[117], w0_s0[117]}), .a ({w1_s1[117], w1_s0[117]}), .c ({new_AGEMA_signal_6085, addc_in[117]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_118_U1 ( .s (p256_sel), .b ({w0_s1[118], w0_s0[118]}), .a ({w1_s1[118], w1_s0[118]}), .c ({new_AGEMA_signal_6088, addc_in[118]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_119_U1 ( .s (p256_sel), .b ({w0_s1[119], w0_s0[119]}), .a ({w1_s1[119], w1_s0[119]}), .c ({new_AGEMA_signal_6091, addc_in[119]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_120_U1 ( .s (p256_sel), .b ({w0_s1[120], w0_s0[120]}), .a ({w1_s1[120], w1_s0[120]}), .c ({new_AGEMA_signal_6094, addc_in[120]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_121_U1 ( .s (p256_sel), .b ({w0_s1[121], w0_s0[121]}), .a ({w1_s1[121], w1_s0[121]}), .c ({new_AGEMA_signal_6097, addc_in[121]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_122_U1 ( .s (p256_sel), .b ({w0_s1[122], w0_s0[122]}), .a ({w1_s1[122], w1_s0[122]}), .c ({new_AGEMA_signal_6100, addc_in[122]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_123_U1 ( .s (p256_sel), .b ({w0_s1[123], w0_s0[123]}), .a ({w1_s1[123], w1_s0[123]}), .c ({new_AGEMA_signal_6103, addc_in[123]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_124_U1 ( .s (p256_sel), .b ({w0_s1[124], w0_s0[124]}), .a ({w1_s1[124], w1_s0[124]}), .c ({new_AGEMA_signal_6106, addc_in[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_125_U1 ( .s (p256_sel), .b ({w0_s1[125], w0_s0[125]}), .a ({w1_s1[125], w1_s0[125]}), .c ({new_AGEMA_signal_6109, addc_in[125]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_126_U1 ( .s (p256_sel), .b ({w0_s1[126], w0_s0[126]}), .a ({w1_s1[126], w1_s0[126]}), .c ({new_AGEMA_signal_6112, addc_in[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst1_MUXInst_127_U1 ( .s (p256_sel), .b ({w0_s1[127], w0_s0[127]}), .a ({w1_s1[127], w1_s0[127]}), .c ({new_AGEMA_signal_6115, addc_in[127]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_U8 ( .a ({new_AGEMA_signal_6116, add_sub1_0_n8}), .b ({1'b0, add_sub1_0_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_6632, add_sub1_0_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_U7 ( .a ({new_AGEMA_signal_6115, addc_in[127]}), .b ({1'b0, p256_sel}), .c ({new_AGEMA_signal_6116, add_sub1_0_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_U6 ( .a ({new_AGEMA_signal_6320, add_sub1_0_n7}), .b ({1'b0, add_sub1_0_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_6633, add_sub1_0_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_U5 ( .a ({new_AGEMA_signal_6112, addc_in[126]}), .b ({1'b0, add_sub1_0_addc_rom_ic_out[2]}), .c ({new_AGEMA_signal_6320, add_sub1_0_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_U4 ( .a ({new_AGEMA_signal_6117, add_sub1_0_n6}), .b ({1'b0, add_sub1_0_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_6634, add_sub1_0_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_U3 ( .a ({new_AGEMA_signal_6109, addc_in[125]}), .b ({1'b0, add_sub1_0_addc_rom_ic_out[1]}), .c ({new_AGEMA_signal_6117, add_sub1_0_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_U2 ( .a ({new_AGEMA_signal_6548, add_sub1_0_n5}), .b ({1'b0, add_sub1_0_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_6635, add_sub1_0_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_U1 ( .a ({new_AGEMA_signal_6106, addc_in[124]}), .b ({1'b0, add_sub1_0_addc_rom_ic_out[0]}), .c ({new_AGEMA_signal_6548, add_sub1_0_n5}) ) ;
    XOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U4 ( .A (1'b0), .B (p256_sel), .Z (add_sub1_0_addc_rom_ic_out[1]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_0_addc_rom_ic1_ANF_0_n2), .B (1'b0), .ZN (add_sub1_0_addc_rom_ic_out[0]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U2 ( .A (1'b0), .B (add_sub1_0_addc_rom_ic_out[2]), .ZN (add_sub1_0_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_0_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_0_addc_rom_ic_out[2]) ) ;
    AND2_X1 add_sub1_0_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b0), .A2 (1'b0), .ZN (add_sub1_0_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n21), .B (add_sub1_0_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_0_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n19), .B (add_sub1_0_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t5), .B (add_sub1_0_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t7), .B (add_sub1_0_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n17), .B (add_sub1_0_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_0_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t6), .B (add_sub1_0_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n14), .B (add_sub1_0_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_0_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t5), .B (add_sub1_0_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_0_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_0_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n12), .B (add_sub1_0_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_0_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t0), .B (add_sub1_0_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t4), .B (add_sub1_0_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_0_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_0_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_0_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_0_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_6632, add_sub1_0_addc_out[3]}), .b ({new_AGEMA_signal_6633, add_sub1_0_addc_out[2]}), .c ({new_AGEMA_signal_6868, add_sub1_0_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_6634, add_sub1_0_addc_out[1]}), .b ({new_AGEMA_signal_6633, add_sub1_0_addc_out[2]}), .c ({new_AGEMA_signal_6869, add_sub1_0_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_6103, addc_in[123]}), .b ({new_AGEMA_signal_6100, addc_in[122]}), .c ({new_AGEMA_signal_6118, add_sub1_0_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_6097, addc_in[121]}), .b ({new_AGEMA_signal_6100, addc_in[122]}), .c ({new_AGEMA_signal_6119, add_sub1_0_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_6091, addc_in[119]}), .b ({new_AGEMA_signal_6088, addc_in[118]}), .c ({new_AGEMA_signal_6125, add_sub1_0_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_6085, addc_in[117]}), .b ({new_AGEMA_signal_6088, addc_in[118]}), .c ({new_AGEMA_signal_6126, add_sub1_0_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_6079, addc_in[115]}), .b ({new_AGEMA_signal_6076, addc_in[114]}), .c ({new_AGEMA_signal_6132, add_sub1_0_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_6073, addc_in[113]}), .b ({new_AGEMA_signal_6076, addc_in[114]}), .c ({new_AGEMA_signal_6133, add_sub1_0_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_6067, addc_in[111]}), .b ({new_AGEMA_signal_6064, addc_in[110]}), .c ({new_AGEMA_signal_6139, add_sub1_0_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_6061, addc_in[109]}), .b ({new_AGEMA_signal_6064, addc_in[110]}), .c ({new_AGEMA_signal_6140, add_sub1_0_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_6055, addc_in[107]}), .b ({new_AGEMA_signal_6052, addc_in[106]}), .c ({new_AGEMA_signal_6146, add_sub1_0_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_6049, addc_in[105]}), .b ({new_AGEMA_signal_6052, addc_in[106]}), .c ({new_AGEMA_signal_6147, add_sub1_0_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_6043, addc_in[103]}), .b ({new_AGEMA_signal_6040, addc_in[102]}), .c ({new_AGEMA_signal_6153, add_sub1_0_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_6037, addc_in[101]}), .b ({new_AGEMA_signal_6040, addc_in[102]}), .c ({new_AGEMA_signal_6154, add_sub1_0_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_6031, addc_in[99]}), .b ({new_AGEMA_signal_6028, addc_in[98]}), .c ({new_AGEMA_signal_6160, add_sub1_0_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_6025, addc_in[97]}), .b ({new_AGEMA_signal_6028, addc_in[98]}), .c ({new_AGEMA_signal_6161, add_sub1_0_subc_rom_sbox_0_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_U8 ( .a ({new_AGEMA_signal_6167, add_sub1_1_n8}), .b ({1'b0, add_sub1_1_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_6643, add_sub1_1_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_U7 ( .a ({new_AGEMA_signal_6019, addc_in[95]}), .b ({1'b0, p256_sel}), .c ({new_AGEMA_signal_6167, add_sub1_1_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_U6 ( .a ({new_AGEMA_signal_6356, add_sub1_1_n7}), .b ({1'b0, add_sub1_1_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_6644, add_sub1_1_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_U5 ( .a ({new_AGEMA_signal_6016, addc_in[94]}), .b ({1'b0, add_sub1_1_addc_rom_ic_out[2]}), .c ({new_AGEMA_signal_6356, add_sub1_1_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_U4 ( .a ({new_AGEMA_signal_6168, add_sub1_1_n6}), .b ({1'b0, add_sub1_1_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_6645, add_sub1_1_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_U3 ( .a ({new_AGEMA_signal_6013, addc_in[93]}), .b ({1'b0, add_sub1_1_addc_rom_ic_out[1]}), .c ({new_AGEMA_signal_6168, add_sub1_1_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_U2 ( .a ({new_AGEMA_signal_6563, add_sub1_1_n5}), .b ({1'b0, add_sub1_1_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_6646, add_sub1_1_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_U1 ( .a ({new_AGEMA_signal_6010, addc_in[92]}), .b ({1'b0, add_sub1_1_addc_rom_ic_out[0]}), .c ({new_AGEMA_signal_6563, add_sub1_1_n5}) ) ;
    XOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U4 ( .A (1'b0), .B (p256_sel), .Z (add_sub1_1_addc_rom_ic_out[1]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_1_addc_rom_ic1_ANF_0_n2), .B (1'b1), .ZN (add_sub1_1_addc_rom_ic_out[0]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U2 ( .A (1'b0), .B (add_sub1_1_addc_rom_ic_out[2]), .ZN (add_sub1_1_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_1_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_1_addc_rom_ic_out[2]) ) ;
    AND2_X1 add_sub1_1_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b1), .A2 (1'b0), .ZN (add_sub1_1_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n21), .B (add_sub1_1_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_1_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n19), .B (add_sub1_1_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t5), .B (add_sub1_1_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t7), .B (add_sub1_1_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n17), .B (add_sub1_1_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_1_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t6), .B (add_sub1_1_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n14), .B (add_sub1_1_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_1_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t5), .B (add_sub1_1_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_1_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_1_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n12), .B (add_sub1_1_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_1_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t0), .B (add_sub1_1_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t4), .B (add_sub1_1_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_1_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_1_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_1_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_1_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_6643, add_sub1_1_addc_out[3]}), .b ({new_AGEMA_signal_6644, add_sub1_1_addc_out[2]}), .c ({new_AGEMA_signal_6889, add_sub1_1_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_6645, add_sub1_1_addc_out[1]}), .b ({new_AGEMA_signal_6644, add_sub1_1_addc_out[2]}), .c ({new_AGEMA_signal_6890, add_sub1_1_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_6007, addc_in[91]}), .b ({new_AGEMA_signal_6004, addc_in[90]}), .c ({new_AGEMA_signal_6169, add_sub1_1_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_6001, addc_in[89]}), .b ({new_AGEMA_signal_6004, addc_in[90]}), .c ({new_AGEMA_signal_6170, add_sub1_1_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_5995, addc_in[87]}), .b ({new_AGEMA_signal_5992, addc_in[86]}), .c ({new_AGEMA_signal_6176, add_sub1_1_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_5989, addc_in[85]}), .b ({new_AGEMA_signal_5992, addc_in[86]}), .c ({new_AGEMA_signal_6177, add_sub1_1_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_5983, addc_in[83]}), .b ({new_AGEMA_signal_5980, addc_in[82]}), .c ({new_AGEMA_signal_6183, add_sub1_1_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_5977, addc_in[81]}), .b ({new_AGEMA_signal_5980, addc_in[82]}), .c ({new_AGEMA_signal_6184, add_sub1_1_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_5971, addc_in[79]}), .b ({new_AGEMA_signal_5968, addc_in[78]}), .c ({new_AGEMA_signal_6190, add_sub1_1_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_5965, addc_in[77]}), .b ({new_AGEMA_signal_5968, addc_in[78]}), .c ({new_AGEMA_signal_6191, add_sub1_1_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_5959, addc_in[75]}), .b ({new_AGEMA_signal_5956, addc_in[74]}), .c ({new_AGEMA_signal_6197, add_sub1_1_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_5953, addc_in[73]}), .b ({new_AGEMA_signal_5956, addc_in[74]}), .c ({new_AGEMA_signal_6198, add_sub1_1_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_5947, addc_in[71]}), .b ({new_AGEMA_signal_5944, addc_in[70]}), .c ({new_AGEMA_signal_6204, add_sub1_1_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_5941, addc_in[69]}), .b ({new_AGEMA_signal_5944, addc_in[70]}), .c ({new_AGEMA_signal_6205, add_sub1_1_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_5935, addc_in[67]}), .b ({new_AGEMA_signal_5932, addc_in[66]}), .c ({new_AGEMA_signal_6211, add_sub1_1_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_5929, addc_in[65]}), .b ({new_AGEMA_signal_5932, addc_in[66]}), .c ({new_AGEMA_signal_6212, add_sub1_1_subc_rom_sbox_0_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_U8 ( .a ({new_AGEMA_signal_6218, add_sub1_2_n8}), .b ({1'b0, add_sub1_2_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_6654, add_sub1_2_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_U7 ( .a ({new_AGEMA_signal_5923, addc_in[63]}), .b ({1'b0, p256_sel}), .c ({new_AGEMA_signal_6218, add_sub1_2_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_U6 ( .a ({new_AGEMA_signal_6392, add_sub1_2_n7}), .b ({1'b0, add_sub1_2_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_6655, add_sub1_2_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_U5 ( .a ({new_AGEMA_signal_5920, addc_in[62]}), .b ({1'b0, add_sub1_2_addc_rom_ic_out[2]}), .c ({new_AGEMA_signal_6392, add_sub1_2_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_U4 ( .a ({new_AGEMA_signal_6219, add_sub1_2_n6}), .b ({1'b0, add_sub1_2_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_6656, add_sub1_2_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_U3 ( .a ({new_AGEMA_signal_5917, addc_in[61]}), .b ({1'b0, add_sub1_2_addc_rom_ic_out[1]}), .c ({new_AGEMA_signal_6219, add_sub1_2_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_U2 ( .a ({new_AGEMA_signal_6578, add_sub1_2_n5}), .b ({1'b0, add_sub1_2_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_6657, add_sub1_2_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_U1 ( .a ({new_AGEMA_signal_5914, addc_in[60]}), .b ({1'b0, add_sub1_2_addc_rom_ic_out[0]}), .c ({new_AGEMA_signal_6578, add_sub1_2_n5}) ) ;
    XOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U4 ( .A (1'b1), .B (p256_sel), .Z (add_sub1_2_addc_rom_ic_out[1]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_2_addc_rom_ic1_ANF_0_n2), .B (1'b0), .ZN (add_sub1_2_addc_rom_ic_out[0]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U2 ( .A (1'b1), .B (add_sub1_2_addc_rom_ic_out[2]), .ZN (add_sub1_2_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_2_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_2_addc_rom_ic_out[2]) ) ;
    AND2_X1 add_sub1_2_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b0), .A2 (1'b1), .ZN (add_sub1_2_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n21), .B (add_sub1_2_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_2_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n19), .B (add_sub1_2_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t5), .B (add_sub1_2_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t7), .B (add_sub1_2_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n17), .B (add_sub1_2_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_2_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t6), .B (add_sub1_2_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n14), .B (add_sub1_2_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_2_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t5), .B (add_sub1_2_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_2_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_2_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n12), .B (add_sub1_2_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_2_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t0), .B (add_sub1_2_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t4), .B (add_sub1_2_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_2_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_2_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_2_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_2_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_6654, add_sub1_2_addc_out[3]}), .b ({new_AGEMA_signal_6655, add_sub1_2_addc_out[2]}), .c ({new_AGEMA_signal_6910, add_sub1_2_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_6656, add_sub1_2_addc_out[1]}), .b ({new_AGEMA_signal_6655, add_sub1_2_addc_out[2]}), .c ({new_AGEMA_signal_6911, add_sub1_2_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_5911, addc_in[59]}), .b ({new_AGEMA_signal_5908, addc_in[58]}), .c ({new_AGEMA_signal_6220, add_sub1_2_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_5905, addc_in[57]}), .b ({new_AGEMA_signal_5908, addc_in[58]}), .c ({new_AGEMA_signal_6221, add_sub1_2_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_5899, addc_in[55]}), .b ({new_AGEMA_signal_5896, addc_in[54]}), .c ({new_AGEMA_signal_6227, add_sub1_2_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_5893, addc_in[53]}), .b ({new_AGEMA_signal_5896, addc_in[54]}), .c ({new_AGEMA_signal_6228, add_sub1_2_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_5887, addc_in[51]}), .b ({new_AGEMA_signal_5884, addc_in[50]}), .c ({new_AGEMA_signal_6234, add_sub1_2_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_5881, addc_in[49]}), .b ({new_AGEMA_signal_5884, addc_in[50]}), .c ({new_AGEMA_signal_6235, add_sub1_2_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_5875, addc_in[47]}), .b ({new_AGEMA_signal_5872, addc_in[46]}), .c ({new_AGEMA_signal_6241, add_sub1_2_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_5869, addc_in[45]}), .b ({new_AGEMA_signal_5872, addc_in[46]}), .c ({new_AGEMA_signal_6242, add_sub1_2_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_5863, addc_in[43]}), .b ({new_AGEMA_signal_5860, addc_in[42]}), .c ({new_AGEMA_signal_6248, add_sub1_2_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_5857, addc_in[41]}), .b ({new_AGEMA_signal_5860, addc_in[42]}), .c ({new_AGEMA_signal_6249, add_sub1_2_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_5851, addc_in[39]}), .b ({new_AGEMA_signal_5848, addc_in[38]}), .c ({new_AGEMA_signal_6255, add_sub1_2_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_5845, addc_in[37]}), .b ({new_AGEMA_signal_5848, addc_in[38]}), .c ({new_AGEMA_signal_6256, add_sub1_2_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_5839, addc_in[35]}), .b ({new_AGEMA_signal_5836, addc_in[34]}), .c ({new_AGEMA_signal_6262, add_sub1_2_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_5833, addc_in[33]}), .b ({new_AGEMA_signal_5836, addc_in[34]}), .c ({new_AGEMA_signal_6263, add_sub1_2_subc_rom_sbox_0_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_U8 ( .a ({new_AGEMA_signal_6269, add_sub1_3_n8}), .b ({1'b0, add_sub1_3_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_6665, add_sub1_3_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_U7 ( .a ({new_AGEMA_signal_5827, addc_in[31]}), .b ({1'b0, p256_sel}), .c ({new_AGEMA_signal_6269, add_sub1_3_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_U6 ( .a ({new_AGEMA_signal_6428, add_sub1_3_n7}), .b ({1'b0, add_sub1_3_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_6666, add_sub1_3_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_U5 ( .a ({new_AGEMA_signal_5824, addc_in[30]}), .b ({1'b0, add_sub1_3_addc_rom_ic_out_2_}), .c ({new_AGEMA_signal_6428, add_sub1_3_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_U4 ( .a ({new_AGEMA_signal_6270, add_sub1_3_n6}), .b ({1'b0, add_sub1_3_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_6667, add_sub1_3_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_U3 ( .a ({new_AGEMA_signal_5821, addc_in[29]}), .b ({1'b0, add_sub1_3_addc_rom_ic_out_1_}), .c ({new_AGEMA_signal_6270, add_sub1_3_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_U2 ( .a ({new_AGEMA_signal_6593, add_sub1_3_n5}), .b ({1'b0, add_sub1_3_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_6668, add_sub1_3_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_U1 ( .a ({new_AGEMA_signal_5818, addc_in[28]}), .b ({1'b0, add_sub1_3_addc_rom_ic_out_0_}), .c ({new_AGEMA_signal_6593, add_sub1_3_n5}) ) ;
    XOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U4 ( .A (1'b1), .B (p256_sel), .Z (add_sub1_3_addc_rom_ic_out_1_) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_3_addc_rom_ic1_ANF_0_n2), .B (1'b1), .ZN (add_sub1_3_addc_rom_ic_out_0_) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U2 ( .A (1'b1), .B (add_sub1_3_addc_rom_ic_out_2_), .ZN (add_sub1_3_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_3_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_3_addc_rom_ic_out_2_) ) ;
    AND2_X1 add_sub1_3_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b1), .A2 (1'b1), .ZN (add_sub1_3_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n21), .B (add_sub1_3_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_3_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n19), .B (add_sub1_3_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t5), .B (add_sub1_3_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t7), .B (add_sub1_3_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n17), .B (add_sub1_3_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_3_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t6), .B (add_sub1_3_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n14), .B (add_sub1_3_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_3_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t5), .B (add_sub1_3_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_3_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_3_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n12), .B (add_sub1_3_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_3_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t0), .B (add_sub1_3_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t4), .B (add_sub1_3_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_3_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_3_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_3_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_3_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_6665, add_sub1_3_addc_out[3]}), .b ({new_AGEMA_signal_6666, add_sub1_3_addc_out[2]}), .c ({new_AGEMA_signal_6931, add_sub1_3_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_6667, add_sub1_3_addc_out[1]}), .b ({new_AGEMA_signal_6666, add_sub1_3_addc_out[2]}), .c ({new_AGEMA_signal_6932, add_sub1_3_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_5815, addc_in[27]}), .b ({new_AGEMA_signal_5812, addc_in[26]}), .c ({new_AGEMA_signal_6271, add_sub1_3_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_5809, addc_in[25]}), .b ({new_AGEMA_signal_5812, addc_in[26]}), .c ({new_AGEMA_signal_6272, add_sub1_3_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_5803, addc_in[23]}), .b ({new_AGEMA_signal_5800, addc_in[22]}), .c ({new_AGEMA_signal_6278, add_sub1_3_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_5797, addc_in[21]}), .b ({new_AGEMA_signal_5800, addc_in[22]}), .c ({new_AGEMA_signal_6279, add_sub1_3_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_5791, addc_in[19]}), .b ({new_AGEMA_signal_5788, addc_in[18]}), .c ({new_AGEMA_signal_6285, add_sub1_3_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_5785, addc_in[17]}), .b ({new_AGEMA_signal_5788, addc_in[18]}), .c ({new_AGEMA_signal_6286, add_sub1_3_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_5779, addc_in[15]}), .b ({new_AGEMA_signal_5776, addc_in[14]}), .c ({new_AGEMA_signal_6292, add_sub1_3_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_5773, addc_in[13]}), .b ({new_AGEMA_signal_5776, addc_in[14]}), .c ({new_AGEMA_signal_6293, add_sub1_3_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_5767, addc_in[11]}), .b ({new_AGEMA_signal_5764, addc_in[10]}), .c ({new_AGEMA_signal_6299, add_sub1_3_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_5761, addc_in[9]}), .b ({new_AGEMA_signal_5764, addc_in[10]}), .c ({new_AGEMA_signal_6300, add_sub1_3_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_5755, addc_in[7]}), .b ({new_AGEMA_signal_5752, addc_in[6]}), .c ({new_AGEMA_signal_6306, add_sub1_3_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_5749, addc_in[5]}), .b ({new_AGEMA_signal_5752, addc_in[6]}), .c ({new_AGEMA_signal_6307, add_sub1_3_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_5743, addc_in[3]}), .b ({new_AGEMA_signal_5740, addc_in[2]}), .c ({new_AGEMA_signal_6313, add_sub1_3_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_5737, addc_in[1]}), .b ({new_AGEMA_signal_5740, addc_in[2]}), .c ({new_AGEMA_signal_6314, add_sub1_3_subc_rom_sbox_0_ANF_2_t5}) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_7175, add_sub1_0_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_7174, add_sub1_0_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_7276, add_sub1_0_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_6871, add_sub1_0_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_6873, add_sub1_0_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_7174, add_sub1_0_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_6874, add_sub1_0_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_6633, add_sub1_0_addc_out[2]}), .c ({new_AGEMA_signal_7175, add_sub1_0_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_6868, add_sub1_0_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_7176, add_sub1_0_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_7278, subc_out[124]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_6870, add_sub1_0_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_6635, add_sub1_0_addc_out[0]}), .c ({new_AGEMA_signal_7176, add_sub1_0_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6634, add_sub1_0_addc_out[1]}), .b ({new_AGEMA_signal_6633, add_sub1_0_addc_out[2]}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_6870, add_sub1_0_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6634, add_sub1_0_addc_out[1]}), .b ({new_AGEMA_signal_6632, add_sub1_0_addc_out[3]}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_6871, add_sub1_0_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6633, add_sub1_0_addc_out[2]}), .b ({new_AGEMA_signal_6632, add_sub1_0_addc_out[3]}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_6872, add_sub1_0_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6635, add_sub1_0_addc_out[0]}), .b ({new_AGEMA_signal_6632, add_sub1_0_addc_out[3]}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_6873, add_sub1_0_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6635, add_sub1_0_addc_out[0]}), .b ({new_AGEMA_signal_6634, add_sub1_0_addc_out[1]}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_6874, add_sub1_0_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_6322, add_sub1_0_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_6321, add_sub1_0_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_6464, add_sub1_0_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_6121, add_sub1_0_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_6123, add_sub1_0_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_6321, add_sub1_0_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_6124, add_sub1_0_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_6100, addc_in[122]}), .c ({new_AGEMA_signal_6322, add_sub1_0_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_6118, add_sub1_0_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_6323, add_sub1_0_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_6466, subc_out[120]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_6120, add_sub1_0_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_6094, addc_in[120]}), .c ({new_AGEMA_signal_6323, add_sub1_0_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6097, addc_in[121]}), .b ({new_AGEMA_signal_6100, addc_in[122]}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_6120, add_sub1_0_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6097, addc_in[121]}), .b ({new_AGEMA_signal_6103, addc_in[123]}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_6121, add_sub1_0_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6100, addc_in[122]}), .b ({new_AGEMA_signal_6103, addc_in[123]}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_6122, add_sub1_0_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6094, addc_in[120]}), .b ({new_AGEMA_signal_6103, addc_in[123]}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_6123, add_sub1_0_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6094, addc_in[120]}), .b ({new_AGEMA_signal_6097, addc_in[121]}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_6124, add_sub1_0_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_6327, add_sub1_0_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_6326, add_sub1_0_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_6467, add_sub1_0_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_6128, add_sub1_0_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_6130, add_sub1_0_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_6326, add_sub1_0_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_6131, add_sub1_0_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_6088, addc_in[118]}), .c ({new_AGEMA_signal_6327, add_sub1_0_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_6125, add_sub1_0_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_6328, add_sub1_0_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_6469, subc_out[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_6127, add_sub1_0_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_6082, addc_in[116]}), .c ({new_AGEMA_signal_6328, add_sub1_0_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6085, addc_in[117]}), .b ({new_AGEMA_signal_6088, addc_in[118]}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_6127, add_sub1_0_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6085, addc_in[117]}), .b ({new_AGEMA_signal_6091, addc_in[119]}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_6128, add_sub1_0_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6088, addc_in[118]}), .b ({new_AGEMA_signal_6091, addc_in[119]}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_6129, add_sub1_0_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6082, addc_in[116]}), .b ({new_AGEMA_signal_6091, addc_in[119]}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_6130, add_sub1_0_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6082, addc_in[116]}), .b ({new_AGEMA_signal_6085, addc_in[117]}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_6131, add_sub1_0_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_6332, add_sub1_0_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_6331, add_sub1_0_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_6470, add_sub1_0_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_6135, add_sub1_0_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_6137, add_sub1_0_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_6331, add_sub1_0_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_6138, add_sub1_0_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_6076, addc_in[114]}), .c ({new_AGEMA_signal_6332, add_sub1_0_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_6132, add_sub1_0_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_6333, add_sub1_0_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_6472, subc_out[112]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_6134, add_sub1_0_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_6070, addc_in[112]}), .c ({new_AGEMA_signal_6333, add_sub1_0_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6073, addc_in[113]}), .b ({new_AGEMA_signal_6076, addc_in[114]}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_6134, add_sub1_0_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6073, addc_in[113]}), .b ({new_AGEMA_signal_6079, addc_in[115]}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_6135, add_sub1_0_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6076, addc_in[114]}), .b ({new_AGEMA_signal_6079, addc_in[115]}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_6136, add_sub1_0_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6070, addc_in[112]}), .b ({new_AGEMA_signal_6079, addc_in[115]}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_6137, add_sub1_0_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6070, addc_in[112]}), .b ({new_AGEMA_signal_6073, addc_in[113]}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_6138, add_sub1_0_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_6337, add_sub1_0_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_6336, add_sub1_0_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_6473, add_sub1_0_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_6142, add_sub1_0_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_6144, add_sub1_0_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_6336, add_sub1_0_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_6145, add_sub1_0_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_6064, addc_in[110]}), .c ({new_AGEMA_signal_6337, add_sub1_0_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_6139, add_sub1_0_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_6338, add_sub1_0_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_6475, subc_out[108]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_6141, add_sub1_0_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_6058, addc_in[108]}), .c ({new_AGEMA_signal_6338, add_sub1_0_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6061, addc_in[109]}), .b ({new_AGEMA_signal_6064, addc_in[110]}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_6141, add_sub1_0_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6061, addc_in[109]}), .b ({new_AGEMA_signal_6067, addc_in[111]}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_6142, add_sub1_0_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6064, addc_in[110]}), .b ({new_AGEMA_signal_6067, addc_in[111]}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_6143, add_sub1_0_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6058, addc_in[108]}), .b ({new_AGEMA_signal_6067, addc_in[111]}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_6144, add_sub1_0_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6058, addc_in[108]}), .b ({new_AGEMA_signal_6061, addc_in[109]}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_6145, add_sub1_0_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_6342, add_sub1_0_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_6341, add_sub1_0_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_6476, add_sub1_0_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_6149, add_sub1_0_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_6151, add_sub1_0_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_6341, add_sub1_0_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_6152, add_sub1_0_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_6052, addc_in[106]}), .c ({new_AGEMA_signal_6342, add_sub1_0_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_6146, add_sub1_0_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_6343, add_sub1_0_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_6478, subc_out[104]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_6148, add_sub1_0_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_6046, addc_in[104]}), .c ({new_AGEMA_signal_6343, add_sub1_0_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6049, addc_in[105]}), .b ({new_AGEMA_signal_6052, addc_in[106]}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_6148, add_sub1_0_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6049, addc_in[105]}), .b ({new_AGEMA_signal_6055, addc_in[107]}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_6149, add_sub1_0_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6052, addc_in[106]}), .b ({new_AGEMA_signal_6055, addc_in[107]}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_6150, add_sub1_0_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6046, addc_in[104]}), .b ({new_AGEMA_signal_6055, addc_in[107]}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_6151, add_sub1_0_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6046, addc_in[104]}), .b ({new_AGEMA_signal_6049, addc_in[105]}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_6152, add_sub1_0_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_6347, add_sub1_0_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_6346, add_sub1_0_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_6479, add_sub1_0_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_6156, add_sub1_0_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_6158, add_sub1_0_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_6346, add_sub1_0_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_6159, add_sub1_0_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_6040, addc_in[102]}), .c ({new_AGEMA_signal_6347, add_sub1_0_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_6153, add_sub1_0_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_6348, add_sub1_0_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_6481, subc_out[100]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_6155, add_sub1_0_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_6034, addc_in[100]}), .c ({new_AGEMA_signal_6348, add_sub1_0_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6037, addc_in[101]}), .b ({new_AGEMA_signal_6040, addc_in[102]}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_6155, add_sub1_0_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6037, addc_in[101]}), .b ({new_AGEMA_signal_6043, addc_in[103]}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_6156, add_sub1_0_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6040, addc_in[102]}), .b ({new_AGEMA_signal_6043, addc_in[103]}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_6157, add_sub1_0_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6034, addc_in[100]}), .b ({new_AGEMA_signal_6043, addc_in[103]}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_6158, add_sub1_0_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6034, addc_in[100]}), .b ({new_AGEMA_signal_6037, addc_in[101]}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_6159, add_sub1_0_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_6352, add_sub1_0_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_6351, add_sub1_0_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_6482, add_sub1_0_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_6163, add_sub1_0_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_6165, add_sub1_0_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_6351, add_sub1_0_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_6166, add_sub1_0_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_6028, addc_in[98]}), .c ({new_AGEMA_signal_6352, add_sub1_0_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_6160, add_sub1_0_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_6353, add_sub1_0_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_6484, subc_out[96]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_6162, add_sub1_0_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_6022, addc_in[96]}), .c ({new_AGEMA_signal_6353, add_sub1_0_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6025, addc_in[97]}), .b ({new_AGEMA_signal_6028, addc_in[98]}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_6162, add_sub1_0_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6025, addc_in[97]}), .b ({new_AGEMA_signal_6031, addc_in[99]}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_6163, add_sub1_0_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6028, addc_in[98]}), .b ({new_AGEMA_signal_6031, addc_in[99]}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_6164, add_sub1_0_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6022, addc_in[96]}), .b ({new_AGEMA_signal_6031, addc_in[99]}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_6165, add_sub1_0_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6022, addc_in[96]}), .b ({new_AGEMA_signal_6025, addc_in[97]}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_6166, add_sub1_0_subc_rom_sbox_0_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_7187, add_sub1_1_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_7186, add_sub1_1_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_7279, add_sub1_1_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_6892, add_sub1_1_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_6894, add_sub1_1_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_7186, add_sub1_1_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_6895, add_sub1_1_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_6644, add_sub1_1_addc_out[2]}), .c ({new_AGEMA_signal_7187, add_sub1_1_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_6889, add_sub1_1_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_7188, add_sub1_1_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_7281, subc_out[92]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_6891, add_sub1_1_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_6646, add_sub1_1_addc_out[0]}), .c ({new_AGEMA_signal_7188, add_sub1_1_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6645, add_sub1_1_addc_out[1]}), .b ({new_AGEMA_signal_6644, add_sub1_1_addc_out[2]}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_6891, add_sub1_1_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6645, add_sub1_1_addc_out[1]}), .b ({new_AGEMA_signal_6643, add_sub1_1_addc_out[3]}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_6892, add_sub1_1_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6644, add_sub1_1_addc_out[2]}), .b ({new_AGEMA_signal_6643, add_sub1_1_addc_out[3]}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_6893, add_sub1_1_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6646, add_sub1_1_addc_out[0]}), .b ({new_AGEMA_signal_6643, add_sub1_1_addc_out[3]}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_6894, add_sub1_1_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6646, add_sub1_1_addc_out[0]}), .b ({new_AGEMA_signal_6645, add_sub1_1_addc_out[1]}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_6895, add_sub1_1_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_6358, add_sub1_1_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_6357, add_sub1_1_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_6485, add_sub1_1_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_6172, add_sub1_1_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_6174, add_sub1_1_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_6357, add_sub1_1_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_6175, add_sub1_1_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_6004, addc_in[90]}), .c ({new_AGEMA_signal_6358, add_sub1_1_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_6169, add_sub1_1_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_6359, add_sub1_1_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_6487, subc_out[88]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_6171, add_sub1_1_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_5998, addc_in[88]}), .c ({new_AGEMA_signal_6359, add_sub1_1_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6001, addc_in[89]}), .b ({new_AGEMA_signal_6004, addc_in[90]}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_6171, add_sub1_1_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6001, addc_in[89]}), .b ({new_AGEMA_signal_6007, addc_in[91]}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_6172, add_sub1_1_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6004, addc_in[90]}), .b ({new_AGEMA_signal_6007, addc_in[91]}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_6173, add_sub1_1_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5998, addc_in[88]}), .b ({new_AGEMA_signal_6007, addc_in[91]}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_6174, add_sub1_1_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5998, addc_in[88]}), .b ({new_AGEMA_signal_6001, addc_in[89]}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_6175, add_sub1_1_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_6363, add_sub1_1_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_6362, add_sub1_1_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_6488, add_sub1_1_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_6179, add_sub1_1_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_6181, add_sub1_1_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_6362, add_sub1_1_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_6182, add_sub1_1_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_5992, addc_in[86]}), .c ({new_AGEMA_signal_6363, add_sub1_1_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_6176, add_sub1_1_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_6364, add_sub1_1_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_6490, subc_out[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_6178, add_sub1_1_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_5986, addc_in[84]}), .c ({new_AGEMA_signal_6364, add_sub1_1_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5989, addc_in[85]}), .b ({new_AGEMA_signal_5992, addc_in[86]}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_6178, add_sub1_1_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5989, addc_in[85]}), .b ({new_AGEMA_signal_5995, addc_in[87]}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_6179, add_sub1_1_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5992, addc_in[86]}), .b ({new_AGEMA_signal_5995, addc_in[87]}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_6180, add_sub1_1_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5986, addc_in[84]}), .b ({new_AGEMA_signal_5995, addc_in[87]}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_6181, add_sub1_1_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5986, addc_in[84]}), .b ({new_AGEMA_signal_5989, addc_in[85]}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_6182, add_sub1_1_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_6368, add_sub1_1_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_6367, add_sub1_1_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_6491, add_sub1_1_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_6186, add_sub1_1_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_6188, add_sub1_1_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_6367, add_sub1_1_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_6189, add_sub1_1_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_5980, addc_in[82]}), .c ({new_AGEMA_signal_6368, add_sub1_1_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_6183, add_sub1_1_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_6369, add_sub1_1_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_6493, subc_out[80]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_6185, add_sub1_1_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_5974, addc_in[80]}), .c ({new_AGEMA_signal_6369, add_sub1_1_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5977, addc_in[81]}), .b ({new_AGEMA_signal_5980, addc_in[82]}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_6185, add_sub1_1_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5977, addc_in[81]}), .b ({new_AGEMA_signal_5983, addc_in[83]}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_6186, add_sub1_1_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5980, addc_in[82]}), .b ({new_AGEMA_signal_5983, addc_in[83]}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_6187, add_sub1_1_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5974, addc_in[80]}), .b ({new_AGEMA_signal_5983, addc_in[83]}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_6188, add_sub1_1_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5974, addc_in[80]}), .b ({new_AGEMA_signal_5977, addc_in[81]}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_6189, add_sub1_1_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_6373, add_sub1_1_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_6372, add_sub1_1_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_6494, add_sub1_1_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_6193, add_sub1_1_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_6195, add_sub1_1_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_6372, add_sub1_1_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_6196, add_sub1_1_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_5968, addc_in[78]}), .c ({new_AGEMA_signal_6373, add_sub1_1_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_6190, add_sub1_1_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_6374, add_sub1_1_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_6496, subc_out[76]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_6192, add_sub1_1_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_5962, addc_in[76]}), .c ({new_AGEMA_signal_6374, add_sub1_1_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5965, addc_in[77]}), .b ({new_AGEMA_signal_5968, addc_in[78]}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_6192, add_sub1_1_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5965, addc_in[77]}), .b ({new_AGEMA_signal_5971, addc_in[79]}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_6193, add_sub1_1_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5968, addc_in[78]}), .b ({new_AGEMA_signal_5971, addc_in[79]}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_6194, add_sub1_1_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5962, addc_in[76]}), .b ({new_AGEMA_signal_5971, addc_in[79]}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_6195, add_sub1_1_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5962, addc_in[76]}), .b ({new_AGEMA_signal_5965, addc_in[77]}), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_6196, add_sub1_1_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_6378, add_sub1_1_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_6377, add_sub1_1_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_6497, add_sub1_1_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_6200, add_sub1_1_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_6202, add_sub1_1_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_6377, add_sub1_1_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_6203, add_sub1_1_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_5956, addc_in[74]}), .c ({new_AGEMA_signal_6378, add_sub1_1_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_6197, add_sub1_1_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_6379, add_sub1_1_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_6499, subc_out[72]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_6199, add_sub1_1_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_5950, addc_in[72]}), .c ({new_AGEMA_signal_6379, add_sub1_1_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5953, addc_in[73]}), .b ({new_AGEMA_signal_5956, addc_in[74]}), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_6199, add_sub1_1_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5953, addc_in[73]}), .b ({new_AGEMA_signal_5959, addc_in[75]}), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_6200, add_sub1_1_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5956, addc_in[74]}), .b ({new_AGEMA_signal_5959, addc_in[75]}), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_6201, add_sub1_1_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5950, addc_in[72]}), .b ({new_AGEMA_signal_5959, addc_in[75]}), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_6202, add_sub1_1_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5950, addc_in[72]}), .b ({new_AGEMA_signal_5953, addc_in[73]}), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_6203, add_sub1_1_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_6383, add_sub1_1_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_6382, add_sub1_1_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_6500, add_sub1_1_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_6207, add_sub1_1_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_6209, add_sub1_1_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_6382, add_sub1_1_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_6210, add_sub1_1_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_5944, addc_in[70]}), .c ({new_AGEMA_signal_6383, add_sub1_1_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_6204, add_sub1_1_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_6384, add_sub1_1_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_6502, subc_out[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_6206, add_sub1_1_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_5938, addc_in[68]}), .c ({new_AGEMA_signal_6384, add_sub1_1_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5941, addc_in[69]}), .b ({new_AGEMA_signal_5944, addc_in[70]}), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_6206, add_sub1_1_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5941, addc_in[69]}), .b ({new_AGEMA_signal_5947, addc_in[71]}), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_6207, add_sub1_1_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5944, addc_in[70]}), .b ({new_AGEMA_signal_5947, addc_in[71]}), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_6208, add_sub1_1_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5938, addc_in[68]}), .b ({new_AGEMA_signal_5947, addc_in[71]}), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_6209, add_sub1_1_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5938, addc_in[68]}), .b ({new_AGEMA_signal_5941, addc_in[69]}), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_6210, add_sub1_1_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_6388, add_sub1_1_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_6387, add_sub1_1_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_6503, add_sub1_1_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_6214, add_sub1_1_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_6216, add_sub1_1_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_6387, add_sub1_1_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_6217, add_sub1_1_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_5932, addc_in[66]}), .c ({new_AGEMA_signal_6388, add_sub1_1_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_6211, add_sub1_1_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_6389, add_sub1_1_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_6505, subc_out[64]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_6213, add_sub1_1_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_5926, addc_in[64]}), .c ({new_AGEMA_signal_6389, add_sub1_1_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5929, addc_in[65]}), .b ({new_AGEMA_signal_5932, addc_in[66]}), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_6213, add_sub1_1_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5929, addc_in[65]}), .b ({new_AGEMA_signal_5935, addc_in[67]}), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_6214, add_sub1_1_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5932, addc_in[66]}), .b ({new_AGEMA_signal_5935, addc_in[67]}), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_6215, add_sub1_1_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5926, addc_in[64]}), .b ({new_AGEMA_signal_5935, addc_in[67]}), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_6216, add_sub1_1_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5926, addc_in[64]}), .b ({new_AGEMA_signal_5929, addc_in[65]}), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_6217, add_sub1_1_subc_rom_sbox_0_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_7199, add_sub1_2_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_7198, add_sub1_2_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_7282, add_sub1_2_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_6913, add_sub1_2_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_6915, add_sub1_2_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_7198, add_sub1_2_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_6916, add_sub1_2_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_6655, add_sub1_2_addc_out[2]}), .c ({new_AGEMA_signal_7199, add_sub1_2_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_6910, add_sub1_2_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_7200, add_sub1_2_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_7284, subc_out[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_6912, add_sub1_2_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_6657, add_sub1_2_addc_out[0]}), .c ({new_AGEMA_signal_7200, add_sub1_2_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6656, add_sub1_2_addc_out[1]}), .b ({new_AGEMA_signal_6655, add_sub1_2_addc_out[2]}), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_6912, add_sub1_2_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6656, add_sub1_2_addc_out[1]}), .b ({new_AGEMA_signal_6654, add_sub1_2_addc_out[3]}), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_6913, add_sub1_2_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6655, add_sub1_2_addc_out[2]}), .b ({new_AGEMA_signal_6654, add_sub1_2_addc_out[3]}), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_6914, add_sub1_2_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6657, add_sub1_2_addc_out[0]}), .b ({new_AGEMA_signal_6654, add_sub1_2_addc_out[3]}), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_6915, add_sub1_2_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6657, add_sub1_2_addc_out[0]}), .b ({new_AGEMA_signal_6656, add_sub1_2_addc_out[1]}), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_6916, add_sub1_2_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_6394, add_sub1_2_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_6393, add_sub1_2_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_6506, add_sub1_2_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_6223, add_sub1_2_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_6225, add_sub1_2_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_6393, add_sub1_2_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_6226, add_sub1_2_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_5908, addc_in[58]}), .c ({new_AGEMA_signal_6394, add_sub1_2_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_6220, add_sub1_2_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_6395, add_sub1_2_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_6508, subc_out[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_6222, add_sub1_2_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_5902, addc_in[56]}), .c ({new_AGEMA_signal_6395, add_sub1_2_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5905, addc_in[57]}), .b ({new_AGEMA_signal_5908, addc_in[58]}), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_6222, add_sub1_2_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5905, addc_in[57]}), .b ({new_AGEMA_signal_5911, addc_in[59]}), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_6223, add_sub1_2_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5908, addc_in[58]}), .b ({new_AGEMA_signal_5911, addc_in[59]}), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_6224, add_sub1_2_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5902, addc_in[56]}), .b ({new_AGEMA_signal_5911, addc_in[59]}), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_6225, add_sub1_2_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5902, addc_in[56]}), .b ({new_AGEMA_signal_5905, addc_in[57]}), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_6226, add_sub1_2_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_6399, add_sub1_2_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_6398, add_sub1_2_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_6509, add_sub1_2_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_6230, add_sub1_2_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_6232, add_sub1_2_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_6398, add_sub1_2_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_6233, add_sub1_2_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_5896, addc_in[54]}), .c ({new_AGEMA_signal_6399, add_sub1_2_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_6227, add_sub1_2_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_6400, add_sub1_2_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_6511, subc_out[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_6229, add_sub1_2_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_5890, addc_in[52]}), .c ({new_AGEMA_signal_6400, add_sub1_2_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5893, addc_in[53]}), .b ({new_AGEMA_signal_5896, addc_in[54]}), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_6229, add_sub1_2_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5893, addc_in[53]}), .b ({new_AGEMA_signal_5899, addc_in[55]}), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_6230, add_sub1_2_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5896, addc_in[54]}), .b ({new_AGEMA_signal_5899, addc_in[55]}), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_6231, add_sub1_2_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5890, addc_in[52]}), .b ({new_AGEMA_signal_5899, addc_in[55]}), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_6232, add_sub1_2_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5890, addc_in[52]}), .b ({new_AGEMA_signal_5893, addc_in[53]}), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_6233, add_sub1_2_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_6404, add_sub1_2_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_6403, add_sub1_2_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_6512, add_sub1_2_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_6237, add_sub1_2_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_6239, add_sub1_2_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_6403, add_sub1_2_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_6240, add_sub1_2_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_5884, addc_in[50]}), .c ({new_AGEMA_signal_6404, add_sub1_2_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_6234, add_sub1_2_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_6405, add_sub1_2_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_6514, subc_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_6236, add_sub1_2_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_5878, addc_in[48]}), .c ({new_AGEMA_signal_6405, add_sub1_2_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5881, addc_in[49]}), .b ({new_AGEMA_signal_5884, addc_in[50]}), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_6236, add_sub1_2_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5881, addc_in[49]}), .b ({new_AGEMA_signal_5887, addc_in[51]}), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_6237, add_sub1_2_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5884, addc_in[50]}), .b ({new_AGEMA_signal_5887, addc_in[51]}), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_6238, add_sub1_2_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5878, addc_in[48]}), .b ({new_AGEMA_signal_5887, addc_in[51]}), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_6239, add_sub1_2_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5878, addc_in[48]}), .b ({new_AGEMA_signal_5881, addc_in[49]}), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_6240, add_sub1_2_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_6409, add_sub1_2_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_6408, add_sub1_2_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_6515, add_sub1_2_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_6244, add_sub1_2_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_6246, add_sub1_2_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_6408, add_sub1_2_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_6247, add_sub1_2_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_5872, addc_in[46]}), .c ({new_AGEMA_signal_6409, add_sub1_2_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_6241, add_sub1_2_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_6410, add_sub1_2_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_6517, subc_out[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_6243, add_sub1_2_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_5866, addc_in[44]}), .c ({new_AGEMA_signal_6410, add_sub1_2_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5869, addc_in[45]}), .b ({new_AGEMA_signal_5872, addc_in[46]}), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_6243, add_sub1_2_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5869, addc_in[45]}), .b ({new_AGEMA_signal_5875, addc_in[47]}), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_6244, add_sub1_2_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5872, addc_in[46]}), .b ({new_AGEMA_signal_5875, addc_in[47]}), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_6245, add_sub1_2_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5866, addc_in[44]}), .b ({new_AGEMA_signal_5875, addc_in[47]}), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_6246, add_sub1_2_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5866, addc_in[44]}), .b ({new_AGEMA_signal_5869, addc_in[45]}), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_6247, add_sub1_2_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_6414, add_sub1_2_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_6413, add_sub1_2_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_6518, add_sub1_2_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_6251, add_sub1_2_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_6253, add_sub1_2_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_6413, add_sub1_2_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_6254, add_sub1_2_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_5860, addc_in[42]}), .c ({new_AGEMA_signal_6414, add_sub1_2_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_6248, add_sub1_2_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_6415, add_sub1_2_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_6520, subc_out[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_6250, add_sub1_2_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_5854, addc_in[40]}), .c ({new_AGEMA_signal_6415, add_sub1_2_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5857, addc_in[41]}), .b ({new_AGEMA_signal_5860, addc_in[42]}), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_6250, add_sub1_2_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5857, addc_in[41]}), .b ({new_AGEMA_signal_5863, addc_in[43]}), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_6251, add_sub1_2_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5860, addc_in[42]}), .b ({new_AGEMA_signal_5863, addc_in[43]}), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_6252, add_sub1_2_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5854, addc_in[40]}), .b ({new_AGEMA_signal_5863, addc_in[43]}), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_6253, add_sub1_2_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5854, addc_in[40]}), .b ({new_AGEMA_signal_5857, addc_in[41]}), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_6254, add_sub1_2_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_6419, add_sub1_2_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_6418, add_sub1_2_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_6521, add_sub1_2_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_6258, add_sub1_2_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_6260, add_sub1_2_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_6418, add_sub1_2_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_6261, add_sub1_2_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_5848, addc_in[38]}), .c ({new_AGEMA_signal_6419, add_sub1_2_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_6255, add_sub1_2_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_6420, add_sub1_2_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_6523, subc_out[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_6257, add_sub1_2_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_5842, addc_in[36]}), .c ({new_AGEMA_signal_6420, add_sub1_2_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5845, addc_in[37]}), .b ({new_AGEMA_signal_5848, addc_in[38]}), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_6257, add_sub1_2_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5845, addc_in[37]}), .b ({new_AGEMA_signal_5851, addc_in[39]}), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_6258, add_sub1_2_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5848, addc_in[38]}), .b ({new_AGEMA_signal_5851, addc_in[39]}), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_6259, add_sub1_2_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5842, addc_in[36]}), .b ({new_AGEMA_signal_5851, addc_in[39]}), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_6260, add_sub1_2_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5842, addc_in[36]}), .b ({new_AGEMA_signal_5845, addc_in[37]}), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_6261, add_sub1_2_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_6424, add_sub1_2_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_6423, add_sub1_2_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_6524, add_sub1_2_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_6265, add_sub1_2_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_6267, add_sub1_2_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_6423, add_sub1_2_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_6268, add_sub1_2_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_5836, addc_in[34]}), .c ({new_AGEMA_signal_6424, add_sub1_2_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_6262, add_sub1_2_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_6425, add_sub1_2_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_6526, subc_out[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_6264, add_sub1_2_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_5830, addc_in[32]}), .c ({new_AGEMA_signal_6425, add_sub1_2_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5833, addc_in[33]}), .b ({new_AGEMA_signal_5836, addc_in[34]}), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_6264, add_sub1_2_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5833, addc_in[33]}), .b ({new_AGEMA_signal_5839, addc_in[35]}), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_6265, add_sub1_2_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5836, addc_in[34]}), .b ({new_AGEMA_signal_5839, addc_in[35]}), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_6266, add_sub1_2_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5830, addc_in[32]}), .b ({new_AGEMA_signal_5839, addc_in[35]}), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_6267, add_sub1_2_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5830, addc_in[32]}), .b ({new_AGEMA_signal_5833, addc_in[33]}), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_6268, add_sub1_2_subc_rom_sbox_0_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_7211, add_sub1_3_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_7210, add_sub1_3_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_7285, add_sub1_3_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_6934, add_sub1_3_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_6936, add_sub1_3_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_7210, add_sub1_3_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_6937, add_sub1_3_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_6666, add_sub1_3_addc_out[2]}), .c ({new_AGEMA_signal_7211, add_sub1_3_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_6931, add_sub1_3_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_7212, add_sub1_3_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_7287, subc_out[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_6933, add_sub1_3_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_6668, add_sub1_3_addc_out[0]}), .c ({new_AGEMA_signal_7212, add_sub1_3_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6667, add_sub1_3_addc_out[1]}), .b ({new_AGEMA_signal_6666, add_sub1_3_addc_out[2]}), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_6933, add_sub1_3_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6667, add_sub1_3_addc_out[1]}), .b ({new_AGEMA_signal_6665, add_sub1_3_addc_out[3]}), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_6934, add_sub1_3_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6666, add_sub1_3_addc_out[2]}), .b ({new_AGEMA_signal_6665, add_sub1_3_addc_out[3]}), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_6935, add_sub1_3_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6668, add_sub1_3_addc_out[0]}), .b ({new_AGEMA_signal_6665, add_sub1_3_addc_out[3]}), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_6936, add_sub1_3_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6668, add_sub1_3_addc_out[0]}), .b ({new_AGEMA_signal_6667, add_sub1_3_addc_out[1]}), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_6937, add_sub1_3_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_6430, add_sub1_3_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_6429, add_sub1_3_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_6527, add_sub1_3_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_6274, add_sub1_3_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_6276, add_sub1_3_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_6429, add_sub1_3_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_6277, add_sub1_3_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_5812, addc_in[26]}), .c ({new_AGEMA_signal_6430, add_sub1_3_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_6271, add_sub1_3_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_6431, add_sub1_3_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_6529, subc_out[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_6273, add_sub1_3_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_5806, addc_in[24]}), .c ({new_AGEMA_signal_6431, add_sub1_3_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5809, addc_in[25]}), .b ({new_AGEMA_signal_5812, addc_in[26]}), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_6273, add_sub1_3_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5809, addc_in[25]}), .b ({new_AGEMA_signal_5815, addc_in[27]}), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_6274, add_sub1_3_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5812, addc_in[26]}), .b ({new_AGEMA_signal_5815, addc_in[27]}), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_6275, add_sub1_3_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5806, addc_in[24]}), .b ({new_AGEMA_signal_5815, addc_in[27]}), .clk (clk), .r (Fresh[128]), .c ({new_AGEMA_signal_6276, add_sub1_3_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5806, addc_in[24]}), .b ({new_AGEMA_signal_5809, addc_in[25]}), .clk (clk), .r (Fresh[129]), .c ({new_AGEMA_signal_6277, add_sub1_3_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_6435, add_sub1_3_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_6434, add_sub1_3_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_6530, add_sub1_3_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_6281, add_sub1_3_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_6283, add_sub1_3_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_6434, add_sub1_3_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_6284, add_sub1_3_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_5800, addc_in[22]}), .c ({new_AGEMA_signal_6435, add_sub1_3_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_6278, add_sub1_3_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_6436, add_sub1_3_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_6532, subc_out[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_6280, add_sub1_3_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_5794, addc_in[20]}), .c ({new_AGEMA_signal_6436, add_sub1_3_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5797, addc_in[21]}), .b ({new_AGEMA_signal_5800, addc_in[22]}), .clk (clk), .r (Fresh[130]), .c ({new_AGEMA_signal_6280, add_sub1_3_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5797, addc_in[21]}), .b ({new_AGEMA_signal_5803, addc_in[23]}), .clk (clk), .r (Fresh[131]), .c ({new_AGEMA_signal_6281, add_sub1_3_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5800, addc_in[22]}), .b ({new_AGEMA_signal_5803, addc_in[23]}), .clk (clk), .r (Fresh[132]), .c ({new_AGEMA_signal_6282, add_sub1_3_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5794, addc_in[20]}), .b ({new_AGEMA_signal_5803, addc_in[23]}), .clk (clk), .r (Fresh[133]), .c ({new_AGEMA_signal_6283, add_sub1_3_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5794, addc_in[20]}), .b ({new_AGEMA_signal_5797, addc_in[21]}), .clk (clk), .r (Fresh[134]), .c ({new_AGEMA_signal_6284, add_sub1_3_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_6440, add_sub1_3_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_6439, add_sub1_3_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_6533, add_sub1_3_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_6288, add_sub1_3_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_6290, add_sub1_3_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_6439, add_sub1_3_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_6291, add_sub1_3_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_5788, addc_in[18]}), .c ({new_AGEMA_signal_6440, add_sub1_3_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_6285, add_sub1_3_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_6441, add_sub1_3_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_6535, subc_out[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_6287, add_sub1_3_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_5782, addc_in[16]}), .c ({new_AGEMA_signal_6441, add_sub1_3_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5785, addc_in[17]}), .b ({new_AGEMA_signal_5788, addc_in[18]}), .clk (clk), .r (Fresh[135]), .c ({new_AGEMA_signal_6287, add_sub1_3_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5785, addc_in[17]}), .b ({new_AGEMA_signal_5791, addc_in[19]}), .clk (clk), .r (Fresh[136]), .c ({new_AGEMA_signal_6288, add_sub1_3_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5788, addc_in[18]}), .b ({new_AGEMA_signal_5791, addc_in[19]}), .clk (clk), .r (Fresh[137]), .c ({new_AGEMA_signal_6289, add_sub1_3_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5782, addc_in[16]}), .b ({new_AGEMA_signal_5791, addc_in[19]}), .clk (clk), .r (Fresh[138]), .c ({new_AGEMA_signal_6290, add_sub1_3_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5782, addc_in[16]}), .b ({new_AGEMA_signal_5785, addc_in[17]}), .clk (clk), .r (Fresh[139]), .c ({new_AGEMA_signal_6291, add_sub1_3_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_6445, add_sub1_3_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_6444, add_sub1_3_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_6536, add_sub1_3_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_6295, add_sub1_3_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_6297, add_sub1_3_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_6444, add_sub1_3_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_6298, add_sub1_3_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_5776, addc_in[14]}), .c ({new_AGEMA_signal_6445, add_sub1_3_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_6292, add_sub1_3_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_6446, add_sub1_3_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_6538, subc_out[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_6294, add_sub1_3_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_5770, addc_in[12]}), .c ({new_AGEMA_signal_6446, add_sub1_3_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5773, addc_in[13]}), .b ({new_AGEMA_signal_5776, addc_in[14]}), .clk (clk), .r (Fresh[140]), .c ({new_AGEMA_signal_6294, add_sub1_3_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5773, addc_in[13]}), .b ({new_AGEMA_signal_5779, addc_in[15]}), .clk (clk), .r (Fresh[141]), .c ({new_AGEMA_signal_6295, add_sub1_3_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5776, addc_in[14]}), .b ({new_AGEMA_signal_5779, addc_in[15]}), .clk (clk), .r (Fresh[142]), .c ({new_AGEMA_signal_6296, add_sub1_3_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5770, addc_in[12]}), .b ({new_AGEMA_signal_5779, addc_in[15]}), .clk (clk), .r (Fresh[143]), .c ({new_AGEMA_signal_6297, add_sub1_3_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5770, addc_in[12]}), .b ({new_AGEMA_signal_5773, addc_in[13]}), .clk (clk), .r (Fresh[144]), .c ({new_AGEMA_signal_6298, add_sub1_3_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_6450, add_sub1_3_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_6449, add_sub1_3_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_6539, add_sub1_3_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_6302, add_sub1_3_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_6304, add_sub1_3_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_6449, add_sub1_3_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_6305, add_sub1_3_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_5764, addc_in[10]}), .c ({new_AGEMA_signal_6450, add_sub1_3_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_6299, add_sub1_3_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_6451, add_sub1_3_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_6541, subc_out[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_6301, add_sub1_3_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_5758, addc_in[8]}), .c ({new_AGEMA_signal_6451, add_sub1_3_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5761, addc_in[9]}), .b ({new_AGEMA_signal_5764, addc_in[10]}), .clk (clk), .r (Fresh[145]), .c ({new_AGEMA_signal_6301, add_sub1_3_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5761, addc_in[9]}), .b ({new_AGEMA_signal_5767, addc_in[11]}), .clk (clk), .r (Fresh[146]), .c ({new_AGEMA_signal_6302, add_sub1_3_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5764, addc_in[10]}), .b ({new_AGEMA_signal_5767, addc_in[11]}), .clk (clk), .r (Fresh[147]), .c ({new_AGEMA_signal_6303, add_sub1_3_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5758, addc_in[8]}), .b ({new_AGEMA_signal_5767, addc_in[11]}), .clk (clk), .r (Fresh[148]), .c ({new_AGEMA_signal_6304, add_sub1_3_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5758, addc_in[8]}), .b ({new_AGEMA_signal_5761, addc_in[9]}), .clk (clk), .r (Fresh[149]), .c ({new_AGEMA_signal_6305, add_sub1_3_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_6455, add_sub1_3_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_6454, add_sub1_3_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_6542, add_sub1_3_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_6309, add_sub1_3_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_6311, add_sub1_3_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_6454, add_sub1_3_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_6312, add_sub1_3_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_5752, addc_in[6]}), .c ({new_AGEMA_signal_6455, add_sub1_3_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_6306, add_sub1_3_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_6456, add_sub1_3_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_6544, subc_out[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_6308, add_sub1_3_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_5746, addc_in[4]}), .c ({new_AGEMA_signal_6456, add_sub1_3_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5749, addc_in[5]}), .b ({new_AGEMA_signal_5752, addc_in[6]}), .clk (clk), .r (Fresh[150]), .c ({new_AGEMA_signal_6308, add_sub1_3_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5749, addc_in[5]}), .b ({new_AGEMA_signal_5755, addc_in[7]}), .clk (clk), .r (Fresh[151]), .c ({new_AGEMA_signal_6309, add_sub1_3_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5752, addc_in[6]}), .b ({new_AGEMA_signal_5755, addc_in[7]}), .clk (clk), .r (Fresh[152]), .c ({new_AGEMA_signal_6310, add_sub1_3_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5746, addc_in[4]}), .b ({new_AGEMA_signal_5755, addc_in[7]}), .clk (clk), .r (Fresh[153]), .c ({new_AGEMA_signal_6311, add_sub1_3_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5746, addc_in[4]}), .b ({new_AGEMA_signal_5749, addc_in[5]}), .clk (clk), .r (Fresh[154]), .c ({new_AGEMA_signal_6312, add_sub1_3_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_6460, add_sub1_3_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_6459, add_sub1_3_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_6545, add_sub1_3_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_6316, add_sub1_3_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_6318, add_sub1_3_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_6459, add_sub1_3_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_6319, add_sub1_3_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_5740, addc_in[2]}), .c ({new_AGEMA_signal_6460, add_sub1_3_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_6313, add_sub1_3_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_6461, add_sub1_3_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_6547, subc_out[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_6315, add_sub1_3_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_5734, addc_in[0]}), .c ({new_AGEMA_signal_6461, add_sub1_3_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5737, addc_in[1]}), .b ({new_AGEMA_signal_5740, addc_in[2]}), .clk (clk), .r (Fresh[155]), .c ({new_AGEMA_signal_6315, add_sub1_3_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5737, addc_in[1]}), .b ({new_AGEMA_signal_5743, addc_in[3]}), .clk (clk), .r (Fresh[156]), .c ({new_AGEMA_signal_6316, add_sub1_3_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5740, addc_in[2]}), .b ({new_AGEMA_signal_5743, addc_in[3]}), .clk (clk), .r (Fresh[157]), .c ({new_AGEMA_signal_6317, add_sub1_3_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5734, addc_in[0]}), .b ({new_AGEMA_signal_5743, addc_in[3]}), .clk (clk), .r (Fresh[158]), .c ({new_AGEMA_signal_6318, add_sub1_3_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5734, addc_in[0]}), .b ({new_AGEMA_signal_5737, addc_in[1]}), .clk (clk), .r (Fresh[159]), .c ({new_AGEMA_signal_6319, add_sub1_3_subc_rom_sbox_0_ANF_2_t7}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6484, subc_out[96]}), .a ({new_AGEMA_signal_6472, subc_out[112]}), .c ({new_AGEMA_signal_6608, shiftr_out[96]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6481, subc_out[100]}), .a ({new_AGEMA_signal_6469, subc_out[116]}), .c ({new_AGEMA_signal_6609, shiftr_out[100]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6478, subc_out[104]}), .a ({new_AGEMA_signal_6466, subc_out[120]}), .c ({new_AGEMA_signal_6610, shiftr_out[104]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6475, subc_out[108]}), .a ({new_AGEMA_signal_7278, subc_out[124]}), .c ({new_AGEMA_signal_7614, shiftr_out[108]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6472, subc_out[112]}), .a ({new_AGEMA_signal_6484, subc_out[96]}), .c ({new_AGEMA_signal_6611, shiftr_out[112]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6469, subc_out[116]}), .a ({new_AGEMA_signal_6481, subc_out[100]}), .c ({new_AGEMA_signal_6612, shiftr_out[116]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6466, subc_out[120]}), .a ({new_AGEMA_signal_6478, subc_out[104]}), .c ({new_AGEMA_signal_6613, shiftr_out[120]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7278, subc_out[124]}), .a ({new_AGEMA_signal_6475, subc_out[108]}), .c ({new_AGEMA_signal_7615, shiftr_out[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7281, subc_out[92]}), .a ({new_AGEMA_signal_6496, subc_out[76]}), .c ({new_AGEMA_signal_7616, shiftr_out[64]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6505, subc_out[64]}), .a ({new_AGEMA_signal_6493, subc_out[80]}), .c ({new_AGEMA_signal_6614, shiftr_out[68]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6502, subc_out[68]}), .a ({new_AGEMA_signal_6490, subc_out[84]}), .c ({new_AGEMA_signal_6615, shiftr_out[72]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6499, subc_out[72]}), .a ({new_AGEMA_signal_6487, subc_out[88]}), .c ({new_AGEMA_signal_6616, shiftr_out[76]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6496, subc_out[76]}), .a ({new_AGEMA_signal_7281, subc_out[92]}), .c ({new_AGEMA_signal_7617, shiftr_out[80]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6493, subc_out[80]}), .a ({new_AGEMA_signal_6505, subc_out[64]}), .c ({new_AGEMA_signal_6617, shiftr_out[84]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6490, subc_out[84]}), .a ({new_AGEMA_signal_6502, subc_out[68]}), .c ({new_AGEMA_signal_6618, shiftr_out[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6487, subc_out[88]}), .a ({new_AGEMA_signal_6499, subc_out[72]}), .c ({new_AGEMA_signal_6619, shiftr_out[92]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6508, subc_out[56]}), .a ({new_AGEMA_signal_6520, subc_out[40]}), .c ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7284, subc_out[60]}), .a ({new_AGEMA_signal_6517, subc_out[44]}), .c ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6526, subc_out[32]}), .a ({new_AGEMA_signal_6514, subc_out[48]}), .c ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6523, subc_out[36]}), .a ({new_AGEMA_signal_6511, subc_out[52]}), .c ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6520, subc_out[40]}), .a ({new_AGEMA_signal_6508, subc_out[56]}), .c ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6517, subc_out[44]}), .a ({new_AGEMA_signal_7284, subc_out[60]}), .c ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6514, subc_out[48]}), .a ({new_AGEMA_signal_6526, subc_out[32]}), .c ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6511, subc_out[52]}), .a ({new_AGEMA_signal_6523, subc_out[36]}), .c ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6532, subc_out[20]}), .a ({new_AGEMA_signal_6544, subc_out[4]}), .c ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6529, subc_out[24]}), .a ({new_AGEMA_signal_6541, subc_out[8]}), .c ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7287, subc_out[28]}), .a ({new_AGEMA_signal_6538, subc_out[12]}), .c ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6547, subc_out[0]}), .a ({new_AGEMA_signal_6535, subc_out[16]}), .c ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6544, subc_out[4]}), .a ({new_AGEMA_signal_6532, subc_out[20]}), .c ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6541, subc_out[8]}), .a ({new_AGEMA_signal_6529, subc_out[24]}), .c ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6538, subc_out[12]}), .a ({new_AGEMA_signal_7287, subc_out[28]}), .c ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6535, subc_out[16]}), .a ({new_AGEMA_signal_6547, subc_out[0]}), .c ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_8090, add_sub1_0_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_7176, add_sub1_0_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_8572, subc_out[127]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_7277, add_sub1_0_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_7276, add_sub1_0_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_7606, subc_out[126]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_8573, add_sub1_0_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_6872, add_sub1_0_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_9048, subc_out[125]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_8090, add_sub1_0_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_6871, add_sub1_0_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_8573, add_sub1_0_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_7607, add_sub1_0_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_6634, add_sub1_0_addc_out[1]}), .c ({new_AGEMA_signal_8090, add_sub1_0_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_7277, add_sub1_0_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_7177, add_sub1_0_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_7607, add_sub1_0_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_7178, add_sub1_0_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_6632, add_sub1_0_addc_out[3]}), .c ({new_AGEMA_signal_7277, add_sub1_0_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6635, add_sub1_0_addc_out[0]}), .b ({new_AGEMA_signal_6870, add_sub1_0_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r (Fresh[160]), .c ({new_AGEMA_signal_7177, add_sub1_0_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6869, add_sub1_0_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_6873, add_sub1_0_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r (Fresh[161]), .c ({new_AGEMA_signal_7178, add_sub1_0_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_6636, add_sub1_0_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6323, add_sub1_0_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_6875, subc_out[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_6465, add_sub1_0_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_6464, add_sub1_0_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_6549, subc_out[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_6876, add_sub1_0_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_6122, add_sub1_0_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_7179, subc_out[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_6636, add_sub1_0_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6121, add_sub1_0_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_6876, add_sub1_0_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_6550, add_sub1_0_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_6097, addc_in[121]}), .c ({new_AGEMA_signal_6636, add_sub1_0_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_6465, add_sub1_0_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_6324, add_sub1_0_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_6550, add_sub1_0_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_6325, add_sub1_0_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_6103, addc_in[123]}), .c ({new_AGEMA_signal_6465, add_sub1_0_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6094, addc_in[120]}), .b ({new_AGEMA_signal_6120, add_sub1_0_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r (Fresh[162]), .c ({new_AGEMA_signal_6324, add_sub1_0_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6119, add_sub1_0_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_6123, add_sub1_0_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r (Fresh[163]), .c ({new_AGEMA_signal_6325, add_sub1_0_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_6637, add_sub1_0_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6328, add_sub1_0_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_6877, subc_out[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_6468, add_sub1_0_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_6467, add_sub1_0_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_6551, subc_out[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_6878, add_sub1_0_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_6129, add_sub1_0_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_7180, subc_out[117]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_6637, add_sub1_0_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6128, add_sub1_0_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_6878, add_sub1_0_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_6552, add_sub1_0_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_6085, addc_in[117]}), .c ({new_AGEMA_signal_6637, add_sub1_0_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_6468, add_sub1_0_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_6329, add_sub1_0_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_6552, add_sub1_0_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_6330, add_sub1_0_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_6091, addc_in[119]}), .c ({new_AGEMA_signal_6468, add_sub1_0_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6082, addc_in[116]}), .b ({new_AGEMA_signal_6127, add_sub1_0_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r (Fresh[164]), .c ({new_AGEMA_signal_6329, add_sub1_0_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6126, add_sub1_0_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_6130, add_sub1_0_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r (Fresh[165]), .c ({new_AGEMA_signal_6330, add_sub1_0_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_6638, add_sub1_0_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6333, add_sub1_0_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_6879, subc_out[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_6471, add_sub1_0_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_6470, add_sub1_0_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_6553, subc_out[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_6880, add_sub1_0_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_6136, add_sub1_0_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_7181, subc_out[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_6638, add_sub1_0_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6135, add_sub1_0_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_6880, add_sub1_0_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_6554, add_sub1_0_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_6073, addc_in[113]}), .c ({new_AGEMA_signal_6638, add_sub1_0_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_6471, add_sub1_0_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_6334, add_sub1_0_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_6554, add_sub1_0_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_6335, add_sub1_0_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_6079, addc_in[115]}), .c ({new_AGEMA_signal_6471, add_sub1_0_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6070, addc_in[112]}), .b ({new_AGEMA_signal_6134, add_sub1_0_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r (Fresh[166]), .c ({new_AGEMA_signal_6334, add_sub1_0_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6133, add_sub1_0_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_6137, add_sub1_0_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r (Fresh[167]), .c ({new_AGEMA_signal_6335, add_sub1_0_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_6639, add_sub1_0_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6338, add_sub1_0_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_6881, subc_out[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_6474, add_sub1_0_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_6473, add_sub1_0_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_6555, subc_out[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_6882, add_sub1_0_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_6143, add_sub1_0_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_7182, subc_out[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_6639, add_sub1_0_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6142, add_sub1_0_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_6882, add_sub1_0_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_6556, add_sub1_0_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_6061, addc_in[109]}), .c ({new_AGEMA_signal_6639, add_sub1_0_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_6474, add_sub1_0_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_6339, add_sub1_0_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_6556, add_sub1_0_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_6340, add_sub1_0_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_6067, addc_in[111]}), .c ({new_AGEMA_signal_6474, add_sub1_0_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6058, addc_in[108]}), .b ({new_AGEMA_signal_6141, add_sub1_0_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r (Fresh[168]), .c ({new_AGEMA_signal_6339, add_sub1_0_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6140, add_sub1_0_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_6144, add_sub1_0_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r (Fresh[169]), .c ({new_AGEMA_signal_6340, add_sub1_0_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_6640, add_sub1_0_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6343, add_sub1_0_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_6883, subc_out[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_6477, add_sub1_0_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_6476, add_sub1_0_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_6557, subc_out[106]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_6884, add_sub1_0_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_6150, add_sub1_0_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_7183, subc_out[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_6640, add_sub1_0_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6149, add_sub1_0_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_6884, add_sub1_0_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_6558, add_sub1_0_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_6049, addc_in[105]}), .c ({new_AGEMA_signal_6640, add_sub1_0_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_6477, add_sub1_0_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_6344, add_sub1_0_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_6558, add_sub1_0_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_6345, add_sub1_0_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_6055, addc_in[107]}), .c ({new_AGEMA_signal_6477, add_sub1_0_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6046, addc_in[104]}), .b ({new_AGEMA_signal_6148, add_sub1_0_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r (Fresh[170]), .c ({new_AGEMA_signal_6344, add_sub1_0_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6147, add_sub1_0_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_6151, add_sub1_0_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r (Fresh[171]), .c ({new_AGEMA_signal_6345, add_sub1_0_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_6641, add_sub1_0_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6348, add_sub1_0_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_6885, subc_out[103]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_6480, add_sub1_0_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_6479, add_sub1_0_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_6559, subc_out[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_6886, add_sub1_0_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_6157, add_sub1_0_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_7184, subc_out[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_6641, add_sub1_0_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6156, add_sub1_0_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_6886, add_sub1_0_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_6560, add_sub1_0_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_6037, addc_in[101]}), .c ({new_AGEMA_signal_6641, add_sub1_0_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_6480, add_sub1_0_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_6349, add_sub1_0_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_6560, add_sub1_0_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_6350, add_sub1_0_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_6043, addc_in[103]}), .c ({new_AGEMA_signal_6480, add_sub1_0_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6034, addc_in[100]}), .b ({new_AGEMA_signal_6155, add_sub1_0_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r (Fresh[172]), .c ({new_AGEMA_signal_6349, add_sub1_0_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6154, add_sub1_0_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_6158, add_sub1_0_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r (Fresh[173]), .c ({new_AGEMA_signal_6350, add_sub1_0_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_6642, add_sub1_0_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6353, add_sub1_0_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_6887, subc_out[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_6483, add_sub1_0_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_6482, add_sub1_0_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_6561, subc_out[98]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_6888, add_sub1_0_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_6164, add_sub1_0_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_7185, subc_out[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_6642, add_sub1_0_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6163, add_sub1_0_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_6888, add_sub1_0_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_6562, add_sub1_0_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_6025, addc_in[97]}), .c ({new_AGEMA_signal_6642, add_sub1_0_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_6483, add_sub1_0_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_6354, add_sub1_0_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_6562, add_sub1_0_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_6355, add_sub1_0_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_6031, addc_in[99]}), .c ({new_AGEMA_signal_6483, add_sub1_0_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6022, addc_in[96]}), .b ({new_AGEMA_signal_6162, add_sub1_0_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r (Fresh[174]), .c ({new_AGEMA_signal_6354, add_sub1_0_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6161, add_sub1_0_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_6165, add_sub1_0_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r (Fresh[175]), .c ({new_AGEMA_signal_6355, add_sub1_0_subc_rom_sbox_0_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_8091, add_sub1_1_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_7188, add_sub1_1_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_8574, subc_out[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_7280, add_sub1_1_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_7279, add_sub1_1_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_7608, subc_out[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_8575, add_sub1_1_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_6893, add_sub1_1_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_9049, subc_out[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_8091, add_sub1_1_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_6892, add_sub1_1_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_8575, add_sub1_1_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_7609, add_sub1_1_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_6645, add_sub1_1_addc_out[1]}), .c ({new_AGEMA_signal_8091, add_sub1_1_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_7280, add_sub1_1_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_7189, add_sub1_1_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_7609, add_sub1_1_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_7190, add_sub1_1_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_6643, add_sub1_1_addc_out[3]}), .c ({new_AGEMA_signal_7280, add_sub1_1_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6646, add_sub1_1_addc_out[0]}), .b ({new_AGEMA_signal_6891, add_sub1_1_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r (Fresh[176]), .c ({new_AGEMA_signal_7189, add_sub1_1_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6890, add_sub1_1_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_6894, add_sub1_1_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r (Fresh[177]), .c ({new_AGEMA_signal_7190, add_sub1_1_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_6647, add_sub1_1_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6359, add_sub1_1_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_6896, subc_out[91]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_6486, add_sub1_1_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_6485, add_sub1_1_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_6564, subc_out[90]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_6897, add_sub1_1_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_6173, add_sub1_1_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_7191, subc_out[89]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_6647, add_sub1_1_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6172, add_sub1_1_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_6897, add_sub1_1_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_6565, add_sub1_1_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_6001, addc_in[89]}), .c ({new_AGEMA_signal_6647, add_sub1_1_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_6486, add_sub1_1_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_6360, add_sub1_1_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_6565, add_sub1_1_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_6361, add_sub1_1_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_6007, addc_in[91]}), .c ({new_AGEMA_signal_6486, add_sub1_1_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5998, addc_in[88]}), .b ({new_AGEMA_signal_6171, add_sub1_1_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r (Fresh[178]), .c ({new_AGEMA_signal_6360, add_sub1_1_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6170, add_sub1_1_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_6174, add_sub1_1_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r (Fresh[179]), .c ({new_AGEMA_signal_6361, add_sub1_1_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_6648, add_sub1_1_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6364, add_sub1_1_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_6898, subc_out[87]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_6489, add_sub1_1_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_6488, add_sub1_1_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_6566, subc_out[86]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_6899, add_sub1_1_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_6180, add_sub1_1_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_7192, subc_out[85]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_6648, add_sub1_1_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6179, add_sub1_1_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_6899, add_sub1_1_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_6567, add_sub1_1_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_5989, addc_in[85]}), .c ({new_AGEMA_signal_6648, add_sub1_1_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_6489, add_sub1_1_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_6365, add_sub1_1_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_6567, add_sub1_1_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_6366, add_sub1_1_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_5995, addc_in[87]}), .c ({new_AGEMA_signal_6489, add_sub1_1_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5986, addc_in[84]}), .b ({new_AGEMA_signal_6178, add_sub1_1_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r (Fresh[180]), .c ({new_AGEMA_signal_6365, add_sub1_1_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6177, add_sub1_1_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_6181, add_sub1_1_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r (Fresh[181]), .c ({new_AGEMA_signal_6366, add_sub1_1_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_6649, add_sub1_1_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6369, add_sub1_1_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_6900, subc_out[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_6492, add_sub1_1_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_6491, add_sub1_1_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_6568, subc_out[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_6901, add_sub1_1_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_6187, add_sub1_1_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_7193, subc_out[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_6649, add_sub1_1_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6186, add_sub1_1_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_6901, add_sub1_1_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_6569, add_sub1_1_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_5977, addc_in[81]}), .c ({new_AGEMA_signal_6649, add_sub1_1_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_6492, add_sub1_1_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_6370, add_sub1_1_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_6569, add_sub1_1_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_6371, add_sub1_1_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_5983, addc_in[83]}), .c ({new_AGEMA_signal_6492, add_sub1_1_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5974, addc_in[80]}), .b ({new_AGEMA_signal_6185, add_sub1_1_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r (Fresh[182]), .c ({new_AGEMA_signal_6370, add_sub1_1_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6184, add_sub1_1_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_6188, add_sub1_1_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r (Fresh[183]), .c ({new_AGEMA_signal_6371, add_sub1_1_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_6650, add_sub1_1_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6374, add_sub1_1_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_6902, subc_out[79]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_6495, add_sub1_1_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_6494, add_sub1_1_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_6570, subc_out[78]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_6903, add_sub1_1_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_6194, add_sub1_1_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_7194, subc_out[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_6650, add_sub1_1_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6193, add_sub1_1_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_6903, add_sub1_1_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_6571, add_sub1_1_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_5965, addc_in[77]}), .c ({new_AGEMA_signal_6650, add_sub1_1_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_6495, add_sub1_1_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_6375, add_sub1_1_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_6571, add_sub1_1_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_6376, add_sub1_1_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_5971, addc_in[79]}), .c ({new_AGEMA_signal_6495, add_sub1_1_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5962, addc_in[76]}), .b ({new_AGEMA_signal_6192, add_sub1_1_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r (Fresh[184]), .c ({new_AGEMA_signal_6375, add_sub1_1_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6191, add_sub1_1_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_6195, add_sub1_1_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r (Fresh[185]), .c ({new_AGEMA_signal_6376, add_sub1_1_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_6651, add_sub1_1_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6379, add_sub1_1_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_6904, subc_out[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_6498, add_sub1_1_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_6497, add_sub1_1_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_6572, subc_out[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_6905, add_sub1_1_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_6201, add_sub1_1_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_7195, subc_out[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_6651, add_sub1_1_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6200, add_sub1_1_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_6905, add_sub1_1_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_6573, add_sub1_1_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_5953, addc_in[73]}), .c ({new_AGEMA_signal_6651, add_sub1_1_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_6498, add_sub1_1_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_6380, add_sub1_1_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_6573, add_sub1_1_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_6381, add_sub1_1_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_5959, addc_in[75]}), .c ({new_AGEMA_signal_6498, add_sub1_1_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5950, addc_in[72]}), .b ({new_AGEMA_signal_6199, add_sub1_1_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r (Fresh[186]), .c ({new_AGEMA_signal_6380, add_sub1_1_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6198, add_sub1_1_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_6202, add_sub1_1_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r (Fresh[187]), .c ({new_AGEMA_signal_6381, add_sub1_1_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_6652, add_sub1_1_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6384, add_sub1_1_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_6906, subc_out[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_6501, add_sub1_1_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_6500, add_sub1_1_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_6574, subc_out[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_6907, add_sub1_1_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_6208, add_sub1_1_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_7196, subc_out[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_6652, add_sub1_1_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6207, add_sub1_1_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_6907, add_sub1_1_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_6575, add_sub1_1_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_5941, addc_in[69]}), .c ({new_AGEMA_signal_6652, add_sub1_1_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_6501, add_sub1_1_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_6385, add_sub1_1_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_6575, add_sub1_1_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_6386, add_sub1_1_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_5947, addc_in[71]}), .c ({new_AGEMA_signal_6501, add_sub1_1_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5938, addc_in[68]}), .b ({new_AGEMA_signal_6206, add_sub1_1_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r (Fresh[188]), .c ({new_AGEMA_signal_6385, add_sub1_1_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6205, add_sub1_1_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_6209, add_sub1_1_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r (Fresh[189]), .c ({new_AGEMA_signal_6386, add_sub1_1_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_6653, add_sub1_1_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6389, add_sub1_1_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_6908, subc_out[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_6504, add_sub1_1_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_6503, add_sub1_1_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_6576, subc_out[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_6909, add_sub1_1_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_6215, add_sub1_1_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_7197, subc_out[65]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_6653, add_sub1_1_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6214, add_sub1_1_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_6909, add_sub1_1_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_6577, add_sub1_1_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_5929, addc_in[65]}), .c ({new_AGEMA_signal_6653, add_sub1_1_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_6504, add_sub1_1_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_6390, add_sub1_1_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_6577, add_sub1_1_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_6391, add_sub1_1_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_5935, addc_in[67]}), .c ({new_AGEMA_signal_6504, add_sub1_1_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5926, addc_in[64]}), .b ({new_AGEMA_signal_6213, add_sub1_1_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r (Fresh[190]), .c ({new_AGEMA_signal_6390, add_sub1_1_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6212, add_sub1_1_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_6216, add_sub1_1_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r (Fresh[191]), .c ({new_AGEMA_signal_6391, add_sub1_1_subc_rom_sbox_0_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_8092, add_sub1_2_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_7200, add_sub1_2_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_8576, subc_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_7283, add_sub1_2_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_7282, add_sub1_2_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_7610, subc_out[62]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_8577, add_sub1_2_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_6914, add_sub1_2_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_9050, subc_out[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_8092, add_sub1_2_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_6913, add_sub1_2_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_8577, add_sub1_2_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_7611, add_sub1_2_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_6656, add_sub1_2_addc_out[1]}), .c ({new_AGEMA_signal_8092, add_sub1_2_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_7283, add_sub1_2_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_7201, add_sub1_2_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_7611, add_sub1_2_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_7202, add_sub1_2_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_6654, add_sub1_2_addc_out[3]}), .c ({new_AGEMA_signal_7283, add_sub1_2_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6657, add_sub1_2_addc_out[0]}), .b ({new_AGEMA_signal_6912, add_sub1_2_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r (Fresh[192]), .c ({new_AGEMA_signal_7201, add_sub1_2_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6911, add_sub1_2_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_6915, add_sub1_2_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r (Fresh[193]), .c ({new_AGEMA_signal_7202, add_sub1_2_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_6658, add_sub1_2_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6395, add_sub1_2_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_6917, subc_out[59]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_6507, add_sub1_2_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_6506, add_sub1_2_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_6579, subc_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_6918, add_sub1_2_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_6224, add_sub1_2_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_7203, subc_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_6658, add_sub1_2_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6223, add_sub1_2_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_6918, add_sub1_2_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_6580, add_sub1_2_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_5905, addc_in[57]}), .c ({new_AGEMA_signal_6658, add_sub1_2_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_6507, add_sub1_2_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_6396, add_sub1_2_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_6580, add_sub1_2_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_6397, add_sub1_2_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_5911, addc_in[59]}), .c ({new_AGEMA_signal_6507, add_sub1_2_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5902, addc_in[56]}), .b ({new_AGEMA_signal_6222, add_sub1_2_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r (Fresh[194]), .c ({new_AGEMA_signal_6396, add_sub1_2_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6221, add_sub1_2_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_6225, add_sub1_2_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r (Fresh[195]), .c ({new_AGEMA_signal_6397, add_sub1_2_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_6659, add_sub1_2_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6400, add_sub1_2_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_6919, subc_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_6510, add_sub1_2_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_6509, add_sub1_2_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_6581, subc_out[54]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_6920, add_sub1_2_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_6231, add_sub1_2_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_7204, subc_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_6659, add_sub1_2_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6230, add_sub1_2_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_6920, add_sub1_2_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_6582, add_sub1_2_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_5893, addc_in[53]}), .c ({new_AGEMA_signal_6659, add_sub1_2_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_6510, add_sub1_2_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_6401, add_sub1_2_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_6582, add_sub1_2_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_6402, add_sub1_2_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_5899, addc_in[55]}), .c ({new_AGEMA_signal_6510, add_sub1_2_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5890, addc_in[52]}), .b ({new_AGEMA_signal_6229, add_sub1_2_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r (Fresh[196]), .c ({new_AGEMA_signal_6401, add_sub1_2_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6228, add_sub1_2_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_6232, add_sub1_2_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r (Fresh[197]), .c ({new_AGEMA_signal_6402, add_sub1_2_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_6660, add_sub1_2_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6405, add_sub1_2_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_6921, subc_out[51]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_6513, add_sub1_2_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_6512, add_sub1_2_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_6583, subc_out[50]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_6922, add_sub1_2_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_6238, add_sub1_2_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_7205, subc_out[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_6660, add_sub1_2_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6237, add_sub1_2_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_6922, add_sub1_2_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_6584, add_sub1_2_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_5881, addc_in[49]}), .c ({new_AGEMA_signal_6660, add_sub1_2_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_6513, add_sub1_2_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_6406, add_sub1_2_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_6584, add_sub1_2_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_6407, add_sub1_2_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_5887, addc_in[51]}), .c ({new_AGEMA_signal_6513, add_sub1_2_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5878, addc_in[48]}), .b ({new_AGEMA_signal_6236, add_sub1_2_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r (Fresh[198]), .c ({new_AGEMA_signal_6406, add_sub1_2_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6235, add_sub1_2_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_6239, add_sub1_2_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r (Fresh[199]), .c ({new_AGEMA_signal_6407, add_sub1_2_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_6661, add_sub1_2_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6410, add_sub1_2_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_6923, subc_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_6516, add_sub1_2_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_6515, add_sub1_2_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_6585, subc_out[46]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_6924, add_sub1_2_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_6245, add_sub1_2_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_7206, subc_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_6661, add_sub1_2_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6244, add_sub1_2_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_6924, add_sub1_2_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_6586, add_sub1_2_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_5869, addc_in[45]}), .c ({new_AGEMA_signal_6661, add_sub1_2_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_6516, add_sub1_2_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_6411, add_sub1_2_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_6586, add_sub1_2_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_6412, add_sub1_2_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_5875, addc_in[47]}), .c ({new_AGEMA_signal_6516, add_sub1_2_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5866, addc_in[44]}), .b ({new_AGEMA_signal_6243, add_sub1_2_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r (Fresh[200]), .c ({new_AGEMA_signal_6411, add_sub1_2_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6242, add_sub1_2_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_6246, add_sub1_2_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r (Fresh[201]), .c ({new_AGEMA_signal_6412, add_sub1_2_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_6662, add_sub1_2_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6415, add_sub1_2_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_6925, subc_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_6519, add_sub1_2_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_6518, add_sub1_2_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_6587, subc_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_6926, add_sub1_2_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_6252, add_sub1_2_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_7207, subc_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_6662, add_sub1_2_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6251, add_sub1_2_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_6926, add_sub1_2_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_6588, add_sub1_2_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_5857, addc_in[41]}), .c ({new_AGEMA_signal_6662, add_sub1_2_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_6519, add_sub1_2_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_6416, add_sub1_2_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_6588, add_sub1_2_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_6417, add_sub1_2_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_5863, addc_in[43]}), .c ({new_AGEMA_signal_6519, add_sub1_2_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5854, addc_in[40]}), .b ({new_AGEMA_signal_6250, add_sub1_2_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r (Fresh[202]), .c ({new_AGEMA_signal_6416, add_sub1_2_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6249, add_sub1_2_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_6253, add_sub1_2_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r (Fresh[203]), .c ({new_AGEMA_signal_6417, add_sub1_2_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_6663, add_sub1_2_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6420, add_sub1_2_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_6927, subc_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_6522, add_sub1_2_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_6521, add_sub1_2_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_6589, subc_out[38]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_6928, add_sub1_2_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_6259, add_sub1_2_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_7208, subc_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_6663, add_sub1_2_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6258, add_sub1_2_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_6928, add_sub1_2_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_6590, add_sub1_2_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_5845, addc_in[37]}), .c ({new_AGEMA_signal_6663, add_sub1_2_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_6522, add_sub1_2_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_6421, add_sub1_2_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_6590, add_sub1_2_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_6422, add_sub1_2_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_5851, addc_in[39]}), .c ({new_AGEMA_signal_6522, add_sub1_2_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5842, addc_in[36]}), .b ({new_AGEMA_signal_6257, add_sub1_2_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r (Fresh[204]), .c ({new_AGEMA_signal_6421, add_sub1_2_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6256, add_sub1_2_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_6260, add_sub1_2_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r (Fresh[205]), .c ({new_AGEMA_signal_6422, add_sub1_2_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_6664, add_sub1_2_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6425, add_sub1_2_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_6929, subc_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_6525, add_sub1_2_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_6524, add_sub1_2_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_6591, subc_out[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_6930, add_sub1_2_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_6266, add_sub1_2_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_7209, subc_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_6664, add_sub1_2_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6265, add_sub1_2_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_6930, add_sub1_2_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_6592, add_sub1_2_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_5833, addc_in[33]}), .c ({new_AGEMA_signal_6664, add_sub1_2_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_6525, add_sub1_2_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_6426, add_sub1_2_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_6592, add_sub1_2_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_6427, add_sub1_2_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_5839, addc_in[35]}), .c ({new_AGEMA_signal_6525, add_sub1_2_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5830, addc_in[32]}), .b ({new_AGEMA_signal_6264, add_sub1_2_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r (Fresh[206]), .c ({new_AGEMA_signal_6426, add_sub1_2_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6263, add_sub1_2_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_6267, add_sub1_2_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r (Fresh[207]), .c ({new_AGEMA_signal_6427, add_sub1_2_subc_rom_sbox_0_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_8093, add_sub1_3_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_7212, add_sub1_3_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_8578, subc_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_7286, add_sub1_3_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_7285, add_sub1_3_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_7612, subc_out[30]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_8579, add_sub1_3_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_6935, add_sub1_3_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_9051, subc_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_8093, add_sub1_3_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_6934, add_sub1_3_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_8579, add_sub1_3_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_7613, add_sub1_3_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_6667, add_sub1_3_addc_out[1]}), .c ({new_AGEMA_signal_8093, add_sub1_3_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_7286, add_sub1_3_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_7213, add_sub1_3_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_7613, add_sub1_3_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_7214, add_sub1_3_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_6665, add_sub1_3_addc_out[3]}), .c ({new_AGEMA_signal_7286, add_sub1_3_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6668, add_sub1_3_addc_out[0]}), .b ({new_AGEMA_signal_6933, add_sub1_3_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r (Fresh[208]), .c ({new_AGEMA_signal_7213, add_sub1_3_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6932, add_sub1_3_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_6936, add_sub1_3_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r (Fresh[209]), .c ({new_AGEMA_signal_7214, add_sub1_3_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_6669, add_sub1_3_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6431, add_sub1_3_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_6938, subc_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_6528, add_sub1_3_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_6527, add_sub1_3_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_6594, subc_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_6939, add_sub1_3_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_6275, add_sub1_3_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_7215, subc_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_6669, add_sub1_3_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6274, add_sub1_3_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_6939, add_sub1_3_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_6595, add_sub1_3_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_5809, addc_in[25]}), .c ({new_AGEMA_signal_6669, add_sub1_3_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_6528, add_sub1_3_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_6432, add_sub1_3_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_6595, add_sub1_3_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_6433, add_sub1_3_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_5815, addc_in[27]}), .c ({new_AGEMA_signal_6528, add_sub1_3_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5806, addc_in[24]}), .b ({new_AGEMA_signal_6273, add_sub1_3_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r (Fresh[210]), .c ({new_AGEMA_signal_6432, add_sub1_3_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6272, add_sub1_3_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_6276, add_sub1_3_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r (Fresh[211]), .c ({new_AGEMA_signal_6433, add_sub1_3_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_6670, add_sub1_3_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6436, add_sub1_3_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_6940, subc_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_6531, add_sub1_3_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_6530, add_sub1_3_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_6596, subc_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_6941, add_sub1_3_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_6282, add_sub1_3_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_7216, subc_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_6670, add_sub1_3_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6281, add_sub1_3_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_6941, add_sub1_3_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_6597, add_sub1_3_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_5797, addc_in[21]}), .c ({new_AGEMA_signal_6670, add_sub1_3_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_6531, add_sub1_3_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_6437, add_sub1_3_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_6597, add_sub1_3_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_6438, add_sub1_3_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_5803, addc_in[23]}), .c ({new_AGEMA_signal_6531, add_sub1_3_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5794, addc_in[20]}), .b ({new_AGEMA_signal_6280, add_sub1_3_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r (Fresh[212]), .c ({new_AGEMA_signal_6437, add_sub1_3_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6279, add_sub1_3_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_6283, add_sub1_3_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r (Fresh[213]), .c ({new_AGEMA_signal_6438, add_sub1_3_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_6671, add_sub1_3_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6441, add_sub1_3_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_6942, subc_out[19]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_6534, add_sub1_3_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_6533, add_sub1_3_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_6598, subc_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_6943, add_sub1_3_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_6289, add_sub1_3_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_7217, subc_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_6671, add_sub1_3_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6288, add_sub1_3_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_6943, add_sub1_3_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_6599, add_sub1_3_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_5785, addc_in[17]}), .c ({new_AGEMA_signal_6671, add_sub1_3_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_6534, add_sub1_3_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_6442, add_sub1_3_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_6599, add_sub1_3_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_6443, add_sub1_3_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_5791, addc_in[19]}), .c ({new_AGEMA_signal_6534, add_sub1_3_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5782, addc_in[16]}), .b ({new_AGEMA_signal_6287, add_sub1_3_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r (Fresh[214]), .c ({new_AGEMA_signal_6442, add_sub1_3_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6286, add_sub1_3_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_6290, add_sub1_3_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r (Fresh[215]), .c ({new_AGEMA_signal_6443, add_sub1_3_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_6672, add_sub1_3_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6446, add_sub1_3_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_6944, subc_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_6537, add_sub1_3_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_6536, add_sub1_3_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_6600, subc_out[14]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_6945, add_sub1_3_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_6296, add_sub1_3_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_7218, subc_out[13]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_6672, add_sub1_3_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6295, add_sub1_3_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_6945, add_sub1_3_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_6601, add_sub1_3_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_5773, addc_in[13]}), .c ({new_AGEMA_signal_6672, add_sub1_3_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_6537, add_sub1_3_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_6447, add_sub1_3_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_6601, add_sub1_3_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_6448, add_sub1_3_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_5779, addc_in[15]}), .c ({new_AGEMA_signal_6537, add_sub1_3_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5770, addc_in[12]}), .b ({new_AGEMA_signal_6294, add_sub1_3_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r (Fresh[216]), .c ({new_AGEMA_signal_6447, add_sub1_3_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6293, add_sub1_3_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_6297, add_sub1_3_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r (Fresh[217]), .c ({new_AGEMA_signal_6448, add_sub1_3_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_6673, add_sub1_3_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6451, add_sub1_3_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_6946, subc_out[11]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_6540, add_sub1_3_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_6539, add_sub1_3_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_6602, subc_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_6947, add_sub1_3_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_6303, add_sub1_3_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_7219, subc_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_6673, add_sub1_3_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6302, add_sub1_3_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_6947, add_sub1_3_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_6603, add_sub1_3_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_5761, addc_in[9]}), .c ({new_AGEMA_signal_6673, add_sub1_3_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_6540, add_sub1_3_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_6452, add_sub1_3_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_6603, add_sub1_3_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_6453, add_sub1_3_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_5767, addc_in[11]}), .c ({new_AGEMA_signal_6540, add_sub1_3_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5758, addc_in[8]}), .b ({new_AGEMA_signal_6301, add_sub1_3_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r (Fresh[218]), .c ({new_AGEMA_signal_6452, add_sub1_3_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6300, add_sub1_3_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_6304, add_sub1_3_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r (Fresh[219]), .c ({new_AGEMA_signal_6453, add_sub1_3_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_6674, add_sub1_3_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6456, add_sub1_3_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_6948, subc_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_6543, add_sub1_3_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_6542, add_sub1_3_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_6604, subc_out[6]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_6949, add_sub1_3_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_6310, add_sub1_3_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_7220, subc_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_6674, add_sub1_3_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6309, add_sub1_3_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_6949, add_sub1_3_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_6605, add_sub1_3_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_5749, addc_in[5]}), .c ({new_AGEMA_signal_6674, add_sub1_3_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_6543, add_sub1_3_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_6457, add_sub1_3_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_6605, add_sub1_3_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_6458, add_sub1_3_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_5755, addc_in[7]}), .c ({new_AGEMA_signal_6543, add_sub1_3_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5746, addc_in[4]}), .b ({new_AGEMA_signal_6308, add_sub1_3_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r (Fresh[220]), .c ({new_AGEMA_signal_6457, add_sub1_3_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6307, add_sub1_3_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_6311, add_sub1_3_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r (Fresh[221]), .c ({new_AGEMA_signal_6458, add_sub1_3_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_6675, add_sub1_3_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6461, add_sub1_3_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_6950, subc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_6546, add_sub1_3_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_6545, add_sub1_3_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_6606, subc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_6951, add_sub1_3_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_6317, add_sub1_3_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_7221, subc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_6675, add_sub1_3_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6316, add_sub1_3_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_6951, add_sub1_3_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_6607, add_sub1_3_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_5737, addc_in[1]}), .c ({new_AGEMA_signal_6675, add_sub1_3_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_6546, add_sub1_3_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_6462, add_sub1_3_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_6607, add_sub1_3_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_6463, add_sub1_3_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_5743, addc_in[3]}), .c ({new_AGEMA_signal_6546, add_sub1_3_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5734, addc_in[0]}), .b ({new_AGEMA_signal_6315, add_sub1_3_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r (Fresh[222]), .c ({new_AGEMA_signal_6462, add_sub1_3_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6314, add_sub1_3_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_6318, add_sub1_3_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r (Fresh[223]), .c ({new_AGEMA_signal_6463, add_sub1_3_subc_rom_sbox_0_ANF_2_t6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7185, subc_out[97]}), .a ({new_AGEMA_signal_7181, subc_out[113]}), .c ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6561, subc_out[98]}), .a ({new_AGEMA_signal_6553, subc_out[114]}), .c ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6887, subc_out[99]}), .a ({new_AGEMA_signal_6879, subc_out[115]}), .c ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7184, subc_out[101]}), .a ({new_AGEMA_signal_7180, subc_out[117]}), .c ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6559, subc_out[102]}), .a ({new_AGEMA_signal_6551, subc_out[118]}), .c ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6885, subc_out[103]}), .a ({new_AGEMA_signal_6877, subc_out[119]}), .c ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7183, subc_out[105]}), .a ({new_AGEMA_signal_7179, subc_out[121]}), .c ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6557, subc_out[106]}), .a ({new_AGEMA_signal_6549, subc_out[122]}), .c ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6883, subc_out[107]}), .a ({new_AGEMA_signal_6875, subc_out[123]}), .c ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7182, subc_out[109]}), .a ({new_AGEMA_signal_9048, subc_out[125]}), .c ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6555, subc_out[110]}), .a ({new_AGEMA_signal_7606, subc_out[126]}), .c ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6881, subc_out[111]}), .a ({new_AGEMA_signal_8572, subc_out[127]}), .c ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7181, subc_out[113]}), .a ({new_AGEMA_signal_7185, subc_out[97]}), .c ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6553, subc_out[114]}), .a ({new_AGEMA_signal_6561, subc_out[98]}), .c ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6879, subc_out[115]}), .a ({new_AGEMA_signal_6887, subc_out[99]}), .c ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7180, subc_out[117]}), .a ({new_AGEMA_signal_7184, subc_out[101]}), .c ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6551, subc_out[118]}), .a ({new_AGEMA_signal_6559, subc_out[102]}), .c ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6877, subc_out[119]}), .a ({new_AGEMA_signal_6885, subc_out[103]}), .c ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7179, subc_out[121]}), .a ({new_AGEMA_signal_7183, subc_out[105]}), .c ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6549, subc_out[122]}), .a ({new_AGEMA_signal_6557, subc_out[106]}), .c ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6875, subc_out[123]}), .a ({new_AGEMA_signal_6883, subc_out[107]}), .c ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9048, subc_out[125]}), .a ({new_AGEMA_signal_7182, subc_out[109]}), .c ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7606, subc_out[126]}), .a ({new_AGEMA_signal_6555, subc_out[110]}), .c ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8572, subc_out[127]}), .a ({new_AGEMA_signal_6881, subc_out[111]}), .c ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9049, subc_out[93]}), .a ({new_AGEMA_signal_7194, subc_out[77]}), .c ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7608, subc_out[94]}), .a ({new_AGEMA_signal_6570, subc_out[78]}), .c ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8574, subc_out[95]}), .a ({new_AGEMA_signal_6902, subc_out[79]}), .c ({new_AGEMA_signal_9054, shiftr_out[67]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7197, subc_out[65]}), .a ({new_AGEMA_signal_7193, subc_out[81]}), .c ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6576, subc_out[66]}), .a ({new_AGEMA_signal_6568, subc_out[82]}), .c ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6908, subc_out[67]}), .a ({new_AGEMA_signal_6900, subc_out[83]}), .c ({new_AGEMA_signal_7228, shiftr_out[71]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7196, subc_out[69]}), .a ({new_AGEMA_signal_7192, subc_out[85]}), .c ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6574, subc_out[70]}), .a ({new_AGEMA_signal_6566, subc_out[86]}), .c ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6906, subc_out[71]}), .a ({new_AGEMA_signal_6898, subc_out[87]}), .c ({new_AGEMA_signal_7229, shiftr_out[75]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7195, subc_out[73]}), .a ({new_AGEMA_signal_7191, subc_out[89]}), .c ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6572, subc_out[74]}), .a ({new_AGEMA_signal_6564, subc_out[90]}), .c ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6904, subc_out[75]}), .a ({new_AGEMA_signal_6896, subc_out[91]}), .c ({new_AGEMA_signal_7230, shiftr_out[79]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7194, subc_out[77]}), .a ({new_AGEMA_signal_9049, subc_out[93]}), .c ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6570, subc_out[78]}), .a ({new_AGEMA_signal_7608, subc_out[94]}), .c ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6902, subc_out[79]}), .a ({new_AGEMA_signal_8574, subc_out[95]}), .c ({new_AGEMA_signal_9055, shiftr_out[83]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7193, subc_out[81]}), .a ({new_AGEMA_signal_7197, subc_out[65]}), .c ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6568, subc_out[82]}), .a ({new_AGEMA_signal_6576, subc_out[66]}), .c ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6900, subc_out[83]}), .a ({new_AGEMA_signal_6908, subc_out[67]}), .c ({new_AGEMA_signal_7231, shiftr_out[87]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7192, subc_out[85]}), .a ({new_AGEMA_signal_7196, subc_out[69]}), .c ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6566, subc_out[86]}), .a ({new_AGEMA_signal_6574, subc_out[70]}), .c ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6898, subc_out[87]}), .a ({new_AGEMA_signal_6906, subc_out[71]}), .c ({new_AGEMA_signal_7232, shiftr_out[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7191, subc_out[89]}), .a ({new_AGEMA_signal_7195, subc_out[73]}), .c ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6564, subc_out[90]}), .a ({new_AGEMA_signal_6572, subc_out[74]}), .c ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6896, subc_out[91]}), .a ({new_AGEMA_signal_6904, subc_out[75]}), .c ({new_AGEMA_signal_7233, shiftr_out[95]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7203, subc_out[57]}), .a ({new_AGEMA_signal_7207, subc_out[41]}), .c ({new_AGEMA_signal_7300, shiftr_out[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6579, subc_out[58]}), .a ({new_AGEMA_signal_6587, subc_out[42]}), .c ({new_AGEMA_signal_6688, shiftr_out[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6917, subc_out[59]}), .a ({new_AGEMA_signal_6925, subc_out[43]}), .c ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9050, subc_out[61]}), .a ({new_AGEMA_signal_7206, subc_out[45]}), .c ({new_AGEMA_signal_9360, shiftr_out[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7610, subc_out[62]}), .a ({new_AGEMA_signal_6585, subc_out[46]}), .c ({new_AGEMA_signal_8098, shiftr_out[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8576, subc_out[63]}), .a ({new_AGEMA_signal_6923, subc_out[47]}), .c ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7209, subc_out[33]}), .a ({new_AGEMA_signal_7205, subc_out[49]}), .c ({new_AGEMA_signal_7301, shiftr_out[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6591, subc_out[34]}), .a ({new_AGEMA_signal_6583, subc_out[50]}), .c ({new_AGEMA_signal_6689, shiftr_out[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6929, subc_out[35]}), .a ({new_AGEMA_signal_6921, subc_out[51]}), .c ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7208, subc_out[37]}), .a ({new_AGEMA_signal_7204, subc_out[53]}), .c ({new_AGEMA_signal_7302, shiftr_out[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6589, subc_out[38]}), .a ({new_AGEMA_signal_6581, subc_out[54]}), .c ({new_AGEMA_signal_6690, shiftr_out[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6927, subc_out[39]}), .a ({new_AGEMA_signal_6919, subc_out[55]}), .c ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7207, subc_out[41]}), .a ({new_AGEMA_signal_7203, subc_out[57]}), .c ({new_AGEMA_signal_7303, shiftr_out[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6587, subc_out[42]}), .a ({new_AGEMA_signal_6579, subc_out[58]}), .c ({new_AGEMA_signal_6691, shiftr_out[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6925, subc_out[43]}), .a ({new_AGEMA_signal_6917, subc_out[59]}), .c ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7206, subc_out[45]}), .a ({new_AGEMA_signal_9050, subc_out[61]}), .c ({new_AGEMA_signal_9361, shiftr_out[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6585, subc_out[46]}), .a ({new_AGEMA_signal_7610, subc_out[62]}), .c ({new_AGEMA_signal_8099, shiftr_out[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6923, subc_out[47]}), .a ({new_AGEMA_signal_8576, subc_out[63]}), .c ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7205, subc_out[49]}), .a ({new_AGEMA_signal_7209, subc_out[33]}), .c ({new_AGEMA_signal_7304, shiftr_out[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6583, subc_out[50]}), .a ({new_AGEMA_signal_6591, subc_out[34]}), .c ({new_AGEMA_signal_6692, shiftr_out[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6921, subc_out[51]}), .a ({new_AGEMA_signal_6929, subc_out[35]}), .c ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7204, subc_out[53]}), .a ({new_AGEMA_signal_7208, subc_out[37]}), .c ({new_AGEMA_signal_7305, shiftr_out[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6581, subc_out[54]}), .a ({new_AGEMA_signal_6589, subc_out[38]}), .c ({new_AGEMA_signal_6693, shiftr_out[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6919, subc_out[55]}), .a ({new_AGEMA_signal_6927, subc_out[39]}), .c ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7216, subc_out[21]}), .a ({new_AGEMA_signal_7220, subc_out[5]}), .c ({new_AGEMA_signal_7306, shiftr_out[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6596, subc_out[22]}), .a ({new_AGEMA_signal_6604, subc_out[6]}), .c ({new_AGEMA_signal_6694, shiftr_out[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6940, subc_out[23]}), .a ({new_AGEMA_signal_6948, subc_out[7]}), .c ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7215, subc_out[25]}), .a ({new_AGEMA_signal_7219, subc_out[9]}), .c ({new_AGEMA_signal_7307, shiftr_out[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6594, subc_out[26]}), .a ({new_AGEMA_signal_6602, subc_out[10]}), .c ({new_AGEMA_signal_6695, shiftr_out[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6938, subc_out[27]}), .a ({new_AGEMA_signal_6946, subc_out[11]}), .c ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9051, subc_out[29]}), .a ({new_AGEMA_signal_7218, subc_out[13]}), .c ({new_AGEMA_signal_9362, shiftr_out[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7612, subc_out[30]}), .a ({new_AGEMA_signal_6600, subc_out[14]}), .c ({new_AGEMA_signal_8100, shiftr_out[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8578, subc_out[31]}), .a ({new_AGEMA_signal_6944, subc_out[15]}), .c ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7221, subc_out[1]}), .a ({new_AGEMA_signal_7217, subc_out[17]}), .c ({new_AGEMA_signal_7308, shiftr_out[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6606, subc_out[2]}), .a ({new_AGEMA_signal_6598, subc_out[18]}), .c ({new_AGEMA_signal_6696, shiftr_out[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6950, subc_out[3]}), .a ({new_AGEMA_signal_6942, subc_out[19]}), .c ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7220, subc_out[5]}), .a ({new_AGEMA_signal_7216, subc_out[21]}), .c ({new_AGEMA_signal_7309, shiftr_out[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6604, subc_out[6]}), .a ({new_AGEMA_signal_6596, subc_out[22]}), .c ({new_AGEMA_signal_6697, shiftr_out[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6948, subc_out[7]}), .a ({new_AGEMA_signal_6940, subc_out[23]}), .c ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7219, subc_out[9]}), .a ({new_AGEMA_signal_7215, subc_out[25]}), .c ({new_AGEMA_signal_7310, shiftr_out[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6602, subc_out[10]}), .a ({new_AGEMA_signal_6594, subc_out[26]}), .c ({new_AGEMA_signal_6698, shiftr_out[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6946, subc_out[11]}), .a ({new_AGEMA_signal_6938, subc_out[27]}), .c ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7218, subc_out[13]}), .a ({new_AGEMA_signal_9051, subc_out[29]}), .c ({new_AGEMA_signal_9363, shiftr_out[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6600, subc_out[14]}), .a ({new_AGEMA_signal_7612, subc_out[30]}), .c ({new_AGEMA_signal_8101, shiftr_out[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6944, subc_out[15]}), .a ({new_AGEMA_signal_8578, subc_out[31]}), .c ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7217, subc_out[17]}), .a ({new_AGEMA_signal_7221, subc_out[1]}), .c ({new_AGEMA_signal_7311, shiftr_out[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6598, subc_out[18]}), .a ({new_AGEMA_signal_6606, subc_out[2]}), .c ({new_AGEMA_signal_6699, shiftr_out[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_6942, subc_out[19]}), .a ({new_AGEMA_signal_6950, subc_out[3]}), .c ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U44 ( .a ({new_AGEMA_signal_7325, mcs1_mcs_mat1_0_mcs_out[90]}), .b ({new_AGEMA_signal_9629, mcs1_mcs_mat1_0_mcs_out[94]}), .c ({new_AGEMA_signal_9863, mcs1_mcs_mat1_0_n93}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({new_AGEMA_signal_7615, shiftr_out[124]}), .c ({new_AGEMA_signal_9380, mcs1_mcs_mat1_0_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_6619, shiftr_out[92]}), .b ({new_AGEMA_signal_6700, mcs1_mcs_mat1_0_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_6952, mcs1_mcs_mat1_0_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6619, shiftr_out[92]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[224]), .c ({new_AGEMA_signal_6700, mcs1_mcs_mat1_0_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_7314, mcs1_mcs_mat1_0_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_7624, mcs1_mcs_mat1_0_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_6701, mcs1_mcs_mat1_0_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_7314, mcs1_mcs_mat1_0_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[225]), .c ({new_AGEMA_signal_6701, mcs1_mcs_mat1_0_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_6702, mcs1_mcs_mat1_0_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_7628, mcs1_mcs_mat1_0_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8106, mcs1_mcs_mat1_0_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_6955, mcs1_mcs_mat1_0_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_7317, mcs1_mcs_mat1_0_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_6699, shiftr_out[30]}), .c ({new_AGEMA_signal_6955, mcs1_mcs_mat1_0_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_7311, shiftr_out[29]}), .b ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_7628, mcs1_mcs_mat1_0_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[226]), .c ({new_AGEMA_signal_6702, mcs1_mcs_mat1_0_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_9626, mcs1_mcs_mat1_0_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_9868, mcs1_mcs_mat1_0_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_8109, mcs1_mcs_mat1_0_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_9626, mcs1_mcs_mat1_0_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[227]), .c ({new_AGEMA_signal_8109, mcs1_mcs_mat1_0_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6619, shiftr_out[92]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[228]), .c ({new_AGEMA_signal_6703, mcs1_mcs_mat1_0_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({new_AGEMA_signal_7321, mcs1_mcs_mat1_0_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_7632, mcs1_mcs_mat1_0_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_6704, mcs1_mcs_mat1_0_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_7321, mcs1_mcs_mat1_0_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_7305, shiftr_out[61]}), .b ({new_AGEMA_signal_6693, shiftr_out[62]}), .c ({new_AGEMA_signal_7633, mcs1_mcs_mat1_0_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[229]), .c ({new_AGEMA_signal_6704, mcs1_mcs_mat1_0_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_6705, mcs1_mcs_mat1_0_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_7323, mcs1_mcs_mat1_0_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_6705, mcs1_mcs_mat1_0_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .c ({new_AGEMA_signal_6959, mcs1_mcs_mat1_0_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[230]), .c ({new_AGEMA_signal_6705, mcs1_mcs_mat1_0_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_9383, mcs1_mcs_mat1_0_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_7615, shiftr_out[124]}), .c ({new_AGEMA_signal_9629, mcs1_mcs_mat1_0_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_8116, mcs1_mcs_mat1_0_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_9383, mcs1_mcs_mat1_0_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_9384, mcs1_mcs_mat1_0_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[231]), .c ({new_AGEMA_signal_8116, mcs1_mcs_mat1_0_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_7233, shiftr_out[95]}), .b ({new_AGEMA_signal_6619, shiftr_out[92]}), .c ({new_AGEMA_signal_7325, mcs1_mcs_mat1_0_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_7233, shiftr_out[95]}), .b ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_7326, mcs1_mcs_mat1_0_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({new_AGEMA_signal_7637, mcs1_mcs_mat1_0_mcs_out[87]}), .c ({new_AGEMA_signal_8117, mcs1_mcs_mat1_0_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_7305, shiftr_out[61]}), .c ({new_AGEMA_signal_7637, mcs1_mcs_mat1_0_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_7311, shiftr_out[29]}), .c ({new_AGEMA_signal_7640, mcs1_mcs_mat1_0_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[232]), .c ({new_AGEMA_signal_6706, mcs1_mcs_mat1_0_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_8122, mcs1_mcs_mat1_0_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_8606, mcs1_mcs_mat1_0_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[233]), .c ({new_AGEMA_signal_8122, mcs1_mcs_mat1_0_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_6707, mcs1_mcs_mat1_0_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_6962, mcs1_mcs_mat1_0_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6619, shiftr_out[92]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[234]), .c ({new_AGEMA_signal_6707, mcs1_mcs_mat1_0_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[235]), .c ({new_AGEMA_signal_6708, mcs1_mcs_mat1_0_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_6709, mcs1_mcs_mat1_0_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7311, shiftr_out[29]}), .c ({new_AGEMA_signal_7648, mcs1_mcs_mat1_0_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[236]), .c ({new_AGEMA_signal_6709, mcs1_mcs_mat1_0_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_10084, mcs1_mcs_mat1_0_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_8128, mcs1_mcs_mat1_0_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_10328, mcs1_mcs_mat1_0_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_9874, mcs1_mcs_mat1_0_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_10084, mcs1_mcs_mat1_0_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_9634, mcs1_mcs_mat1_0_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_9874, mcs1_mcs_mat1_0_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_9634, mcs1_mcs_mat1_0_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[237]), .c ({new_AGEMA_signal_8128, mcs1_mcs_mat1_0_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_7651, mcs1_mcs_mat1_0_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_6966, mcs1_mcs_mat1_0_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_8129, mcs1_mcs_mat1_0_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_6710, mcs1_mcs_mat1_0_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_6619, shiftr_out[92]}), .c ({new_AGEMA_signal_6966, mcs1_mcs_mat1_0_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_6619, shiftr_out[92]}), .c ({new_AGEMA_signal_6967, mcs1_mcs_mat1_0_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_7233, shiftr_out[95]}), .c ({new_AGEMA_signal_7651, mcs1_mcs_mat1_0_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_6710, mcs1_mcs_mat1_0_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_7652, mcs1_mcs_mat1_0_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6619, shiftr_out[92]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[238]), .c ({new_AGEMA_signal_6710, mcs1_mcs_mat1_0_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_7305, shiftr_out[61]}), .b ({new_AGEMA_signal_6711, mcs1_mcs_mat1_0_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_7656, mcs1_mcs_mat1_0_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[239]), .c ({new_AGEMA_signal_6711, mcs1_mcs_mat1_0_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({new_AGEMA_signal_7658, mcs1_mcs_mat1_0_mcs_out[51]}), .c ({new_AGEMA_signal_8134, mcs1_mcs_mat1_0_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_7311, shiftr_out[29]}), .c ({new_AGEMA_signal_7658, mcs1_mcs_mat1_0_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_8135, mcs1_mcs_mat1_0_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_9389, mcs1_mcs_mat1_0_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[240]), .c ({new_AGEMA_signal_8135, mcs1_mcs_mat1_0_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_7659, mcs1_mcs_mat1_0_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_8137, mcs1_mcs_mat1_0_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_6619, shiftr_out[92]}), .b ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_7659, mcs1_mcs_mat1_0_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_7334, mcs1_mcs_mat1_0_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_7660, mcs1_mcs_mat1_0_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_7233, shiftr_out[95]}), .c ({new_AGEMA_signal_7334, mcs1_mcs_mat1_0_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6619, shiftr_out[92]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[241]), .c ({new_AGEMA_signal_6712, mcs1_mcs_mat1_0_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({new_AGEMA_signal_6713, mcs1_mcs_mat1_0_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_7336, mcs1_mcs_mat1_0_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_7305, shiftr_out[61]}), .b ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_7663, mcs1_mcs_mat1_0_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[242]), .c ({new_AGEMA_signal_6713, mcs1_mcs_mat1_0_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_8625, mcs1_mcs_mat1_0_mcs_out[35]}), .b ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_9085, mcs1_mcs_mat1_0_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_8143, mcs1_mcs_mat1_0_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_6714, mcs1_mcs_mat1_0_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_8625, mcs1_mcs_mat1_0_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_7665, mcs1_mcs_mat1_0_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_6699, shiftr_out[30]}), .c ({new_AGEMA_signal_8143, mcs1_mcs_mat1_0_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_7311, shiftr_out[29]}), .c ({new_AGEMA_signal_7665, mcs1_mcs_mat1_0_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[243]), .c ({new_AGEMA_signal_6714, mcs1_mcs_mat1_0_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_8144, mcs1_mcs_mat1_0_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_8626, mcs1_mcs_mat1_0_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({new_AGEMA_signal_9638, mcs1_mcs_mat1_0_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_9877, mcs1_mcs_mat1_0_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_8144, mcs1_mcs_mat1_0_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_9638, mcs1_mcs_mat1_0_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[244]), .c ({new_AGEMA_signal_8144, mcs1_mcs_mat1_0_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6619, shiftr_out[92]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[245]), .c ({new_AGEMA_signal_6715, mcs1_mcs_mat1_0_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[246]), .c ({new_AGEMA_signal_6716, mcs1_mcs_mat1_0_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_7342, mcs1_mcs_mat1_0_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_7673, mcs1_mcs_mat1_0_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_7342, mcs1_mcs_mat1_0_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_7311, shiftr_out[29]}), .c ({new_AGEMA_signal_7675, mcs1_mcs_mat1_0_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[247]), .c ({new_AGEMA_signal_6717, mcs1_mcs_mat1_0_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[248]), .c ({new_AGEMA_signal_8154, mcs1_mcs_mat1_0_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6619, shiftr_out[92]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[249]), .c ({new_AGEMA_signal_6718, mcs1_mcs_mat1_0_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_6719, mcs1_mcs_mat1_0_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_7346, mcs1_mcs_mat1_0_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_6719, mcs1_mcs_mat1_0_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_6977, mcs1_mcs_mat1_0_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[250]), .c ({new_AGEMA_signal_6719, mcs1_mcs_mat1_0_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_7681, mcs1_mcs_mat1_0_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_6720, mcs1_mcs_mat1_0_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8158, mcs1_mcs_mat1_0_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_7681, mcs1_mcs_mat1_0_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7311, shiftr_out[29]}), .c ({new_AGEMA_signal_8160, mcs1_mcs_mat1_0_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_7348, mcs1_mcs_mat1_0_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_7681, mcs1_mcs_mat1_0_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_7348, mcs1_mcs_mat1_0_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_7311, shiftr_out[29]}), .c ({new_AGEMA_signal_7682, mcs1_mcs_mat1_0_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[251]), .c ({new_AGEMA_signal_6720, mcs1_mcs_mat1_0_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U44 ( .a ({new_AGEMA_signal_7364, mcs1_mcs_mat1_1_mcs_out[90]}), .b ({new_AGEMA_signal_7697, mcs1_mcs_mat1_1_mcs_out[94]}), .c ({new_AGEMA_signal_8163, mcs1_mcs_mat1_1_n93}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({new_AGEMA_signal_6613, shiftr_out[120]}), .c ({new_AGEMA_signal_7350, mcs1_mcs_mat1_1_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_6618, shiftr_out[88]}), .b ({new_AGEMA_signal_6721, mcs1_mcs_mat1_1_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_6980, mcs1_mcs_mat1_1_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6618, shiftr_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[252]), .c ({new_AGEMA_signal_6721, mcs1_mcs_mat1_1_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_7353, mcs1_mcs_mat1_1_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_7686, mcs1_mcs_mat1_1_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_6722, mcs1_mcs_mat1_1_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_7353, mcs1_mcs_mat1_1_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[253]), .c ({new_AGEMA_signal_6722, mcs1_mcs_mat1_1_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_8169, mcs1_mcs_mat1_1_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9650, mcs1_mcs_mat1_1_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_9887, mcs1_mcs_mat1_1_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_8650, mcs1_mcs_mat1_1_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_9409, mcs1_mcs_mat1_1_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_8101, shiftr_out[26]}), .c ({new_AGEMA_signal_8650, mcs1_mcs_mat1_1_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_9363, shiftr_out[25]}), .b ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_9650, mcs1_mcs_mat1_1_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[254]), .c ({new_AGEMA_signal_8169, mcs1_mcs_mat1_1_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_7689, mcs1_mcs_mat1_1_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_8170, mcs1_mcs_mat1_1_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_6723, mcs1_mcs_mat1_1_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_7689, mcs1_mcs_mat1_1_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[255]), .c ({new_AGEMA_signal_6723, mcs1_mcs_mat1_1_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6618, shiftr_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[256]), .c ({new_AGEMA_signal_6724, mcs1_mcs_mat1_1_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({new_AGEMA_signal_7359, mcs1_mcs_mat1_1_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_7693, mcs1_mcs_mat1_1_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_6725, mcs1_mcs_mat1_1_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_7359, mcs1_mcs_mat1_1_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_7304, shiftr_out[57]}), .b ({new_AGEMA_signal_6692, shiftr_out[58]}), .c ({new_AGEMA_signal_7694, mcs1_mcs_mat1_1_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[257]), .c ({new_AGEMA_signal_6725, mcs1_mcs_mat1_1_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_8177, mcs1_mcs_mat1_1_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_9411, mcs1_mcs_mat1_1_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_8177, mcs1_mcs_mat1_1_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .c ({new_AGEMA_signal_8660, mcs1_mcs_mat1_1_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[258]), .c ({new_AGEMA_signal_8177, mcs1_mcs_mat1_1_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_7361, mcs1_mcs_mat1_1_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_6613, shiftr_out[120]}), .c ({new_AGEMA_signal_7697, mcs1_mcs_mat1_1_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_6726, mcs1_mcs_mat1_1_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_7361, mcs1_mcs_mat1_1_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_7362, mcs1_mcs_mat1_1_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[259]), .c ({new_AGEMA_signal_6726, mcs1_mcs_mat1_1_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_7232, shiftr_out[91]}), .b ({new_AGEMA_signal_6618, shiftr_out[88]}), .c ({new_AGEMA_signal_7364, mcs1_mcs_mat1_1_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_7232, shiftr_out[91]}), .b ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_7365, mcs1_mcs_mat1_1_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({new_AGEMA_signal_7700, mcs1_mcs_mat1_1_mcs_out[87]}), .c ({new_AGEMA_signal_8179, mcs1_mcs_mat1_1_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_7304, shiftr_out[57]}), .c ({new_AGEMA_signal_7700, mcs1_mcs_mat1_1_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_9363, shiftr_out[25]}), .c ({new_AGEMA_signal_9655, mcs1_mcs_mat1_1_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[260]), .c ({new_AGEMA_signal_8180, mcs1_mcs_mat1_1_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_6727, mcs1_mcs_mat1_1_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_6987, mcs1_mcs_mat1_1_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[261]), .c ({new_AGEMA_signal_6727, mcs1_mcs_mat1_1_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_6728, mcs1_mcs_mat1_1_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_6989, mcs1_mcs_mat1_1_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6618, shiftr_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[262]), .c ({new_AGEMA_signal_6728, mcs1_mcs_mat1_1_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[263]), .c ({new_AGEMA_signal_6729, mcs1_mcs_mat1_1_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_8186, mcs1_mcs_mat1_1_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_9363, shiftr_out[25]}), .c ({new_AGEMA_signal_9657, mcs1_mcs_mat1_1_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[264]), .c ({new_AGEMA_signal_8186, mcs1_mcs_mat1_1_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_8674, mcs1_mcs_mat1_1_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_6730, mcs1_mcs_mat1_1_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_9119, mcs1_mcs_mat1_1_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_8189, mcs1_mcs_mat1_1_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_8674, mcs1_mcs_mat1_1_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_7709, mcs1_mcs_mat1_1_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8189, mcs1_mcs_mat1_1_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_7709, mcs1_mcs_mat1_1_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[265]), .c ({new_AGEMA_signal_6730, mcs1_mcs_mat1_1_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_7712, mcs1_mcs_mat1_1_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_6993, mcs1_mcs_mat1_1_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_8190, mcs1_mcs_mat1_1_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_6731, mcs1_mcs_mat1_1_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_6618, shiftr_out[88]}), .c ({new_AGEMA_signal_6993, mcs1_mcs_mat1_1_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_6618, shiftr_out[88]}), .c ({new_AGEMA_signal_6994, mcs1_mcs_mat1_1_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_7232, shiftr_out[91]}), .c ({new_AGEMA_signal_7712, mcs1_mcs_mat1_1_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_6731, mcs1_mcs_mat1_1_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_7713, mcs1_mcs_mat1_1_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6618, shiftr_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[266]), .c ({new_AGEMA_signal_6731, mcs1_mcs_mat1_1_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_7304, shiftr_out[57]}), .b ({new_AGEMA_signal_6732, mcs1_mcs_mat1_1_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_7717, mcs1_mcs_mat1_1_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[267]), .c ({new_AGEMA_signal_6732, mcs1_mcs_mat1_1_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({new_AGEMA_signal_9659, mcs1_mcs_mat1_1_mcs_out[51]}), .c ({new_AGEMA_signal_9896, mcs1_mcs_mat1_1_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_9363, shiftr_out[25]}), .c ({new_AGEMA_signal_9659, mcs1_mcs_mat1_1_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_6733, mcs1_mcs_mat1_1_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_7373, mcs1_mcs_mat1_1_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[268]), .c ({new_AGEMA_signal_6733, mcs1_mcs_mat1_1_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_7721, mcs1_mcs_mat1_1_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_8197, mcs1_mcs_mat1_1_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_6618, shiftr_out[88]}), .b ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_7721, mcs1_mcs_mat1_1_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_7375, mcs1_mcs_mat1_1_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_7722, mcs1_mcs_mat1_1_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_7232, shiftr_out[91]}), .c ({new_AGEMA_signal_7375, mcs1_mcs_mat1_1_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6618, shiftr_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[269]), .c ({new_AGEMA_signal_6734, mcs1_mcs_mat1_1_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({new_AGEMA_signal_6735, mcs1_mcs_mat1_1_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_7377, mcs1_mcs_mat1_1_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_7304, shiftr_out[57]}), .b ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_7725, mcs1_mcs_mat1_1_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[270]), .c ({new_AGEMA_signal_6735, mcs1_mcs_mat1_1_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_10112, mcs1_mcs_mat1_1_mcs_out[35]}), .b ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_10356, mcs1_mcs_mat1_1_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_9898, mcs1_mcs_mat1_1_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_8202, mcs1_mcs_mat1_1_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_10112, mcs1_mcs_mat1_1_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_9660, mcs1_mcs_mat1_1_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_8101, shiftr_out[26]}), .c ({new_AGEMA_signal_9898, mcs1_mcs_mat1_1_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_9363, shiftr_out[25]}), .c ({new_AGEMA_signal_9660, mcs1_mcs_mat1_1_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[271]), .c ({new_AGEMA_signal_8202, mcs1_mcs_mat1_1_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_6736, mcs1_mcs_mat1_1_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_7000, mcs1_mcs_mat1_1_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({new_AGEMA_signal_7727, mcs1_mcs_mat1_1_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_8204, mcs1_mcs_mat1_1_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_6736, mcs1_mcs_mat1_1_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_7727, mcs1_mcs_mat1_1_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[272]), .c ({new_AGEMA_signal_6736, mcs1_mcs_mat1_1_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6618, shiftr_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[273]), .c ({new_AGEMA_signal_6737, mcs1_mcs_mat1_1_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[274]), .c ({new_AGEMA_signal_6738, mcs1_mcs_mat1_1_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_9417, mcs1_mcs_mat1_1_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_9662, mcs1_mcs_mat1_1_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_9417, mcs1_mcs_mat1_1_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_9363, shiftr_out[25]}), .c ({new_AGEMA_signal_9664, mcs1_mcs_mat1_1_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[275]), .c ({new_AGEMA_signal_8212, mcs1_mcs_mat1_1_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[276]), .c ({new_AGEMA_signal_6739, mcs1_mcs_mat1_1_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6618, shiftr_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[277]), .c ({new_AGEMA_signal_6740, mcs1_mcs_mat1_1_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_6741, mcs1_mcs_mat1_1_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_7386, mcs1_mcs_mat1_1_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_6741, mcs1_mcs_mat1_1_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_7006, mcs1_mcs_mat1_1_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[278]), .c ({new_AGEMA_signal_6741, mcs1_mcs_mat1_1_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_9668, mcs1_mcs_mat1_1_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8219, mcs1_mcs_mat1_1_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_9902, mcs1_mcs_mat1_1_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_9668, mcs1_mcs_mat1_1_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_9363, shiftr_out[25]}), .c ({new_AGEMA_signal_9904, mcs1_mcs_mat1_1_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_9421, mcs1_mcs_mat1_1_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_9668, mcs1_mcs_mat1_1_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_9421, mcs1_mcs_mat1_1_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_9363, shiftr_out[25]}), .c ({new_AGEMA_signal_9669, mcs1_mcs_mat1_1_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[279]), .c ({new_AGEMA_signal_8219, mcs1_mcs_mat1_1_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U44 ( .a ({new_AGEMA_signal_7401, mcs1_mcs_mat1_2_mcs_out[90]}), .b ({new_AGEMA_signal_7751, mcs1_mcs_mat1_2_mcs_out[94]}), .c ({new_AGEMA_signal_8221, mcs1_mcs_mat1_2_n93}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({new_AGEMA_signal_6612, shiftr_out[116]}), .c ({new_AGEMA_signal_7388, mcs1_mcs_mat1_2_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_6617, shiftr_out[84]}), .b ({new_AGEMA_signal_6742, mcs1_mcs_mat1_2_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_7008, mcs1_mcs_mat1_2_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6617, shiftr_out[84]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[280]), .c ({new_AGEMA_signal_6742, mcs1_mcs_mat1_2_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_9437, mcs1_mcs_mat1_2_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_9675, mcs1_mcs_mat1_2_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_8225, mcs1_mcs_mat1_2_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_9437, mcs1_mcs_mat1_2_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[281]), .c ({new_AGEMA_signal_8225, mcs1_mcs_mat1_2_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_6743, mcs1_mcs_mat1_2_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_7744, mcs1_mcs_mat1_2_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8226, mcs1_mcs_mat1_2_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_7010, mcs1_mcs_mat1_2_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_7391, mcs1_mcs_mat1_2_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_6698, shiftr_out[22]}), .c ({new_AGEMA_signal_7010, mcs1_mcs_mat1_2_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_7310, shiftr_out[21]}), .b ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_7744, mcs1_mcs_mat1_2_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[282]), .c ({new_AGEMA_signal_6743, mcs1_mcs_mat1_2_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_7746, mcs1_mcs_mat1_2_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_8229, mcs1_mcs_mat1_2_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_6744, mcs1_mcs_mat1_2_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_7746, mcs1_mcs_mat1_2_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[283]), .c ({new_AGEMA_signal_6744, mcs1_mcs_mat1_2_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6617, shiftr_out[84]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[284]), .c ({new_AGEMA_signal_6745, mcs1_mcs_mat1_2_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({new_AGEMA_signal_9440, mcs1_mcs_mat1_2_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_9678, mcs1_mcs_mat1_2_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_8233, mcs1_mcs_mat1_2_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_9440, mcs1_mcs_mat1_2_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_9361, shiftr_out[53]}), .b ({new_AGEMA_signal_8099, shiftr_out[54]}), .c ({new_AGEMA_signal_9679, mcs1_mcs_mat1_2_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[285]), .c ({new_AGEMA_signal_8233, mcs1_mcs_mat1_2_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_6746, mcs1_mcs_mat1_2_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_7396, mcs1_mcs_mat1_2_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_6746, mcs1_mcs_mat1_2_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .c ({new_AGEMA_signal_7014, mcs1_mcs_mat1_2_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[286]), .c ({new_AGEMA_signal_6746, mcs1_mcs_mat1_2_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_7398, mcs1_mcs_mat1_2_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_6612, shiftr_out[116]}), .c ({new_AGEMA_signal_7751, mcs1_mcs_mat1_2_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_6747, mcs1_mcs_mat1_2_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_7398, mcs1_mcs_mat1_2_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_7399, mcs1_mcs_mat1_2_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[287]), .c ({new_AGEMA_signal_6747, mcs1_mcs_mat1_2_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_7231, shiftr_out[87]}), .b ({new_AGEMA_signal_6617, shiftr_out[84]}), .c ({new_AGEMA_signal_7401, mcs1_mcs_mat1_2_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_7231, shiftr_out[87]}), .b ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_7402, mcs1_mcs_mat1_2_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({new_AGEMA_signal_9683, mcs1_mcs_mat1_2_mcs_out[87]}), .c ({new_AGEMA_signal_9916, mcs1_mcs_mat1_2_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_9361, shiftr_out[53]}), .c ({new_AGEMA_signal_9683, mcs1_mcs_mat1_2_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_7310, shiftr_out[21]}), .c ({new_AGEMA_signal_7756, mcs1_mcs_mat1_2_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[288]), .c ({new_AGEMA_signal_6748, mcs1_mcs_mat1_2_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_6749, mcs1_mcs_mat1_2_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_7018, mcs1_mcs_mat1_2_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[289]), .c ({new_AGEMA_signal_6749, mcs1_mcs_mat1_2_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_6750, mcs1_mcs_mat1_2_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_7020, mcs1_mcs_mat1_2_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6617, shiftr_out[84]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[290]), .c ({new_AGEMA_signal_6750, mcs1_mcs_mat1_2_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[291]), .c ({new_AGEMA_signal_8243, mcs1_mcs_mat1_2_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_6751, mcs1_mcs_mat1_2_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7310, shiftr_out[21]}), .c ({new_AGEMA_signal_7763, mcs1_mcs_mat1_2_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[292]), .c ({new_AGEMA_signal_6751, mcs1_mcs_mat1_2_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_8729, mcs1_mcs_mat1_2_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_6752, mcs1_mcs_mat1_2_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_9160, mcs1_mcs_mat1_2_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_8247, mcs1_mcs_mat1_2_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_8729, mcs1_mcs_mat1_2_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_7765, mcs1_mcs_mat1_2_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8247, mcs1_mcs_mat1_2_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_7765, mcs1_mcs_mat1_2_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[293]), .c ({new_AGEMA_signal_6752, mcs1_mcs_mat1_2_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_7768, mcs1_mcs_mat1_2_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_7024, mcs1_mcs_mat1_2_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_8248, mcs1_mcs_mat1_2_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_6753, mcs1_mcs_mat1_2_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_6617, shiftr_out[84]}), .c ({new_AGEMA_signal_7024, mcs1_mcs_mat1_2_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_6617, shiftr_out[84]}), .c ({new_AGEMA_signal_7025, mcs1_mcs_mat1_2_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_7231, shiftr_out[87]}), .c ({new_AGEMA_signal_7768, mcs1_mcs_mat1_2_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_6753, mcs1_mcs_mat1_2_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_7769, mcs1_mcs_mat1_2_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6617, shiftr_out[84]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[294]), .c ({new_AGEMA_signal_6753, mcs1_mcs_mat1_2_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_9361, shiftr_out[53]}), .b ({new_AGEMA_signal_8251, mcs1_mcs_mat1_2_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_9689, mcs1_mcs_mat1_2_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[295]), .c ({new_AGEMA_signal_8251, mcs1_mcs_mat1_2_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({new_AGEMA_signal_7771, mcs1_mcs_mat1_2_mcs_out[51]}), .c ({new_AGEMA_signal_8252, mcs1_mcs_mat1_2_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_7310, shiftr_out[21]}), .c ({new_AGEMA_signal_7771, mcs1_mcs_mat1_2_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_6754, mcs1_mcs_mat1_2_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_7409, mcs1_mcs_mat1_2_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[296]), .c ({new_AGEMA_signal_6754, mcs1_mcs_mat1_2_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_7774, mcs1_mcs_mat1_2_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_8255, mcs1_mcs_mat1_2_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_6617, shiftr_out[84]}), .b ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_7774, mcs1_mcs_mat1_2_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_7411, mcs1_mcs_mat1_2_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_7775, mcs1_mcs_mat1_2_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_7231, shiftr_out[87]}), .c ({new_AGEMA_signal_7411, mcs1_mcs_mat1_2_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6617, shiftr_out[84]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[297]), .c ({new_AGEMA_signal_6755, mcs1_mcs_mat1_2_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({new_AGEMA_signal_8258, mcs1_mcs_mat1_2_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9448, mcs1_mcs_mat1_2_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_9361, shiftr_out[53]}), .b ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_9692, mcs1_mcs_mat1_2_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[298]), .c ({new_AGEMA_signal_8258, mcs1_mcs_mat1_2_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_8737, mcs1_mcs_mat1_2_mcs_out[35]}), .b ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_9163, mcs1_mcs_mat1_2_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_8260, mcs1_mcs_mat1_2_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_6756, mcs1_mcs_mat1_2_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_8737, mcs1_mcs_mat1_2_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_7777, mcs1_mcs_mat1_2_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_6698, shiftr_out[22]}), .c ({new_AGEMA_signal_8260, mcs1_mcs_mat1_2_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_7310, shiftr_out[21]}), .c ({new_AGEMA_signal_7777, mcs1_mcs_mat1_2_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[299]), .c ({new_AGEMA_signal_6756, mcs1_mcs_mat1_2_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_6757, mcs1_mcs_mat1_2_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_7030, mcs1_mcs_mat1_2_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({new_AGEMA_signal_7779, mcs1_mcs_mat1_2_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_8262, mcs1_mcs_mat1_2_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_6757, mcs1_mcs_mat1_2_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_7779, mcs1_mcs_mat1_2_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[300]), .c ({new_AGEMA_signal_6757, mcs1_mcs_mat1_2_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6617, shiftr_out[84]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[301]), .c ({new_AGEMA_signal_6758, mcs1_mcs_mat1_2_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[302]), .c ({new_AGEMA_signal_8267, mcs1_mcs_mat1_2_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_7416, mcs1_mcs_mat1_2_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_7785, mcs1_mcs_mat1_2_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_7416, mcs1_mcs_mat1_2_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_7310, shiftr_out[21]}), .c ({new_AGEMA_signal_7787, mcs1_mcs_mat1_2_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[303]), .c ({new_AGEMA_signal_6759, mcs1_mcs_mat1_2_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[304]), .c ({new_AGEMA_signal_6760, mcs1_mcs_mat1_2_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6617, shiftr_out[84]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[305]), .c ({new_AGEMA_signal_6761, mcs1_mcs_mat1_2_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_8276, mcs1_mcs_mat1_2_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_9454, mcs1_mcs_mat1_2_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_8276, mcs1_mcs_mat1_2_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_8751, mcs1_mcs_mat1_2_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[306]), .c ({new_AGEMA_signal_8276, mcs1_mcs_mat1_2_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_7794, mcs1_mcs_mat1_2_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_6762, mcs1_mcs_mat1_2_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8277, mcs1_mcs_mat1_2_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_7794, mcs1_mcs_mat1_2_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7310, shiftr_out[21]}), .c ({new_AGEMA_signal_8279, mcs1_mcs_mat1_2_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_7421, mcs1_mcs_mat1_2_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_7794, mcs1_mcs_mat1_2_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_7421, mcs1_mcs_mat1_2_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_7310, shiftr_out[21]}), .c ({new_AGEMA_signal_7795, mcs1_mcs_mat1_2_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[307]), .c ({new_AGEMA_signal_6762, mcs1_mcs_mat1_2_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U44 ( .a ({new_AGEMA_signal_9477, mcs1_mcs_mat1_3_mcs_out[90]}), .b ({new_AGEMA_signal_7810, mcs1_mcs_mat1_3_mcs_out[94]}), .c ({new_AGEMA_signal_9701, mcs1_mcs_mat1_3_n93}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({new_AGEMA_signal_6611, shiftr_out[112]}), .c ({new_AGEMA_signal_7423, mcs1_mcs_mat1_3_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_7617, shiftr_out[80]}), .b ({new_AGEMA_signal_8281, mcs1_mcs_mat1_3_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8762, mcs1_mcs_mat1_3_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7617, shiftr_out[80]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[308]), .c ({new_AGEMA_signal_8281, mcs1_mcs_mat1_3_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_7424, mcs1_mcs_mat1_3_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_7797, mcs1_mcs_mat1_3_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_6763, mcs1_mcs_mat1_3_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_7424, mcs1_mcs_mat1_3_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[309]), .c ({new_AGEMA_signal_6763, mcs1_mcs_mat1_3_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_6764, mcs1_mcs_mat1_3_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_7801, mcs1_mcs_mat1_3_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8284, mcs1_mcs_mat1_3_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_7038, mcs1_mcs_mat1_3_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_7427, mcs1_mcs_mat1_3_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_6697, shiftr_out[18]}), .c ({new_AGEMA_signal_7038, mcs1_mcs_mat1_3_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_7309, shiftr_out[17]}), .b ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_7801, mcs1_mcs_mat1_3_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[310]), .c ({new_AGEMA_signal_6764, mcs1_mcs_mat1_3_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_7803, mcs1_mcs_mat1_3_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_8287, mcs1_mcs_mat1_3_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_6765, mcs1_mcs_mat1_3_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_7803, mcs1_mcs_mat1_3_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[311]), .c ({new_AGEMA_signal_6765, mcs1_mcs_mat1_3_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7617, shiftr_out[80]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[312]), .c ({new_AGEMA_signal_8289, mcs1_mcs_mat1_3_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({new_AGEMA_signal_7430, mcs1_mcs_mat1_3_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_7805, mcs1_mcs_mat1_3_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_6766, mcs1_mcs_mat1_3_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_7430, mcs1_mcs_mat1_3_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_7303, shiftr_out[49]}), .b ({new_AGEMA_signal_6691, shiftr_out[50]}), .c ({new_AGEMA_signal_7806, mcs1_mcs_mat1_3_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[313]), .c ({new_AGEMA_signal_6766, mcs1_mcs_mat1_3_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_6767, mcs1_mcs_mat1_3_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_7432, mcs1_mcs_mat1_3_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_6767, mcs1_mcs_mat1_3_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .c ({new_AGEMA_signal_7042, mcs1_mcs_mat1_3_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[314]), .c ({new_AGEMA_signal_6767, mcs1_mcs_mat1_3_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_7434, mcs1_mcs_mat1_3_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_6611, shiftr_out[112]}), .c ({new_AGEMA_signal_7810, mcs1_mcs_mat1_3_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_6768, mcs1_mcs_mat1_3_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_7434, mcs1_mcs_mat1_3_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_7435, mcs1_mcs_mat1_3_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[315]), .c ({new_AGEMA_signal_6768, mcs1_mcs_mat1_3_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_9055, shiftr_out[83]}), .b ({new_AGEMA_signal_7617, shiftr_out[80]}), .c ({new_AGEMA_signal_9477, mcs1_mcs_mat1_3_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_9055, shiftr_out[83]}), .b ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_9478, mcs1_mcs_mat1_3_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({new_AGEMA_signal_7813, mcs1_mcs_mat1_3_mcs_out[87]}), .c ({new_AGEMA_signal_8295, mcs1_mcs_mat1_3_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_7303, shiftr_out[49]}), .c ({new_AGEMA_signal_7813, mcs1_mcs_mat1_3_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_7309, shiftr_out[17]}), .c ({new_AGEMA_signal_7816, mcs1_mcs_mat1_3_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[316]), .c ({new_AGEMA_signal_6769, mcs1_mcs_mat1_3_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_6770, mcs1_mcs_mat1_3_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_7046, mcs1_mcs_mat1_3_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[317]), .c ({new_AGEMA_signal_6770, mcs1_mcs_mat1_3_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_8301, mcs1_mcs_mat1_3_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_8780, mcs1_mcs_mat1_3_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7617, shiftr_out[80]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[318]), .c ({new_AGEMA_signal_8301, mcs1_mcs_mat1_3_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[319]), .c ({new_AGEMA_signal_6771, mcs1_mcs_mat1_3_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_6772, mcs1_mcs_mat1_3_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7309, shiftr_out[17]}), .c ({new_AGEMA_signal_7823, mcs1_mcs_mat1_3_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[320]), .c ({new_AGEMA_signal_6772, mcs1_mcs_mat1_3_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_8788, mcs1_mcs_mat1_3_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_6773, mcs1_mcs_mat1_3_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_9192, mcs1_mcs_mat1_3_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_8307, mcs1_mcs_mat1_3_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_8788, mcs1_mcs_mat1_3_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_7825, mcs1_mcs_mat1_3_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8307, mcs1_mcs_mat1_3_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_7825, mcs1_mcs_mat1_3_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[321]), .c ({new_AGEMA_signal_6773, mcs1_mcs_mat1_3_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_9715, mcs1_mcs_mat1_3_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_8789, mcs1_mcs_mat1_3_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_9941, mcs1_mcs_mat1_3_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_8308, mcs1_mcs_mat1_3_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_7617, shiftr_out[80]}), .c ({new_AGEMA_signal_8789, mcs1_mcs_mat1_3_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_7617, shiftr_out[80]}), .c ({new_AGEMA_signal_8790, mcs1_mcs_mat1_3_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_9055, shiftr_out[83]}), .c ({new_AGEMA_signal_9715, mcs1_mcs_mat1_3_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_8308, mcs1_mcs_mat1_3_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_9716, mcs1_mcs_mat1_3_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7617, shiftr_out[80]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[322]), .c ({new_AGEMA_signal_8308, mcs1_mcs_mat1_3_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_7303, shiftr_out[49]}), .b ({new_AGEMA_signal_6774, mcs1_mcs_mat1_3_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_7829, mcs1_mcs_mat1_3_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[323]), .c ({new_AGEMA_signal_6774, mcs1_mcs_mat1_3_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({new_AGEMA_signal_7831, mcs1_mcs_mat1_3_mcs_out[51]}), .c ({new_AGEMA_signal_8311, mcs1_mcs_mat1_3_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_7309, shiftr_out[17]}), .c ({new_AGEMA_signal_7831, mcs1_mcs_mat1_3_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_6775, mcs1_mcs_mat1_3_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_7444, mcs1_mcs_mat1_3_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[324]), .c ({new_AGEMA_signal_6775, mcs1_mcs_mat1_3_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_9718, mcs1_mcs_mat1_3_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_9945, mcs1_mcs_mat1_3_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_7617, shiftr_out[80]}), .b ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_9718, mcs1_mcs_mat1_3_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_9483, mcs1_mcs_mat1_3_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_9719, mcs1_mcs_mat1_3_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_9055, shiftr_out[83]}), .c ({new_AGEMA_signal_9483, mcs1_mcs_mat1_3_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7617, shiftr_out[80]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[325]), .c ({new_AGEMA_signal_8313, mcs1_mcs_mat1_3_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({new_AGEMA_signal_6776, mcs1_mcs_mat1_3_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_7446, mcs1_mcs_mat1_3_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_7303, shiftr_out[49]}), .b ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_7835, mcs1_mcs_mat1_3_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[326]), .c ({new_AGEMA_signal_6776, mcs1_mcs_mat1_3_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_8798, mcs1_mcs_mat1_3_mcs_out[35]}), .b ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_9198, mcs1_mcs_mat1_3_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_8317, mcs1_mcs_mat1_3_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_6777, mcs1_mcs_mat1_3_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_8798, mcs1_mcs_mat1_3_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_7837, mcs1_mcs_mat1_3_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_6697, shiftr_out[18]}), .c ({new_AGEMA_signal_8317, mcs1_mcs_mat1_3_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_7309, shiftr_out[17]}), .c ({new_AGEMA_signal_7837, mcs1_mcs_mat1_3_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[327]), .c ({new_AGEMA_signal_6777, mcs1_mcs_mat1_3_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_6778, mcs1_mcs_mat1_3_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_7055, mcs1_mcs_mat1_3_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({new_AGEMA_signal_7839, mcs1_mcs_mat1_3_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_8319, mcs1_mcs_mat1_3_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_6778, mcs1_mcs_mat1_3_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_7839, mcs1_mcs_mat1_3_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[328]), .c ({new_AGEMA_signal_6778, mcs1_mcs_mat1_3_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7617, shiftr_out[80]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[329]), .c ({new_AGEMA_signal_8321, mcs1_mcs_mat1_3_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[330]), .c ({new_AGEMA_signal_6779, mcs1_mcs_mat1_3_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_7452, mcs1_mcs_mat1_3_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_7845, mcs1_mcs_mat1_3_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_7452, mcs1_mcs_mat1_3_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_7309, shiftr_out[17]}), .c ({new_AGEMA_signal_7847, mcs1_mcs_mat1_3_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[331]), .c ({new_AGEMA_signal_6780, mcs1_mcs_mat1_3_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[332]), .c ({new_AGEMA_signal_6781, mcs1_mcs_mat1_3_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7617, shiftr_out[80]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[333]), .c ({new_AGEMA_signal_8331, mcs1_mcs_mat1_3_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_6782, mcs1_mcs_mat1_3_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_7455, mcs1_mcs_mat1_3_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_6782, mcs1_mcs_mat1_3_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_7060, mcs1_mcs_mat1_3_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[334]), .c ({new_AGEMA_signal_6782, mcs1_mcs_mat1_3_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_7853, mcs1_mcs_mat1_3_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_6783, mcs1_mcs_mat1_3_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8333, mcs1_mcs_mat1_3_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_7853, mcs1_mcs_mat1_3_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7309, shiftr_out[17]}), .c ({new_AGEMA_signal_8335, mcs1_mcs_mat1_3_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_7457, mcs1_mcs_mat1_3_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_7853, mcs1_mcs_mat1_3_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_7457, mcs1_mcs_mat1_3_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_7309, shiftr_out[17]}), .c ({new_AGEMA_signal_7854, mcs1_mcs_mat1_3_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[335]), .c ({new_AGEMA_signal_6783, mcs1_mcs_mat1_3_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U44 ( .a ({new_AGEMA_signal_7472, mcs1_mcs_mat1_4_mcs_out[90]}), .b ({new_AGEMA_signal_9738, mcs1_mcs_mat1_4_mcs_out[94]}), .c ({new_AGEMA_signal_9956, mcs1_mcs_mat1_4_n93}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({new_AGEMA_signal_7614, shiftr_out[108]}), .c ({new_AGEMA_signal_9507, mcs1_mcs_mat1_4_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_6616, shiftr_out[76]}), .b ({new_AGEMA_signal_6784, mcs1_mcs_mat1_4_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_7063, mcs1_mcs_mat1_4_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6616, shiftr_out[76]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[336]), .c ({new_AGEMA_signal_6784, mcs1_mcs_mat1_4_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_7461, mcs1_mcs_mat1_4_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_7858, mcs1_mcs_mat1_4_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_6785, mcs1_mcs_mat1_4_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_7461, mcs1_mcs_mat1_4_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[337]), .c ({new_AGEMA_signal_6785, mcs1_mcs_mat1_4_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_6786, mcs1_mcs_mat1_4_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_7862, mcs1_mcs_mat1_4_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8341, mcs1_mcs_mat1_4_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_7066, mcs1_mcs_mat1_4_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_7464, mcs1_mcs_mat1_4_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_6696, shiftr_out[14]}), .c ({new_AGEMA_signal_7066, mcs1_mcs_mat1_4_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_7308, shiftr_out[13]}), .b ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_7862, mcs1_mcs_mat1_4_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[338]), .c ({new_AGEMA_signal_6786, mcs1_mcs_mat1_4_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_9735, mcs1_mcs_mat1_4_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_9961, mcs1_mcs_mat1_4_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_8344, mcs1_mcs_mat1_4_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_9735, mcs1_mcs_mat1_4_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[339]), .c ({new_AGEMA_signal_8344, mcs1_mcs_mat1_4_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6616, shiftr_out[76]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[340]), .c ({new_AGEMA_signal_6787, mcs1_mcs_mat1_4_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({new_AGEMA_signal_7468, mcs1_mcs_mat1_4_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_7866, mcs1_mcs_mat1_4_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_6788, mcs1_mcs_mat1_4_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_7468, mcs1_mcs_mat1_4_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_7302, shiftr_out[45]}), .b ({new_AGEMA_signal_6690, shiftr_out[46]}), .c ({new_AGEMA_signal_7867, mcs1_mcs_mat1_4_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[341]), .c ({new_AGEMA_signal_6788, mcs1_mcs_mat1_4_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_6789, mcs1_mcs_mat1_4_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_7470, mcs1_mcs_mat1_4_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_6789, mcs1_mcs_mat1_4_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .c ({new_AGEMA_signal_7070, mcs1_mcs_mat1_4_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[342]), .c ({new_AGEMA_signal_6789, mcs1_mcs_mat1_4_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_9510, mcs1_mcs_mat1_4_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_7614, shiftr_out[108]}), .c ({new_AGEMA_signal_9738, mcs1_mcs_mat1_4_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_8351, mcs1_mcs_mat1_4_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_9510, mcs1_mcs_mat1_4_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_9511, mcs1_mcs_mat1_4_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[343]), .c ({new_AGEMA_signal_8351, mcs1_mcs_mat1_4_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_7230, shiftr_out[79]}), .b ({new_AGEMA_signal_6616, shiftr_out[76]}), .c ({new_AGEMA_signal_7472, mcs1_mcs_mat1_4_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_7230, shiftr_out[79]}), .b ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_7473, mcs1_mcs_mat1_4_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({new_AGEMA_signal_7871, mcs1_mcs_mat1_4_mcs_out[87]}), .c ({new_AGEMA_signal_8352, mcs1_mcs_mat1_4_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_7302, shiftr_out[45]}), .c ({new_AGEMA_signal_7871, mcs1_mcs_mat1_4_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_7308, shiftr_out[13]}), .c ({new_AGEMA_signal_7874, mcs1_mcs_mat1_4_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[344]), .c ({new_AGEMA_signal_6790, mcs1_mcs_mat1_4_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_8357, mcs1_mcs_mat1_4_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_8840, mcs1_mcs_mat1_4_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[345]), .c ({new_AGEMA_signal_8357, mcs1_mcs_mat1_4_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_6791, mcs1_mcs_mat1_4_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_7073, mcs1_mcs_mat1_4_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6616, shiftr_out[76]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[346]), .c ({new_AGEMA_signal_6791, mcs1_mcs_mat1_4_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[347]), .c ({new_AGEMA_signal_6792, mcs1_mcs_mat1_4_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_6793, mcs1_mcs_mat1_4_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7308, shiftr_out[13]}), .c ({new_AGEMA_signal_7882, mcs1_mcs_mat1_4_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[348]), .c ({new_AGEMA_signal_6793, mcs1_mcs_mat1_4_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_10183, mcs1_mcs_mat1_4_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_8363, mcs1_mcs_mat1_4_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_10423, mcs1_mcs_mat1_4_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_9967, mcs1_mcs_mat1_4_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_10183, mcs1_mcs_mat1_4_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_9743, mcs1_mcs_mat1_4_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_9967, mcs1_mcs_mat1_4_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_9743, mcs1_mcs_mat1_4_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[349]), .c ({new_AGEMA_signal_8363, mcs1_mcs_mat1_4_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_7885, mcs1_mcs_mat1_4_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_7077, mcs1_mcs_mat1_4_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_8364, mcs1_mcs_mat1_4_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_6794, mcs1_mcs_mat1_4_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_6616, shiftr_out[76]}), .c ({new_AGEMA_signal_7077, mcs1_mcs_mat1_4_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_6616, shiftr_out[76]}), .c ({new_AGEMA_signal_7078, mcs1_mcs_mat1_4_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_7230, shiftr_out[79]}), .c ({new_AGEMA_signal_7885, mcs1_mcs_mat1_4_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_6794, mcs1_mcs_mat1_4_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_7886, mcs1_mcs_mat1_4_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6616, shiftr_out[76]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[350]), .c ({new_AGEMA_signal_6794, mcs1_mcs_mat1_4_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_7302, shiftr_out[45]}), .b ({new_AGEMA_signal_6795, mcs1_mcs_mat1_4_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_7890, mcs1_mcs_mat1_4_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[351]), .c ({new_AGEMA_signal_6795, mcs1_mcs_mat1_4_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({new_AGEMA_signal_7892, mcs1_mcs_mat1_4_mcs_out[51]}), .c ({new_AGEMA_signal_8369, mcs1_mcs_mat1_4_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_7308, shiftr_out[13]}), .c ({new_AGEMA_signal_7892, mcs1_mcs_mat1_4_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_8370, mcs1_mcs_mat1_4_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_9516, mcs1_mcs_mat1_4_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[352]), .c ({new_AGEMA_signal_8370, mcs1_mcs_mat1_4_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_7893, mcs1_mcs_mat1_4_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_8372, mcs1_mcs_mat1_4_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_6616, shiftr_out[76]}), .b ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_7893, mcs1_mcs_mat1_4_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_7481, mcs1_mcs_mat1_4_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_7894, mcs1_mcs_mat1_4_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_7230, shiftr_out[79]}), .c ({new_AGEMA_signal_7481, mcs1_mcs_mat1_4_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6616, shiftr_out[76]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[353]), .c ({new_AGEMA_signal_6796, mcs1_mcs_mat1_4_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({new_AGEMA_signal_6797, mcs1_mcs_mat1_4_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_7483, mcs1_mcs_mat1_4_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_7302, shiftr_out[45]}), .b ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_7897, mcs1_mcs_mat1_4_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[354]), .c ({new_AGEMA_signal_6797, mcs1_mcs_mat1_4_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_8859, mcs1_mcs_mat1_4_mcs_out[35]}), .b ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_9232, mcs1_mcs_mat1_4_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_8378, mcs1_mcs_mat1_4_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_6798, mcs1_mcs_mat1_4_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_8859, mcs1_mcs_mat1_4_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_7899, mcs1_mcs_mat1_4_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_6696, shiftr_out[14]}), .c ({new_AGEMA_signal_8378, mcs1_mcs_mat1_4_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_7308, shiftr_out[13]}), .c ({new_AGEMA_signal_7899, mcs1_mcs_mat1_4_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[355]), .c ({new_AGEMA_signal_6798, mcs1_mcs_mat1_4_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_8379, mcs1_mcs_mat1_4_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({new_AGEMA_signal_9747, mcs1_mcs_mat1_4_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_9970, mcs1_mcs_mat1_4_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_8379, mcs1_mcs_mat1_4_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_9747, mcs1_mcs_mat1_4_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[356]), .c ({new_AGEMA_signal_8379, mcs1_mcs_mat1_4_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6616, shiftr_out[76]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[357]), .c ({new_AGEMA_signal_6799, mcs1_mcs_mat1_4_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[358]), .c ({new_AGEMA_signal_6800, mcs1_mcs_mat1_4_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_7489, mcs1_mcs_mat1_4_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_7907, mcs1_mcs_mat1_4_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_7489, mcs1_mcs_mat1_4_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_7308, shiftr_out[13]}), .c ({new_AGEMA_signal_7909, mcs1_mcs_mat1_4_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[359]), .c ({new_AGEMA_signal_6801, mcs1_mcs_mat1_4_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[360]), .c ({new_AGEMA_signal_8389, mcs1_mcs_mat1_4_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6616, shiftr_out[76]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[361]), .c ({new_AGEMA_signal_6802, mcs1_mcs_mat1_4_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_6803, mcs1_mcs_mat1_4_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_7493, mcs1_mcs_mat1_4_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_6803, mcs1_mcs_mat1_4_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_7088, mcs1_mcs_mat1_4_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[362]), .c ({new_AGEMA_signal_6803, mcs1_mcs_mat1_4_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_7915, mcs1_mcs_mat1_4_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_6804, mcs1_mcs_mat1_4_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8393, mcs1_mcs_mat1_4_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_7915, mcs1_mcs_mat1_4_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7308, shiftr_out[13]}), .c ({new_AGEMA_signal_8395, mcs1_mcs_mat1_4_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_7495, mcs1_mcs_mat1_4_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_7915, mcs1_mcs_mat1_4_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_7495, mcs1_mcs_mat1_4_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_7308, shiftr_out[13]}), .c ({new_AGEMA_signal_7916, mcs1_mcs_mat1_4_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[363]), .c ({new_AGEMA_signal_6804, mcs1_mcs_mat1_4_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U44 ( .a ({new_AGEMA_signal_7511, mcs1_mcs_mat1_5_mcs_out[90]}), .b ({new_AGEMA_signal_7931, mcs1_mcs_mat1_5_mcs_out[94]}), .c ({new_AGEMA_signal_8398, mcs1_mcs_mat1_5_n93}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({new_AGEMA_signal_6610, shiftr_out[104]}), .c ({new_AGEMA_signal_7497, mcs1_mcs_mat1_5_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_6615, shiftr_out[72]}), .b ({new_AGEMA_signal_6805, mcs1_mcs_mat1_5_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_7091, mcs1_mcs_mat1_5_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6615, shiftr_out[72]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[364]), .c ({new_AGEMA_signal_6805, mcs1_mcs_mat1_5_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_7500, mcs1_mcs_mat1_5_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_7920, mcs1_mcs_mat1_5_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_6806, mcs1_mcs_mat1_5_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_7500, mcs1_mcs_mat1_5_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[365]), .c ({new_AGEMA_signal_6806, mcs1_mcs_mat1_5_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_8404, mcs1_mcs_mat1_5_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9759, mcs1_mcs_mat1_5_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_9980, mcs1_mcs_mat1_5_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_8884, mcs1_mcs_mat1_5_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_9536, mcs1_mcs_mat1_5_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_8100, shiftr_out[10]}), .c ({new_AGEMA_signal_8884, mcs1_mcs_mat1_5_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_9362, shiftr_out[9]}), .b ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_9759, mcs1_mcs_mat1_5_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[366]), .c ({new_AGEMA_signal_8404, mcs1_mcs_mat1_5_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_7923, mcs1_mcs_mat1_5_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_8405, mcs1_mcs_mat1_5_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_6807, mcs1_mcs_mat1_5_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_7923, mcs1_mcs_mat1_5_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[367]), .c ({new_AGEMA_signal_6807, mcs1_mcs_mat1_5_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6615, shiftr_out[72]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[368]), .c ({new_AGEMA_signal_6808, mcs1_mcs_mat1_5_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({new_AGEMA_signal_7506, mcs1_mcs_mat1_5_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_7927, mcs1_mcs_mat1_5_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_6809, mcs1_mcs_mat1_5_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_7506, mcs1_mcs_mat1_5_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_7301, shiftr_out[41]}), .b ({new_AGEMA_signal_6689, shiftr_out[42]}), .c ({new_AGEMA_signal_7928, mcs1_mcs_mat1_5_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[369]), .c ({new_AGEMA_signal_6809, mcs1_mcs_mat1_5_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_8412, mcs1_mcs_mat1_5_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_9538, mcs1_mcs_mat1_5_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_8412, mcs1_mcs_mat1_5_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .c ({new_AGEMA_signal_8894, mcs1_mcs_mat1_5_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[370]), .c ({new_AGEMA_signal_8412, mcs1_mcs_mat1_5_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_7508, mcs1_mcs_mat1_5_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_6610, shiftr_out[104]}), .c ({new_AGEMA_signal_7931, mcs1_mcs_mat1_5_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_6810, mcs1_mcs_mat1_5_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_7508, mcs1_mcs_mat1_5_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_7509, mcs1_mcs_mat1_5_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[371]), .c ({new_AGEMA_signal_6810, mcs1_mcs_mat1_5_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_7229, shiftr_out[75]}), .b ({new_AGEMA_signal_6615, shiftr_out[72]}), .c ({new_AGEMA_signal_7511, mcs1_mcs_mat1_5_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_7229, shiftr_out[75]}), .b ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_7512, mcs1_mcs_mat1_5_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({new_AGEMA_signal_7934, mcs1_mcs_mat1_5_mcs_out[87]}), .c ({new_AGEMA_signal_8414, mcs1_mcs_mat1_5_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_7301, shiftr_out[41]}), .c ({new_AGEMA_signal_7934, mcs1_mcs_mat1_5_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_9362, shiftr_out[9]}), .c ({new_AGEMA_signal_9764, mcs1_mcs_mat1_5_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[372]), .c ({new_AGEMA_signal_8415, mcs1_mcs_mat1_5_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_6811, mcs1_mcs_mat1_5_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_7098, mcs1_mcs_mat1_5_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[373]), .c ({new_AGEMA_signal_6811, mcs1_mcs_mat1_5_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_6812, mcs1_mcs_mat1_5_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_7100, mcs1_mcs_mat1_5_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6615, shiftr_out[72]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[374]), .c ({new_AGEMA_signal_6812, mcs1_mcs_mat1_5_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[375]), .c ({new_AGEMA_signal_6813, mcs1_mcs_mat1_5_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_8421, mcs1_mcs_mat1_5_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_9362, shiftr_out[9]}), .c ({new_AGEMA_signal_9766, mcs1_mcs_mat1_5_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[376]), .c ({new_AGEMA_signal_8421, mcs1_mcs_mat1_5_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_8908, mcs1_mcs_mat1_5_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_6814, mcs1_mcs_mat1_5_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_9266, mcs1_mcs_mat1_5_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_8424, mcs1_mcs_mat1_5_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_8908, mcs1_mcs_mat1_5_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_7943, mcs1_mcs_mat1_5_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8424, mcs1_mcs_mat1_5_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_7943, mcs1_mcs_mat1_5_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[377]), .c ({new_AGEMA_signal_6814, mcs1_mcs_mat1_5_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_7946, mcs1_mcs_mat1_5_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_7104, mcs1_mcs_mat1_5_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_8425, mcs1_mcs_mat1_5_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_6815, mcs1_mcs_mat1_5_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_6615, shiftr_out[72]}), .c ({new_AGEMA_signal_7104, mcs1_mcs_mat1_5_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_6615, shiftr_out[72]}), .c ({new_AGEMA_signal_7105, mcs1_mcs_mat1_5_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_7229, shiftr_out[75]}), .c ({new_AGEMA_signal_7946, mcs1_mcs_mat1_5_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_6815, mcs1_mcs_mat1_5_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_7947, mcs1_mcs_mat1_5_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6615, shiftr_out[72]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[378]), .c ({new_AGEMA_signal_6815, mcs1_mcs_mat1_5_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_7301, shiftr_out[41]}), .b ({new_AGEMA_signal_6816, mcs1_mcs_mat1_5_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_7951, mcs1_mcs_mat1_5_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[379]), .c ({new_AGEMA_signal_6816, mcs1_mcs_mat1_5_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({new_AGEMA_signal_9768, mcs1_mcs_mat1_5_mcs_out[51]}), .c ({new_AGEMA_signal_9989, mcs1_mcs_mat1_5_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_9362, shiftr_out[9]}), .c ({new_AGEMA_signal_9768, mcs1_mcs_mat1_5_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_6817, mcs1_mcs_mat1_5_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_7520, mcs1_mcs_mat1_5_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[380]), .c ({new_AGEMA_signal_6817, mcs1_mcs_mat1_5_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_7955, mcs1_mcs_mat1_5_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_8432, mcs1_mcs_mat1_5_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_6615, shiftr_out[72]}), .b ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_7955, mcs1_mcs_mat1_5_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_7522, mcs1_mcs_mat1_5_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_7956, mcs1_mcs_mat1_5_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_7229, shiftr_out[75]}), .c ({new_AGEMA_signal_7522, mcs1_mcs_mat1_5_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6615, shiftr_out[72]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[381]), .c ({new_AGEMA_signal_6818, mcs1_mcs_mat1_5_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({new_AGEMA_signal_6819, mcs1_mcs_mat1_5_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_7524, mcs1_mcs_mat1_5_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_7301, shiftr_out[41]}), .b ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_7959, mcs1_mcs_mat1_5_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[382]), .c ({new_AGEMA_signal_6819, mcs1_mcs_mat1_5_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_10211, mcs1_mcs_mat1_5_mcs_out[35]}), .b ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_10451, mcs1_mcs_mat1_5_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_9991, mcs1_mcs_mat1_5_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_8437, mcs1_mcs_mat1_5_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_10211, mcs1_mcs_mat1_5_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_9769, mcs1_mcs_mat1_5_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_8100, shiftr_out[10]}), .c ({new_AGEMA_signal_9991, mcs1_mcs_mat1_5_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_9362, shiftr_out[9]}), .c ({new_AGEMA_signal_9769, mcs1_mcs_mat1_5_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[383]), .c ({new_AGEMA_signal_8437, mcs1_mcs_mat1_5_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_6820, mcs1_mcs_mat1_5_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_7111, mcs1_mcs_mat1_5_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({new_AGEMA_signal_7961, mcs1_mcs_mat1_5_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_8439, mcs1_mcs_mat1_5_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_6820, mcs1_mcs_mat1_5_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_7961, mcs1_mcs_mat1_5_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[384]), .c ({new_AGEMA_signal_6820, mcs1_mcs_mat1_5_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6615, shiftr_out[72]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[385]), .c ({new_AGEMA_signal_6821, mcs1_mcs_mat1_5_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[386]), .c ({new_AGEMA_signal_6822, mcs1_mcs_mat1_5_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_9544, mcs1_mcs_mat1_5_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_9771, mcs1_mcs_mat1_5_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_9544, mcs1_mcs_mat1_5_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_9362, shiftr_out[9]}), .c ({new_AGEMA_signal_9773, mcs1_mcs_mat1_5_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[387]), .c ({new_AGEMA_signal_8447, mcs1_mcs_mat1_5_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[388]), .c ({new_AGEMA_signal_6823, mcs1_mcs_mat1_5_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6615, shiftr_out[72]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[389]), .c ({new_AGEMA_signal_6824, mcs1_mcs_mat1_5_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_6825, mcs1_mcs_mat1_5_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_7533, mcs1_mcs_mat1_5_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_6825, mcs1_mcs_mat1_5_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_7117, mcs1_mcs_mat1_5_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[390]), .c ({new_AGEMA_signal_6825, mcs1_mcs_mat1_5_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_9777, mcs1_mcs_mat1_5_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8454, mcs1_mcs_mat1_5_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_9995, mcs1_mcs_mat1_5_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_9777, mcs1_mcs_mat1_5_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_9362, shiftr_out[9]}), .c ({new_AGEMA_signal_9997, mcs1_mcs_mat1_5_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_9548, mcs1_mcs_mat1_5_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_9777, mcs1_mcs_mat1_5_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_9548, mcs1_mcs_mat1_5_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_9362, shiftr_out[9]}), .c ({new_AGEMA_signal_9778, mcs1_mcs_mat1_5_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[391]), .c ({new_AGEMA_signal_8454, mcs1_mcs_mat1_5_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U44 ( .a ({new_AGEMA_signal_7548, mcs1_mcs_mat1_6_mcs_out[90]}), .b ({new_AGEMA_signal_7985, mcs1_mcs_mat1_6_mcs_out[94]}), .c ({new_AGEMA_signal_8456, mcs1_mcs_mat1_6_n93}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({new_AGEMA_signal_6609, shiftr_out[100]}), .c ({new_AGEMA_signal_7535, mcs1_mcs_mat1_6_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_6614, shiftr_out[68]}), .b ({new_AGEMA_signal_6826, mcs1_mcs_mat1_6_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_7119, mcs1_mcs_mat1_6_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6614, shiftr_out[68]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[392]), .c ({new_AGEMA_signal_6826, mcs1_mcs_mat1_6_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_9564, mcs1_mcs_mat1_6_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_9784, mcs1_mcs_mat1_6_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_8460, mcs1_mcs_mat1_6_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_9564, mcs1_mcs_mat1_6_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[393]), .c ({new_AGEMA_signal_8460, mcs1_mcs_mat1_6_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_6827, mcs1_mcs_mat1_6_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_7978, mcs1_mcs_mat1_6_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8461, mcs1_mcs_mat1_6_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_7121, mcs1_mcs_mat1_6_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_7538, mcs1_mcs_mat1_6_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_6695, shiftr_out[6]}), .c ({new_AGEMA_signal_7121, mcs1_mcs_mat1_6_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_7307, shiftr_out[5]}), .b ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_7978, mcs1_mcs_mat1_6_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[394]), .c ({new_AGEMA_signal_6827, mcs1_mcs_mat1_6_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_7980, mcs1_mcs_mat1_6_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_8464, mcs1_mcs_mat1_6_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_6828, mcs1_mcs_mat1_6_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_7980, mcs1_mcs_mat1_6_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[395]), .c ({new_AGEMA_signal_6828, mcs1_mcs_mat1_6_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6614, shiftr_out[68]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[396]), .c ({new_AGEMA_signal_6829, mcs1_mcs_mat1_6_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({new_AGEMA_signal_9567, mcs1_mcs_mat1_6_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_9787, mcs1_mcs_mat1_6_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_8468, mcs1_mcs_mat1_6_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_9567, mcs1_mcs_mat1_6_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_9360, shiftr_out[37]}), .b ({new_AGEMA_signal_8098, shiftr_out[38]}), .c ({new_AGEMA_signal_9788, mcs1_mcs_mat1_6_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[397]), .c ({new_AGEMA_signal_8468, mcs1_mcs_mat1_6_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_6830, mcs1_mcs_mat1_6_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_7543, mcs1_mcs_mat1_6_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_6830, mcs1_mcs_mat1_6_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .c ({new_AGEMA_signal_7125, mcs1_mcs_mat1_6_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[398]), .c ({new_AGEMA_signal_6830, mcs1_mcs_mat1_6_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_7545, mcs1_mcs_mat1_6_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_6609, shiftr_out[100]}), .c ({new_AGEMA_signal_7985, mcs1_mcs_mat1_6_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_6831, mcs1_mcs_mat1_6_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_7545, mcs1_mcs_mat1_6_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_7546, mcs1_mcs_mat1_6_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[399]), .c ({new_AGEMA_signal_6831, mcs1_mcs_mat1_6_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_7228, shiftr_out[71]}), .b ({new_AGEMA_signal_6614, shiftr_out[68]}), .c ({new_AGEMA_signal_7548, mcs1_mcs_mat1_6_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_7228, shiftr_out[71]}), .b ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_7549, mcs1_mcs_mat1_6_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({new_AGEMA_signal_9792, mcs1_mcs_mat1_6_mcs_out[87]}), .c ({new_AGEMA_signal_10009, mcs1_mcs_mat1_6_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_9360, shiftr_out[37]}), .c ({new_AGEMA_signal_9792, mcs1_mcs_mat1_6_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_7307, shiftr_out[5]}), .c ({new_AGEMA_signal_7990, mcs1_mcs_mat1_6_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[400]), .c ({new_AGEMA_signal_6832, mcs1_mcs_mat1_6_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_6833, mcs1_mcs_mat1_6_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_7129, mcs1_mcs_mat1_6_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[401]), .c ({new_AGEMA_signal_6833, mcs1_mcs_mat1_6_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_6834, mcs1_mcs_mat1_6_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_7131, mcs1_mcs_mat1_6_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6614, shiftr_out[68]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[402]), .c ({new_AGEMA_signal_6834, mcs1_mcs_mat1_6_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[403]), .c ({new_AGEMA_signal_8478, mcs1_mcs_mat1_6_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_6835, mcs1_mcs_mat1_6_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7307, shiftr_out[5]}), .c ({new_AGEMA_signal_7997, mcs1_mcs_mat1_6_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[404]), .c ({new_AGEMA_signal_6835, mcs1_mcs_mat1_6_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_8963, mcs1_mcs_mat1_6_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_6836, mcs1_mcs_mat1_6_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_9307, mcs1_mcs_mat1_6_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_8482, mcs1_mcs_mat1_6_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_8963, mcs1_mcs_mat1_6_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_7999, mcs1_mcs_mat1_6_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8482, mcs1_mcs_mat1_6_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_7999, mcs1_mcs_mat1_6_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[405]), .c ({new_AGEMA_signal_6836, mcs1_mcs_mat1_6_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_8002, mcs1_mcs_mat1_6_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_7135, mcs1_mcs_mat1_6_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_8483, mcs1_mcs_mat1_6_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_6837, mcs1_mcs_mat1_6_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_6614, shiftr_out[68]}), .c ({new_AGEMA_signal_7135, mcs1_mcs_mat1_6_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_6614, shiftr_out[68]}), .c ({new_AGEMA_signal_7136, mcs1_mcs_mat1_6_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_7228, shiftr_out[71]}), .c ({new_AGEMA_signal_8002, mcs1_mcs_mat1_6_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_6837, mcs1_mcs_mat1_6_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_8003, mcs1_mcs_mat1_6_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6614, shiftr_out[68]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[406]), .c ({new_AGEMA_signal_6837, mcs1_mcs_mat1_6_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_9360, shiftr_out[37]}), .b ({new_AGEMA_signal_8486, mcs1_mcs_mat1_6_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_9798, mcs1_mcs_mat1_6_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[407]), .c ({new_AGEMA_signal_8486, mcs1_mcs_mat1_6_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({new_AGEMA_signal_8005, mcs1_mcs_mat1_6_mcs_out[51]}), .c ({new_AGEMA_signal_8487, mcs1_mcs_mat1_6_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_7307, shiftr_out[5]}), .c ({new_AGEMA_signal_8005, mcs1_mcs_mat1_6_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_6838, mcs1_mcs_mat1_6_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_7556, mcs1_mcs_mat1_6_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[408]), .c ({new_AGEMA_signal_6838, mcs1_mcs_mat1_6_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_8008, mcs1_mcs_mat1_6_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_8490, mcs1_mcs_mat1_6_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_6614, shiftr_out[68]}), .b ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_8008, mcs1_mcs_mat1_6_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_7558, mcs1_mcs_mat1_6_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_8009, mcs1_mcs_mat1_6_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_7228, shiftr_out[71]}), .c ({new_AGEMA_signal_7558, mcs1_mcs_mat1_6_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6614, shiftr_out[68]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[409]), .c ({new_AGEMA_signal_6839, mcs1_mcs_mat1_6_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({new_AGEMA_signal_8493, mcs1_mcs_mat1_6_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9575, mcs1_mcs_mat1_6_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_9360, shiftr_out[37]}), .b ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_9801, mcs1_mcs_mat1_6_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[410]), .c ({new_AGEMA_signal_8493, mcs1_mcs_mat1_6_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_8971, mcs1_mcs_mat1_6_mcs_out[35]}), .b ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_9310, mcs1_mcs_mat1_6_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_8495, mcs1_mcs_mat1_6_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_6840, mcs1_mcs_mat1_6_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_8971, mcs1_mcs_mat1_6_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_8011, mcs1_mcs_mat1_6_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_6695, shiftr_out[6]}), .c ({new_AGEMA_signal_8495, mcs1_mcs_mat1_6_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_7307, shiftr_out[5]}), .c ({new_AGEMA_signal_8011, mcs1_mcs_mat1_6_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[411]), .c ({new_AGEMA_signal_6840, mcs1_mcs_mat1_6_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_6841, mcs1_mcs_mat1_6_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_7141, mcs1_mcs_mat1_6_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({new_AGEMA_signal_8013, mcs1_mcs_mat1_6_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_8497, mcs1_mcs_mat1_6_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_6841, mcs1_mcs_mat1_6_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_8013, mcs1_mcs_mat1_6_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[412]), .c ({new_AGEMA_signal_6841, mcs1_mcs_mat1_6_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6614, shiftr_out[68]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[413]), .c ({new_AGEMA_signal_6842, mcs1_mcs_mat1_6_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[414]), .c ({new_AGEMA_signal_8502, mcs1_mcs_mat1_6_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_7563, mcs1_mcs_mat1_6_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_8019, mcs1_mcs_mat1_6_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_7563, mcs1_mcs_mat1_6_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_7307, shiftr_out[5]}), .c ({new_AGEMA_signal_8021, mcs1_mcs_mat1_6_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[415]), .c ({new_AGEMA_signal_6843, mcs1_mcs_mat1_6_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[416]), .c ({new_AGEMA_signal_6844, mcs1_mcs_mat1_6_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6614, shiftr_out[68]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[417]), .c ({new_AGEMA_signal_6845, mcs1_mcs_mat1_6_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_8511, mcs1_mcs_mat1_6_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_9581, mcs1_mcs_mat1_6_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_8511, mcs1_mcs_mat1_6_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_8985, mcs1_mcs_mat1_6_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[418]), .c ({new_AGEMA_signal_8511, mcs1_mcs_mat1_6_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_8028, mcs1_mcs_mat1_6_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_6846, mcs1_mcs_mat1_6_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8512, mcs1_mcs_mat1_6_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_8028, mcs1_mcs_mat1_6_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7307, shiftr_out[5]}), .c ({new_AGEMA_signal_8514, mcs1_mcs_mat1_6_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_7568, mcs1_mcs_mat1_6_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_8028, mcs1_mcs_mat1_6_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_7568, mcs1_mcs_mat1_6_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_7307, shiftr_out[5]}), .c ({new_AGEMA_signal_8029, mcs1_mcs_mat1_6_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[419]), .c ({new_AGEMA_signal_6846, mcs1_mcs_mat1_6_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U44 ( .a ({new_AGEMA_signal_9604, mcs1_mcs_mat1_7_mcs_out[90]}), .b ({new_AGEMA_signal_8044, mcs1_mcs_mat1_7_mcs_out[94]}), .c ({new_AGEMA_signal_9810, mcs1_mcs_mat1_7_n93}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({new_AGEMA_signal_6608, shiftr_out[96]}), .c ({new_AGEMA_signal_7570, mcs1_mcs_mat1_7_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_7616, shiftr_out[64]}), .b ({new_AGEMA_signal_8516, mcs1_mcs_mat1_7_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8996, mcs1_mcs_mat1_7_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7616, shiftr_out[64]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[420]), .c ({new_AGEMA_signal_8516, mcs1_mcs_mat1_7_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_7571, mcs1_mcs_mat1_7_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_8031, mcs1_mcs_mat1_7_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_6847, mcs1_mcs_mat1_7_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_7571, mcs1_mcs_mat1_7_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[421]), .c ({new_AGEMA_signal_6847, mcs1_mcs_mat1_7_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_6848, mcs1_mcs_mat1_7_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_8035, mcs1_mcs_mat1_7_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8519, mcs1_mcs_mat1_7_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_7149, mcs1_mcs_mat1_7_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_7574, mcs1_mcs_mat1_7_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_6694, shiftr_out[2]}), .c ({new_AGEMA_signal_7149, mcs1_mcs_mat1_7_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_7306, shiftr_out[1]}), .b ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_8035, mcs1_mcs_mat1_7_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[422]), .c ({new_AGEMA_signal_6848, mcs1_mcs_mat1_7_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_8037, mcs1_mcs_mat1_7_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_8522, mcs1_mcs_mat1_7_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_6849, mcs1_mcs_mat1_7_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_8037, mcs1_mcs_mat1_7_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[423]), .c ({new_AGEMA_signal_6849, mcs1_mcs_mat1_7_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7616, shiftr_out[64]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[424]), .c ({new_AGEMA_signal_8524, mcs1_mcs_mat1_7_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({new_AGEMA_signal_7577, mcs1_mcs_mat1_7_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_8039, mcs1_mcs_mat1_7_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_6850, mcs1_mcs_mat1_7_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_7577, mcs1_mcs_mat1_7_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_7300, shiftr_out[33]}), .b ({new_AGEMA_signal_6688, shiftr_out[34]}), .c ({new_AGEMA_signal_8040, mcs1_mcs_mat1_7_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[425]), .c ({new_AGEMA_signal_6850, mcs1_mcs_mat1_7_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_6851, mcs1_mcs_mat1_7_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_7579, mcs1_mcs_mat1_7_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_6851, mcs1_mcs_mat1_7_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .c ({new_AGEMA_signal_7153, mcs1_mcs_mat1_7_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[426]), .c ({new_AGEMA_signal_6851, mcs1_mcs_mat1_7_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_7581, mcs1_mcs_mat1_7_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_6608, shiftr_out[96]}), .c ({new_AGEMA_signal_8044, mcs1_mcs_mat1_7_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_6852, mcs1_mcs_mat1_7_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_7581, mcs1_mcs_mat1_7_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_7582, mcs1_mcs_mat1_7_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[427]), .c ({new_AGEMA_signal_6852, mcs1_mcs_mat1_7_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_9054, shiftr_out[67]}), .b ({new_AGEMA_signal_7616, shiftr_out[64]}), .c ({new_AGEMA_signal_9604, mcs1_mcs_mat1_7_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_9054, shiftr_out[67]}), .b ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_9605, mcs1_mcs_mat1_7_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({new_AGEMA_signal_8047, mcs1_mcs_mat1_7_mcs_out[87]}), .c ({new_AGEMA_signal_8530, mcs1_mcs_mat1_7_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_7300, shiftr_out[33]}), .c ({new_AGEMA_signal_8047, mcs1_mcs_mat1_7_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_7306, shiftr_out[1]}), .c ({new_AGEMA_signal_8050, mcs1_mcs_mat1_7_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[428]), .c ({new_AGEMA_signal_6853, mcs1_mcs_mat1_7_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_6854, mcs1_mcs_mat1_7_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_7157, mcs1_mcs_mat1_7_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[429]), .c ({new_AGEMA_signal_6854, mcs1_mcs_mat1_7_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_8536, mcs1_mcs_mat1_7_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_9014, mcs1_mcs_mat1_7_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7616, shiftr_out[64]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[430]), .c ({new_AGEMA_signal_8536, mcs1_mcs_mat1_7_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[431]), .c ({new_AGEMA_signal_6855, mcs1_mcs_mat1_7_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_6856, mcs1_mcs_mat1_7_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7306, shiftr_out[1]}), .c ({new_AGEMA_signal_8057, mcs1_mcs_mat1_7_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[432]), .c ({new_AGEMA_signal_6856, mcs1_mcs_mat1_7_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_9022, mcs1_mcs_mat1_7_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_6857, mcs1_mcs_mat1_7_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_9339, mcs1_mcs_mat1_7_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_8542, mcs1_mcs_mat1_7_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_9022, mcs1_mcs_mat1_7_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_8059, mcs1_mcs_mat1_7_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8542, mcs1_mcs_mat1_7_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_8059, mcs1_mcs_mat1_7_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[433]), .c ({new_AGEMA_signal_6857, mcs1_mcs_mat1_7_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_9824, mcs1_mcs_mat1_7_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_9023, mcs1_mcs_mat1_7_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_10034, mcs1_mcs_mat1_7_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_8543, mcs1_mcs_mat1_7_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_7616, shiftr_out[64]}), .c ({new_AGEMA_signal_9023, mcs1_mcs_mat1_7_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_7616, shiftr_out[64]}), .c ({new_AGEMA_signal_9024, mcs1_mcs_mat1_7_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_9054, shiftr_out[67]}), .c ({new_AGEMA_signal_9824, mcs1_mcs_mat1_7_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_8543, mcs1_mcs_mat1_7_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_9825, mcs1_mcs_mat1_7_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7616, shiftr_out[64]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[434]), .c ({new_AGEMA_signal_8543, mcs1_mcs_mat1_7_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_7300, shiftr_out[33]}), .b ({new_AGEMA_signal_6858, mcs1_mcs_mat1_7_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_8063, mcs1_mcs_mat1_7_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[435]), .c ({new_AGEMA_signal_6858, mcs1_mcs_mat1_7_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({new_AGEMA_signal_8065, mcs1_mcs_mat1_7_mcs_out[51]}), .c ({new_AGEMA_signal_8546, mcs1_mcs_mat1_7_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_7306, shiftr_out[1]}), .c ({new_AGEMA_signal_8065, mcs1_mcs_mat1_7_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_6859, mcs1_mcs_mat1_7_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_7591, mcs1_mcs_mat1_7_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[436]), .c ({new_AGEMA_signal_6859, mcs1_mcs_mat1_7_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_9827, mcs1_mcs_mat1_7_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_10038, mcs1_mcs_mat1_7_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_7616, shiftr_out[64]}), .b ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_9827, mcs1_mcs_mat1_7_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_9610, mcs1_mcs_mat1_7_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_9828, mcs1_mcs_mat1_7_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_9054, shiftr_out[67]}), .c ({new_AGEMA_signal_9610, mcs1_mcs_mat1_7_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7616, shiftr_out[64]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[437]), .c ({new_AGEMA_signal_8548, mcs1_mcs_mat1_7_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({new_AGEMA_signal_6860, mcs1_mcs_mat1_7_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_7593, mcs1_mcs_mat1_7_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_7300, shiftr_out[33]}), .b ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_8069, mcs1_mcs_mat1_7_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[438]), .c ({new_AGEMA_signal_6860, mcs1_mcs_mat1_7_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_9032, mcs1_mcs_mat1_7_mcs_out[35]}), .b ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_9345, mcs1_mcs_mat1_7_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_8552, mcs1_mcs_mat1_7_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_6861, mcs1_mcs_mat1_7_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_9032, mcs1_mcs_mat1_7_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_8071, mcs1_mcs_mat1_7_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_6694, shiftr_out[2]}), .c ({new_AGEMA_signal_8552, mcs1_mcs_mat1_7_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_7306, shiftr_out[1]}), .c ({new_AGEMA_signal_8071, mcs1_mcs_mat1_7_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[439]), .c ({new_AGEMA_signal_6861, mcs1_mcs_mat1_7_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_6862, mcs1_mcs_mat1_7_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_7166, mcs1_mcs_mat1_7_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({new_AGEMA_signal_8073, mcs1_mcs_mat1_7_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_8554, mcs1_mcs_mat1_7_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_6862, mcs1_mcs_mat1_7_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_8073, mcs1_mcs_mat1_7_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[440]), .c ({new_AGEMA_signal_6862, mcs1_mcs_mat1_7_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7616, shiftr_out[64]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[441]), .c ({new_AGEMA_signal_8556, mcs1_mcs_mat1_7_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[442]), .c ({new_AGEMA_signal_6863, mcs1_mcs_mat1_7_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_7599, mcs1_mcs_mat1_7_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_8079, mcs1_mcs_mat1_7_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_7599, mcs1_mcs_mat1_7_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_7306, shiftr_out[1]}), .c ({new_AGEMA_signal_8081, mcs1_mcs_mat1_7_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[443]), .c ({new_AGEMA_signal_6864, mcs1_mcs_mat1_7_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[444]), .c ({new_AGEMA_signal_6865, mcs1_mcs_mat1_7_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7616, shiftr_out[64]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[445]), .c ({new_AGEMA_signal_8566, mcs1_mcs_mat1_7_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_6866, mcs1_mcs_mat1_7_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_7602, mcs1_mcs_mat1_7_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_6866, mcs1_mcs_mat1_7_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_7171, mcs1_mcs_mat1_7_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[446]), .c ({new_AGEMA_signal_6866, mcs1_mcs_mat1_7_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_8087, mcs1_mcs_mat1_7_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_6867, mcs1_mcs_mat1_7_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8568, mcs1_mcs_mat1_7_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_8087, mcs1_mcs_mat1_7_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7306, shiftr_out[1]}), .c ({new_AGEMA_signal_8570, mcs1_mcs_mat1_7_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_7604, mcs1_mcs_mat1_7_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_8087, mcs1_mcs_mat1_7_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_7604, mcs1_mcs_mat1_7_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_7306, shiftr_out[1]}), .c ({new_AGEMA_signal_8088, mcs1_mcs_mat1_7_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[447]), .c ({new_AGEMA_signal_6867, mcs1_mcs_mat1_7_mcs_rom0_31_x0x4}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) U515 ( .a ({new_AGEMA_signal_10936, mcs_out[128]}), .b ({w0_s1[0], w0_s0[0]}), .c ({new_AGEMA_signal_10956, y0_1[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U516 ( .a ({new_AGEMA_signal_10459, mcs_out[228]}), .b ({w0_s1[100], w0_s0[100]}), .c ({new_AGEMA_signal_10514, y0_1[100]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U517 ( .a ({new_AGEMA_signal_10716, mcs_out[229]}), .b ({w0_s1[101], w0_s0[101]}), .c ({new_AGEMA_signal_10764, y0_1[101]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U518 ( .a ({new_AGEMA_signal_10924, mcs_out[230]}), .b ({w0_s1[102], w0_s0[102]}), .c ({new_AGEMA_signal_10957, y0_1[102]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U519 ( .a ({new_AGEMA_signal_10923, mcs_out[231]}), .b ({w0_s1[103], w0_s0[103]}), .c ({new_AGEMA_signal_10958, y0_1[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U520 ( .a ({new_AGEMA_signal_10915, mcs_out[232]}), .b ({w0_s1[104], w0_s0[104]}), .c ({new_AGEMA_signal_10959, y0_1[104]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U521 ( .a ({new_AGEMA_signal_10196, mcs_out[233]}), .b ({w0_s1[105], w0_s0[105]}), .c ({new_AGEMA_signal_10278, y0_1[105]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U522 ( .a ({new_AGEMA_signal_10434, mcs_out[234]}), .b ({w0_s1[106], w0_s0[106]}), .c ({new_AGEMA_signal_10515, y0_1[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U523 ( .a ({new_AGEMA_signal_10698, mcs_out[235]}), .b ({w0_s1[107], w0_s0[107]}), .c ({new_AGEMA_signal_10765, y0_1[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U524 ( .a ({new_AGEMA_signal_9731, mcs_out[236]}), .b ({w0_s1[108], w0_s0[108]}), .c ({new_AGEMA_signal_9838, y0_1[108]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U525 ( .a ({new_AGEMA_signal_9955, mcs_out[237]}), .b ({w0_s1[109], w0_s0[109]}), .c ({new_AGEMA_signal_10046, y0_1[109]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U526 ( .a ({new_AGEMA_signal_10704, mcs_out[138]}), .b ({w0_s1[10], w0_s0[10]}), .c ({new_AGEMA_signal_10766, y0_1[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U527 ( .a ({new_AGEMA_signal_9954, mcs_out[238]}), .b ({w0_s1[110], w0_s0[110]}), .c ({new_AGEMA_signal_10047, y0_1[110]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U528 ( .a ({new_AGEMA_signal_9728, mcs_out[239]}), .b ({w0_s1[111], w0_s0[111]}), .c ({new_AGEMA_signal_9839, y0_1[111]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U529 ( .a ({new_AGEMA_signal_10666, mcs_out[240]}), .b ({w0_s1[112], w0_s0[112]}), .c ({new_AGEMA_signal_10767, y0_1[112]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U530 ( .a ({new_AGEMA_signal_10896, mcs_out[241]}), .b ({w0_s1[113], w0_s0[113]}), .c ({new_AGEMA_signal_10960, y0_1[113]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U531 ( .a ({new_AGEMA_signal_10145, mcs_out[242]}), .b ({w0_s1[114], w0_s0[114]}), .c ({new_AGEMA_signal_10279, y0_1[114]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U532 ( .a ({new_AGEMA_signal_10895, mcs_out[243]}), .b ({w0_s1[115], w0_s0[115]}), .c ({new_AGEMA_signal_10961, y0_1[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U533 ( .a ({new_AGEMA_signal_10364, mcs_out[244]}), .b ({w0_s1[116], w0_s0[116]}), .c ({new_AGEMA_signal_10516, y0_1[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U534 ( .a ({new_AGEMA_signal_10647, mcs_out[245]}), .b ({w0_s1[117], w0_s0[117]}), .c ({new_AGEMA_signal_10768, y0_1[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U535 ( .a ({new_AGEMA_signal_10887, mcs_out[246]}), .b ({w0_s1[118], w0_s0[118]}), .c ({new_AGEMA_signal_10962, y0_1[118]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U536 ( .a ({new_AGEMA_signal_10886, mcs_out[247]}), .b ({w0_s1[119], w0_s0[119]}), .c ({new_AGEMA_signal_10963, y0_1[119]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U537 ( .a ({new_AGEMA_signal_10917, mcs_out[139]}), .b ({w0_s1[11], w0_s0[11]}), .c ({new_AGEMA_signal_10964, y0_1[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U538 ( .a ({new_AGEMA_signal_10878, mcs_out[248]}), .b ({w0_s1[120], w0_s0[120]}), .c ({new_AGEMA_signal_10965, y0_1[120]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U539 ( .a ({new_AGEMA_signal_10097, mcs_out[249]}), .b ({w0_s1[121], w0_s0[121]}), .c ({new_AGEMA_signal_10280, y0_1[121]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U540 ( .a ({new_AGEMA_signal_10339, mcs_out[250]}), .b ({w0_s1[122], w0_s0[122]}), .c ({new_AGEMA_signal_10517, y0_1[122]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U541 ( .a ({new_AGEMA_signal_10629, mcs_out[251]}), .b ({w0_s1[123], w0_s0[123]}), .c ({new_AGEMA_signal_10769, y0_1[123]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U542 ( .a ({new_AGEMA_signal_9622, mcs_out[252]}), .b ({w0_s1[124], w0_s0[124]}), .c ({new_AGEMA_signal_9840, y0_1[124]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U543 ( .a ({new_AGEMA_signal_9862, mcs_out[253]}), .b ({w0_s1[125], w0_s0[125]}), .c ({new_AGEMA_signal_10048, y0_1[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U544 ( .a ({new_AGEMA_signal_9861, mcs_out[254]}), .b ({w0_s1[126], w0_s0[126]}), .c ({new_AGEMA_signal_10049, y0_1[126]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U545 ( .a ({new_AGEMA_signal_9619, mcs_out[255]}), .b ({w0_s1[127], w0_s0[127]}), .c ({new_AGEMA_signal_9841, y0_1[127]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U546 ( .a ({new_AGEMA_signal_10910, mcs_out[140]}), .b ({w0_s1[12], w0_s0[12]}), .c ({new_AGEMA_signal_10966, y0_1[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U547 ( .a ({new_AGEMA_signal_10173, mcs_out[141]}), .b ({w0_s1[13], w0_s0[13]}), .c ({new_AGEMA_signal_10281, y0_1[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U548 ( .a ({new_AGEMA_signal_9732, mcs_out[142]}), .b ({w0_s1[14], w0_s0[14]}), .c ({new_AGEMA_signal_9842, y0_1[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U549 ( .a ({new_AGEMA_signal_10689, mcs_out[143]}), .b ({w0_s1[15], w0_s0[15]}), .c ({new_AGEMA_signal_10770, y0_1[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U550 ( .a ({new_AGEMA_signal_10899, mcs_out[144]}), .b ({w0_s1[16], w0_s0[16]}), .c ({new_AGEMA_signal_10967, y0_1[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U551 ( .a ({new_AGEMA_signal_10394, mcs_out[145]}), .b ({w0_s1[17], w0_s0[17]}), .c ({new_AGEMA_signal_10518, y0_1[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U552 ( .a ({new_AGEMA_signal_10898, mcs_out[146]}), .b ({w0_s1[18], w0_s0[18]}), .c ({new_AGEMA_signal_10968, y0_1[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U553 ( .a ({new_AGEMA_signal_10147, mcs_out[147]}), .b ({w0_s1[19], w0_s0[19]}), .c ({new_AGEMA_signal_10282, y0_1[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U554 ( .a ({new_AGEMA_signal_10489, mcs_out[129]}), .b ({w0_s1[1], w0_s0[1]}), .c ({new_AGEMA_signal_10519, y0_1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U555 ( .a ({new_AGEMA_signal_10653, mcs_out[148]}), .b ({w0_s1[20], w0_s0[20]}), .c ({new_AGEMA_signal_10771, y0_1[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U556 ( .a ({new_AGEMA_signal_10889, mcs_out[149]}), .b ({w0_s1[21], w0_s0[21]}), .c ({new_AGEMA_signal_10969, y0_1[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U557 ( .a ({new_AGEMA_signal_10888, mcs_out[150]}), .b ({w0_s1[22], w0_s0[22]}), .c ({new_AGEMA_signal_10970, y0_1[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U558 ( .a ({new_AGEMA_signal_10650, mcs_out[151]}), .b ({w0_s1[23], w0_s0[23]}), .c ({new_AGEMA_signal_10772, y0_1[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U559 ( .a ({new_AGEMA_signal_11048, mcs_out[152]}), .b ({w0_s1[24], w0_s0[24]}), .c ({new_AGEMA_signal_11084, y0_1[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U560 ( .a ({new_AGEMA_signal_10102, mcs_out[153]}), .b ({w0_s1[25], w0_s0[25]}), .c ({new_AGEMA_signal_10283, y0_1[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U561 ( .a ({new_AGEMA_signal_10635, mcs_out[154]}), .b ({w0_s1[26], w0_s0[26]}), .c ({new_AGEMA_signal_10773, y0_1[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U562 ( .a ({new_AGEMA_signal_10880, mcs_out[155]}), .b ({w0_s1[27], w0_s0[27]}), .c ({new_AGEMA_signal_10971, y0_1[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U563 ( .a ({new_AGEMA_signal_10873, mcs_out[156]}), .b ({w0_s1[28], w0_s0[28]}), .c ({new_AGEMA_signal_10972, y0_1[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U564 ( .a ({new_AGEMA_signal_10074, mcs_out[157]}), .b ({w0_s1[29], w0_s0[29]}), .c ({new_AGEMA_signal_10284, y0_1[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U565 ( .a ({new_AGEMA_signal_10935, mcs_out[130]}), .b ({w0_s1[2], w0_s0[2]}), .c ({new_AGEMA_signal_10973, y0_1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U566 ( .a ({new_AGEMA_signal_9623, mcs_out[158]}), .b ({w0_s1[30], w0_s0[30]}), .c ({new_AGEMA_signal_9843, y0_1[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U567 ( .a ({new_AGEMA_signal_10620, mcs_out[159]}), .b ({w0_s1[31], w0_s0[31]}), .c ({new_AGEMA_signal_10774, y0_1[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U568 ( .a ({new_AGEMA_signal_9812, mcs_out[160]}), .b ({w0_s1[32], w0_s0[32]}), .c ({new_AGEMA_signal_9844, y0_1[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U569 ( .a ({new_AGEMA_signal_10025, mcs_out[161]}), .b ({w0_s1[33], w0_s0[33]}), .c ({new_AGEMA_signal_10050, y0_1[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U570 ( .a ({new_AGEMA_signal_10024, mcs_out[162]}), .b ({w0_s1[34], w0_s0[34]}), .c ({new_AGEMA_signal_10051, y0_1[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U571 ( .a ({new_AGEMA_signal_10023, mcs_out[163]}), .b ({w0_s1[35], w0_s0[35]}), .c ({new_AGEMA_signal_10052, y0_1[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U572 ( .a ({new_AGEMA_signal_10463, mcs_out[164]}), .b ({w0_s1[36], w0_s0[36]}), .c ({new_AGEMA_signal_10520, y0_1[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U573 ( .a ({new_AGEMA_signal_9781, mcs_out[165]}), .b ({w0_s1[37], w0_s0[37]}), .c ({new_AGEMA_signal_9845, y0_1[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U574 ( .a ({new_AGEMA_signal_9286, mcs_out[166]}), .b ({w0_s1[38], w0_s0[38]}), .c ({new_AGEMA_signal_9354, y0_1[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U575 ( .a ({new_AGEMA_signal_10223, mcs_out[167]}), .b ({w0_s1[39], w0_s0[39]}), .c ({new_AGEMA_signal_10285, y0_1[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U576 ( .a ({new_AGEMA_signal_10246, mcs_out[131]}), .b ({w0_s1[3], w0_s0[3]}), .c ({new_AGEMA_signal_10286, y0_1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U577 ( .a ({new_AGEMA_signal_10701, mcs_out[168]}), .b ({w0_s1[40], w0_s0[40]}), .c ({new_AGEMA_signal_10775, y0_1[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U578 ( .a ({new_AGEMA_signal_10439, mcs_out[169]}), .b ({w0_s1[41], w0_s0[41]}), .c ({new_AGEMA_signal_10521, y0_1[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U579 ( .a ({new_AGEMA_signal_10438, mcs_out[170]}), .b ({w0_s1[42], w0_s0[42]}), .c ({new_AGEMA_signal_10522, y0_1[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U580 ( .a ({new_AGEMA_signal_10437, mcs_out[171]}), .b ({w0_s1[43], w0_s0[43]}), .c ({new_AGEMA_signal_10523, y0_1[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U581 ( .a ({new_AGEMA_signal_10909, mcs_out[172]}), .b ({w0_s1[44], w0_s0[44]}), .c ({new_AGEMA_signal_10974, y0_1[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U582 ( .a ({new_AGEMA_signal_10172, mcs_out[173]}), .b ({w0_s1[45], w0_s0[45]}), .c ({new_AGEMA_signal_10287, y0_1[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U583 ( .a ({new_AGEMA_signal_10171, mcs_out[174]}), .b ({w0_s1[46], w0_s0[46]}), .c ({new_AGEMA_signal_10288, y0_1[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U584 ( .a ({new_AGEMA_signal_10686, mcs_out[175]}), .b ({w0_s1[47], w0_s0[47]}), .c ({new_AGEMA_signal_10776, y0_1[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U585 ( .a ({new_AGEMA_signal_9703, mcs_out[176]}), .b ({w0_s1[48], w0_s0[48]}), .c ({new_AGEMA_signal_9846, y0_1[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U586 ( .a ({new_AGEMA_signal_9932, mcs_out[177]}), .b ({w0_s1[49], w0_s0[49]}), .c ({new_AGEMA_signal_10053, y0_1[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U587 ( .a ({new_AGEMA_signal_10722, mcs_out[132]}), .b ({w0_s1[4], w0_s0[4]}), .c ({new_AGEMA_signal_10777, y0_1[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U588 ( .a ({new_AGEMA_signal_9931, mcs_out[178]}), .b ({w0_s1[50], w0_s0[50]}), .c ({new_AGEMA_signal_10054, y0_1[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U589 ( .a ({new_AGEMA_signal_9930, mcs_out[179]}), .b ({w0_s1[51], w0_s0[51]}), .c ({new_AGEMA_signal_10055, y0_1[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U590 ( .a ({new_AGEMA_signal_10368, mcs_out[180]}), .b ({w0_s1[52], w0_s0[52]}), .c ({new_AGEMA_signal_10524, y0_1[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U591 ( .a ({new_AGEMA_signal_9672, mcs_out[181]}), .b ({w0_s1[53], w0_s0[53]}), .c ({new_AGEMA_signal_9847, y0_1[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U592 ( .a ({new_AGEMA_signal_9139, mcs_out[182]}), .b ({w0_s1[54], w0_s0[54]}), .c ({new_AGEMA_signal_9355, y0_1[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U593 ( .a ({new_AGEMA_signal_10124, mcs_out[183]}), .b ({w0_s1[55], w0_s0[55]}), .c ({new_AGEMA_signal_10289, y0_1[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U594 ( .a ({new_AGEMA_signal_10632, mcs_out[184]}), .b ({w0_s1[56], w0_s0[56]}), .c ({new_AGEMA_signal_10778, y0_1[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U595 ( .a ({new_AGEMA_signal_10344, mcs_out[185]}), .b ({w0_s1[57], w0_s0[57]}), .c ({new_AGEMA_signal_10525, y0_1[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U596 ( .a ({new_AGEMA_signal_10343, mcs_out[186]}), .b ({w0_s1[58], w0_s0[58]}), .c ({new_AGEMA_signal_10526, y0_1[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U597 ( .a ({new_AGEMA_signal_10342, mcs_out[187]}), .b ({w0_s1[59], w0_s0[59]}), .c ({new_AGEMA_signal_10527, y0_1[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U598 ( .a ({new_AGEMA_signal_10926, mcs_out[133]}), .b ({w0_s1[5], w0_s0[5]}), .c ({new_AGEMA_signal_10975, y0_1[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U599 ( .a ({new_AGEMA_signal_10872, mcs_out[188]}), .b ({w0_s1[60], w0_s0[60]}), .c ({new_AGEMA_signal_10976, y0_1[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U600 ( .a ({new_AGEMA_signal_10073, mcs_out[189]}), .b ({w0_s1[61], w0_s0[61]}), .c ({new_AGEMA_signal_10290, y0_1[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U601 ( .a ({new_AGEMA_signal_10072, mcs_out[190]}), .b ({w0_s1[62], w0_s0[62]}), .c ({new_AGEMA_signal_10291, y0_1[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U602 ( .a ({new_AGEMA_signal_10617, mcs_out[191]}), .b ({w0_s1[63], w0_s0[63]}), .c ({new_AGEMA_signal_10779, y0_1[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U603 ( .a ({new_AGEMA_signal_10934, mcs_out[192]}), .b ({w0_s1[64], w0_s0[64]}), .c ({new_AGEMA_signal_10977, y0_1[64]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U604 ( .a ({new_AGEMA_signal_10738, mcs_out[193]}), .b ({w0_s1[65], w0_s0[65]}), .c ({new_AGEMA_signal_10780, y0_1[65]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U605 ( .a ({new_AGEMA_signal_10737, mcs_out[194]}), .b ({w0_s1[66], w0_s0[66]}), .c ({new_AGEMA_signal_10781, y0_1[66]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U606 ( .a ({new_AGEMA_signal_10736, mcs_out[195]}), .b ({w0_s1[67], w0_s0[67]}), .c ({new_AGEMA_signal_10782, y0_1[67]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U607 ( .a ({new_AGEMA_signal_10718, mcs_out[196]}), .b ({w0_s1[68], w0_s0[68]}), .c ({new_AGEMA_signal_10783, y0_1[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U608 ( .a ({new_AGEMA_signal_10461, mcs_out[197]}), .b ({w0_s1[69], w0_s0[69]}), .c ({new_AGEMA_signal_10528, y0_1[69]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U609 ( .a ({new_AGEMA_signal_10925, mcs_out[134]}), .b ({w0_s1[6], w0_s0[6]}), .c ({new_AGEMA_signal_10978, y0_1[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U610 ( .a ({new_AGEMA_signal_10221, mcs_out[198]}), .b ({w0_s1[70], w0_s0[70]}), .c ({new_AGEMA_signal_10292, y0_1[70]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U611 ( .a ({new_AGEMA_signal_10717, mcs_out[199]}), .b ({w0_s1[71], w0_s0[71]}), .c ({new_AGEMA_signal_10784, y0_1[71]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U612 ( .a ({new_AGEMA_signal_11100, mcs_out[200]}), .b ({w0_s1[72], w0_s0[72]}), .c ({new_AGEMA_signal_11138, y0_1[72]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U613 ( .a ({new_AGEMA_signal_9976, mcs_out[201]}), .b ({w0_s1[73], w0_s0[73]}), .c ({new_AGEMA_signal_10056, y0_1[73]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U614 ( .a ({new_AGEMA_signal_10436, mcs_out[202]}), .b ({w0_s1[74], w0_s0[74]}), .c ({new_AGEMA_signal_10529, y0_1[74]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U615 ( .a ({new_AGEMA_signal_10916, mcs_out[203]}), .b ({w0_s1[75], w0_s0[75]}), .c ({new_AGEMA_signal_10979, y0_1[75]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U616 ( .a ({new_AGEMA_signal_10908, mcs_out[204]}), .b ({w0_s1[76], w0_s0[76]}), .c ({new_AGEMA_signal_10980, y0_1[76]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U617 ( .a ({new_AGEMA_signal_10907, mcs_out[205]}), .b ({w0_s1[77], w0_s0[77]}), .c ({new_AGEMA_signal_10981, y0_1[77]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U618 ( .a ({new_AGEMA_signal_10906, mcs_out[206]}), .b ({w0_s1[78], w0_s0[78]}), .c ({new_AGEMA_signal_10982, y0_1[78]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U619 ( .a ({new_AGEMA_signal_10905, mcs_out[207]}), .b ({w0_s1[79], w0_s0[79]}), .c ({new_AGEMA_signal_10983, y0_1[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U620 ( .a ({new_AGEMA_signal_10719, mcs_out[135]}), .b ({w0_s1[7], w0_s0[7]}), .c ({new_AGEMA_signal_10785, y0_1[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U621 ( .a ({new_AGEMA_signal_10897, mcs_out[208]}), .b ({w0_s1[80], w0_s0[80]}), .c ({new_AGEMA_signal_10984, y0_1[80]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U622 ( .a ({new_AGEMA_signal_10669, mcs_out[209]}), .b ({w0_s1[81], w0_s0[81]}), .c ({new_AGEMA_signal_10786, y0_1[81]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U623 ( .a ({new_AGEMA_signal_10668, mcs_out[210]}), .b ({w0_s1[82], w0_s0[82]}), .c ({new_AGEMA_signal_10787, y0_1[82]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U624 ( .a ({new_AGEMA_signal_10667, mcs_out[211]}), .b ({w0_s1[83], w0_s0[83]}), .c ({new_AGEMA_signal_10788, y0_1[83]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U625 ( .a ({new_AGEMA_signal_10649, mcs_out[212]}), .b ({w0_s1[84], w0_s0[84]}), .c ({new_AGEMA_signal_10789, y0_1[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U626 ( .a ({new_AGEMA_signal_10366, mcs_out[213]}), .b ({w0_s1[85], w0_s0[85]}), .c ({new_AGEMA_signal_10530, y0_1[85]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U627 ( .a ({new_AGEMA_signal_10122, mcs_out[214]}), .b ({w0_s1[86], w0_s0[86]}), .c ({new_AGEMA_signal_10293, y0_1[86]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U628 ( .a ({new_AGEMA_signal_10648, mcs_out[215]}), .b ({w0_s1[87], w0_s0[87]}), .c ({new_AGEMA_signal_10790, y0_1[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U629 ( .a ({new_AGEMA_signal_11098, mcs_out[216]}), .b ({w0_s1[88], w0_s0[88]}), .c ({new_AGEMA_signal_11139, y0_1[88]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U630 ( .a ({new_AGEMA_signal_9883, mcs_out[217]}), .b ({w0_s1[89], w0_s0[89]}), .c ({new_AGEMA_signal_10057, y0_1[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U631 ( .a ({new_AGEMA_signal_11054, mcs_out[136]}), .b ({w0_s1[8], w0_s0[8]}), .c ({new_AGEMA_signal_11085, y0_1[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U632 ( .a ({new_AGEMA_signal_10341, mcs_out[218]}), .b ({w0_s1[90], w0_s0[90]}), .c ({new_AGEMA_signal_10531, y0_1[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U633 ( .a ({new_AGEMA_signal_10879, mcs_out[219]}), .b ({w0_s1[91], w0_s0[91]}), .c ({new_AGEMA_signal_10985, y0_1[91]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U634 ( .a ({new_AGEMA_signal_10871, mcs_out[220]}), .b ({w0_s1[92], w0_s0[92]}), .c ({new_AGEMA_signal_10986, y0_1[92]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U635 ( .a ({new_AGEMA_signal_10870, mcs_out[221]}), .b ({w0_s1[93], w0_s0[93]}), .c ({new_AGEMA_signal_10987, y0_1[93]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U636 ( .a ({new_AGEMA_signal_10869, mcs_out[222]}), .b ({w0_s1[94], w0_s0[94]}), .c ({new_AGEMA_signal_10988, y0_1[94]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U637 ( .a ({new_AGEMA_signal_10868, mcs_out[223]}), .b ({w0_s1[95], w0_s0[95]}), .c ({new_AGEMA_signal_10989, y0_1[95]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U638 ( .a ({new_AGEMA_signal_10735, mcs_out[224]}), .b ({w0_s1[96], w0_s0[96]}), .c ({new_AGEMA_signal_10791, y0_1[96]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U639 ( .a ({new_AGEMA_signal_10933, mcs_out[225]}), .b ({w0_s1[97], w0_s0[97]}), .c ({new_AGEMA_signal_10990, y0_1[97]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U640 ( .a ({new_AGEMA_signal_10244, mcs_out[226]}), .b ({w0_s1[98], w0_s0[98]}), .c ({new_AGEMA_signal_10294, y0_1[98]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U641 ( .a ({new_AGEMA_signal_10932, mcs_out[227]}), .b ({w0_s1[99], w0_s0[99]}), .c ({new_AGEMA_signal_10991, y0_1[99]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U642 ( .a ({new_AGEMA_signal_10201, mcs_out[137]}), .b ({w0_s1[9], w0_s0[9]}), .c ({new_AGEMA_signal_10295, y0_1[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U643 ( .a ({temp_s1[0], temp_s0[0]}), .b ({temp_next_s1[0], temp_next_s0[0]}), .c ({y1_s1[0], y1_s0[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U644 ( .a ({temp_s1[100], temp_s0[100]}), .b ({temp_next_s1[100], temp_next_s0[100]}), .c ({y1_s1[100], y1_s0[100]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U645 ( .a ({temp_s1[101], temp_s0[101]}), .b ({temp_next_s1[101], temp_next_s0[101]}), .c ({y1_s1[101], y1_s0[101]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U646 ( .a ({temp_s1[102], temp_s0[102]}), .b ({temp_next_s1[102], temp_next_s0[102]}), .c ({y1_s1[102], y1_s0[102]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U647 ( .a ({temp_s1[103], temp_s0[103]}), .b ({temp_next_s1[103], temp_next_s0[103]}), .c ({y1_s1[103], y1_s0[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U648 ( .a ({temp_s1[104], temp_s0[104]}), .b ({temp_next_s1[104], temp_next_s0[104]}), .c ({y1_s1[104], y1_s0[104]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U649 ( .a ({temp_s1[105], temp_s0[105]}), .b ({temp_next_s1[105], temp_next_s0[105]}), .c ({y1_s1[105], y1_s0[105]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U650 ( .a ({temp_s1[106], temp_s0[106]}), .b ({temp_next_s1[106], temp_next_s0[106]}), .c ({y1_s1[106], y1_s0[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U651 ( .a ({temp_s1[107], temp_s0[107]}), .b ({temp_next_s1[107], temp_next_s0[107]}), .c ({y1_s1[107], y1_s0[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U652 ( .a ({temp_s1[108], temp_s0[108]}), .b ({temp_next_s1[108], temp_next_s0[108]}), .c ({y1_s1[108], y1_s0[108]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U653 ( .a ({temp_s1[109], temp_s0[109]}), .b ({temp_next_s1[109], temp_next_s0[109]}), .c ({y1_s1[109], y1_s0[109]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U654 ( .a ({temp_s1[10], temp_s0[10]}), .b ({temp_next_s1[10], temp_next_s0[10]}), .c ({y1_s1[10], y1_s0[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U655 ( .a ({temp_s1[110], temp_s0[110]}), .b ({temp_next_s1[110], temp_next_s0[110]}), .c ({y1_s1[110], y1_s0[110]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U656 ( .a ({temp_s1[111], temp_s0[111]}), .b ({temp_next_s1[111], temp_next_s0[111]}), .c ({y1_s1[111], y1_s0[111]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U657 ( .a ({temp_s1[112], temp_s0[112]}), .b ({temp_next_s1[112], temp_next_s0[112]}), .c ({y1_s1[112], y1_s0[112]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U658 ( .a ({temp_s1[113], temp_s0[113]}), .b ({temp_next_s1[113], temp_next_s0[113]}), .c ({y1_s1[113], y1_s0[113]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U659 ( .a ({temp_s1[114], temp_s0[114]}), .b ({temp_next_s1[114], temp_next_s0[114]}), .c ({y1_s1[114], y1_s0[114]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U660 ( .a ({temp_s1[115], temp_s0[115]}), .b ({temp_next_s1[115], temp_next_s0[115]}), .c ({y1_s1[115], y1_s0[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U661 ( .a ({temp_s1[116], temp_s0[116]}), .b ({temp_next_s1[116], temp_next_s0[116]}), .c ({y1_s1[116], y1_s0[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U662 ( .a ({temp_s1[117], temp_s0[117]}), .b ({temp_next_s1[117], temp_next_s0[117]}), .c ({y1_s1[117], y1_s0[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U663 ( .a ({temp_s1[118], temp_s0[118]}), .b ({temp_next_s1[118], temp_next_s0[118]}), .c ({y1_s1[118], y1_s0[118]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U664 ( .a ({temp_s1[119], temp_s0[119]}), .b ({temp_next_s1[119], temp_next_s0[119]}), .c ({y1_s1[119], y1_s0[119]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U665 ( .a ({temp_s1[11], temp_s0[11]}), .b ({temp_next_s1[11], temp_next_s0[11]}), .c ({y1_s1[11], y1_s0[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U666 ( .a ({temp_s1[120], temp_s0[120]}), .b ({temp_next_s1[120], temp_next_s0[120]}), .c ({y1_s1[120], y1_s0[120]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U667 ( .a ({temp_s1[121], temp_s0[121]}), .b ({temp_next_s1[121], temp_next_s0[121]}), .c ({y1_s1[121], y1_s0[121]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U668 ( .a ({temp_s1[122], temp_s0[122]}), .b ({temp_next_s1[122], temp_next_s0[122]}), .c ({y1_s1[122], y1_s0[122]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U669 ( .a ({temp_s1[123], temp_s0[123]}), .b ({temp_next_s1[123], temp_next_s0[123]}), .c ({y1_s1[123], y1_s0[123]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U670 ( .a ({temp_s1[124], temp_s0[124]}), .b ({temp_next_s1[124], temp_next_s0[124]}), .c ({y1_s1[124], y1_s0[124]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U671 ( .a ({temp_s1[125], temp_s0[125]}), .b ({temp_next_s1[125], temp_next_s0[125]}), .c ({y1_s1[125], y1_s0[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U672 ( .a ({temp_s1[126], temp_s0[126]}), .b ({temp_next_s1[126], temp_next_s0[126]}), .c ({y1_s1[126], y1_s0[126]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U673 ( .a ({temp_s1[127], temp_s0[127]}), .b ({temp_next_s1[127], temp_next_s0[127]}), .c ({y1_s1[127], y1_s0[127]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U674 ( .a ({temp_s1[12], temp_s0[12]}), .b ({temp_next_s1[12], temp_next_s0[12]}), .c ({y1_s1[12], y1_s0[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U675 ( .a ({temp_s1[13], temp_s0[13]}), .b ({temp_next_s1[13], temp_next_s0[13]}), .c ({y1_s1[13], y1_s0[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U676 ( .a ({temp_s1[14], temp_s0[14]}), .b ({temp_next_s1[14], temp_next_s0[14]}), .c ({y1_s1[14], y1_s0[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U677 ( .a ({temp_s1[15], temp_s0[15]}), .b ({temp_next_s1[15], temp_next_s0[15]}), .c ({y1_s1[15], y1_s0[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U678 ( .a ({temp_s1[16], temp_s0[16]}), .b ({temp_next_s1[16], temp_next_s0[16]}), .c ({y1_s1[16], y1_s0[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U679 ( .a ({temp_s1[17], temp_s0[17]}), .b ({temp_next_s1[17], temp_next_s0[17]}), .c ({y1_s1[17], y1_s0[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U680 ( .a ({temp_s1[18], temp_s0[18]}), .b ({temp_next_s1[18], temp_next_s0[18]}), .c ({y1_s1[18], y1_s0[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U681 ( .a ({temp_s1[19], temp_s0[19]}), .b ({temp_next_s1[19], temp_next_s0[19]}), .c ({y1_s1[19], y1_s0[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U682 ( .a ({temp_s1[1], temp_s0[1]}), .b ({temp_next_s1[1], temp_next_s0[1]}), .c ({y1_s1[1], y1_s0[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U683 ( .a ({temp_s1[20], temp_s0[20]}), .b ({temp_next_s1[20], temp_next_s0[20]}), .c ({y1_s1[20], y1_s0[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U684 ( .a ({temp_s1[21], temp_s0[21]}), .b ({temp_next_s1[21], temp_next_s0[21]}), .c ({y1_s1[21], y1_s0[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U685 ( .a ({temp_s1[22], temp_s0[22]}), .b ({temp_next_s1[22], temp_next_s0[22]}), .c ({y1_s1[22], y1_s0[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U686 ( .a ({temp_s1[23], temp_s0[23]}), .b ({temp_next_s1[23], temp_next_s0[23]}), .c ({y1_s1[23], y1_s0[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U687 ( .a ({temp_s1[24], temp_s0[24]}), .b ({temp_next_s1[24], temp_next_s0[24]}), .c ({y1_s1[24], y1_s0[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U688 ( .a ({temp_s1[25], temp_s0[25]}), .b ({temp_next_s1[25], temp_next_s0[25]}), .c ({y1_s1[25], y1_s0[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U689 ( .a ({temp_s1[26], temp_s0[26]}), .b ({temp_next_s1[26], temp_next_s0[26]}), .c ({y1_s1[26], y1_s0[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U690 ( .a ({temp_s1[27], temp_s0[27]}), .b ({temp_next_s1[27], temp_next_s0[27]}), .c ({y1_s1[27], y1_s0[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U691 ( .a ({temp_s1[28], temp_s0[28]}), .b ({temp_next_s1[28], temp_next_s0[28]}), .c ({y1_s1[28], y1_s0[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U692 ( .a ({temp_s1[29], temp_s0[29]}), .b ({temp_next_s1[29], temp_next_s0[29]}), .c ({y1_s1[29], y1_s0[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U693 ( .a ({temp_s1[2], temp_s0[2]}), .b ({temp_next_s1[2], temp_next_s0[2]}), .c ({y1_s1[2], y1_s0[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U694 ( .a ({temp_s1[30], temp_s0[30]}), .b ({temp_next_s1[30], temp_next_s0[30]}), .c ({y1_s1[30], y1_s0[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U695 ( .a ({temp_s1[31], temp_s0[31]}), .b ({temp_next_s1[31], temp_next_s0[31]}), .c ({y1_s1[31], y1_s0[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U696 ( .a ({temp_s1[32], temp_s0[32]}), .b ({temp_next_s1[32], temp_next_s0[32]}), .c ({y1_s1[32], y1_s0[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U697 ( .a ({temp_s1[33], temp_s0[33]}), .b ({temp_next_s1[33], temp_next_s0[33]}), .c ({y1_s1[33], y1_s0[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U698 ( .a ({temp_s1[34], temp_s0[34]}), .b ({temp_next_s1[34], temp_next_s0[34]}), .c ({y1_s1[34], y1_s0[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U699 ( .a ({temp_s1[35], temp_s0[35]}), .b ({temp_next_s1[35], temp_next_s0[35]}), .c ({y1_s1[35], y1_s0[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U700 ( .a ({temp_s1[36], temp_s0[36]}), .b ({temp_next_s1[36], temp_next_s0[36]}), .c ({y1_s1[36], y1_s0[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U701 ( .a ({temp_s1[37], temp_s0[37]}), .b ({temp_next_s1[37], temp_next_s0[37]}), .c ({y1_s1[37], y1_s0[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U702 ( .a ({temp_s1[38], temp_s0[38]}), .b ({temp_next_s1[38], temp_next_s0[38]}), .c ({y1_s1[38], y1_s0[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U703 ( .a ({temp_s1[39], temp_s0[39]}), .b ({temp_next_s1[39], temp_next_s0[39]}), .c ({y1_s1[39], y1_s0[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U704 ( .a ({temp_s1[3], temp_s0[3]}), .b ({temp_next_s1[3], temp_next_s0[3]}), .c ({y1_s1[3], y1_s0[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U705 ( .a ({temp_s1[40], temp_s0[40]}), .b ({temp_next_s1[40], temp_next_s0[40]}), .c ({y1_s1[40], y1_s0[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U706 ( .a ({temp_s1[41], temp_s0[41]}), .b ({temp_next_s1[41], temp_next_s0[41]}), .c ({y1_s1[41], y1_s0[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U707 ( .a ({temp_s1[42], temp_s0[42]}), .b ({temp_next_s1[42], temp_next_s0[42]}), .c ({y1_s1[42], y1_s0[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U708 ( .a ({temp_s1[43], temp_s0[43]}), .b ({temp_next_s1[43], temp_next_s0[43]}), .c ({y1_s1[43], y1_s0[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U709 ( .a ({temp_s1[44], temp_s0[44]}), .b ({temp_next_s1[44], temp_next_s0[44]}), .c ({y1_s1[44], y1_s0[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U710 ( .a ({temp_s1[45], temp_s0[45]}), .b ({temp_next_s1[45], temp_next_s0[45]}), .c ({y1_s1[45], y1_s0[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U711 ( .a ({temp_s1[46], temp_s0[46]}), .b ({temp_next_s1[46], temp_next_s0[46]}), .c ({y1_s1[46], y1_s0[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U712 ( .a ({temp_s1[47], temp_s0[47]}), .b ({temp_next_s1[47], temp_next_s0[47]}), .c ({y1_s1[47], y1_s0[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U713 ( .a ({temp_s1[48], temp_s0[48]}), .b ({temp_next_s1[48], temp_next_s0[48]}), .c ({y1_s1[48], y1_s0[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U714 ( .a ({temp_s1[49], temp_s0[49]}), .b ({temp_next_s1[49], temp_next_s0[49]}), .c ({y1_s1[49], y1_s0[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U715 ( .a ({temp_s1[4], temp_s0[4]}), .b ({temp_next_s1[4], temp_next_s0[4]}), .c ({y1_s1[4], y1_s0[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U716 ( .a ({temp_s1[50], temp_s0[50]}), .b ({temp_next_s1[50], temp_next_s0[50]}), .c ({y1_s1[50], y1_s0[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U717 ( .a ({temp_s1[51], temp_s0[51]}), .b ({temp_next_s1[51], temp_next_s0[51]}), .c ({y1_s1[51], y1_s0[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U718 ( .a ({temp_s1[52], temp_s0[52]}), .b ({temp_next_s1[52], temp_next_s0[52]}), .c ({y1_s1[52], y1_s0[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U719 ( .a ({temp_s1[53], temp_s0[53]}), .b ({temp_next_s1[53], temp_next_s0[53]}), .c ({y1_s1[53], y1_s0[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U720 ( .a ({temp_s1[54], temp_s0[54]}), .b ({temp_next_s1[54], temp_next_s0[54]}), .c ({y1_s1[54], y1_s0[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U721 ( .a ({temp_s1[55], temp_s0[55]}), .b ({temp_next_s1[55], temp_next_s0[55]}), .c ({y1_s1[55], y1_s0[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U722 ( .a ({temp_s1[56], temp_s0[56]}), .b ({temp_next_s1[56], temp_next_s0[56]}), .c ({y1_s1[56], y1_s0[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U723 ( .a ({temp_s1[57], temp_s0[57]}), .b ({temp_next_s1[57], temp_next_s0[57]}), .c ({y1_s1[57], y1_s0[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U724 ( .a ({temp_s1[58], temp_s0[58]}), .b ({temp_next_s1[58], temp_next_s0[58]}), .c ({y1_s1[58], y1_s0[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U725 ( .a ({temp_s1[59], temp_s0[59]}), .b ({temp_next_s1[59], temp_next_s0[59]}), .c ({y1_s1[59], y1_s0[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U726 ( .a ({temp_s1[5], temp_s0[5]}), .b ({temp_next_s1[5], temp_next_s0[5]}), .c ({y1_s1[5], y1_s0[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U727 ( .a ({temp_s1[60], temp_s0[60]}), .b ({temp_next_s1[60], temp_next_s0[60]}), .c ({y1_s1[60], y1_s0[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U728 ( .a ({temp_s1[61], temp_s0[61]}), .b ({temp_next_s1[61], temp_next_s0[61]}), .c ({y1_s1[61], y1_s0[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U729 ( .a ({temp_s1[62], temp_s0[62]}), .b ({temp_next_s1[62], temp_next_s0[62]}), .c ({y1_s1[62], y1_s0[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U730 ( .a ({temp_s1[63], temp_s0[63]}), .b ({temp_next_s1[63], temp_next_s0[63]}), .c ({y1_s1[63], y1_s0[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U731 ( .a ({temp_s1[64], temp_s0[64]}), .b ({temp_next_s1[64], temp_next_s0[64]}), .c ({y1_s1[64], y1_s0[64]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U732 ( .a ({temp_s1[65], temp_s0[65]}), .b ({temp_next_s1[65], temp_next_s0[65]}), .c ({y1_s1[65], y1_s0[65]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U733 ( .a ({temp_s1[66], temp_s0[66]}), .b ({temp_next_s1[66], temp_next_s0[66]}), .c ({y1_s1[66], y1_s0[66]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U734 ( .a ({temp_s1[67], temp_s0[67]}), .b ({temp_next_s1[67], temp_next_s0[67]}), .c ({y1_s1[67], y1_s0[67]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U735 ( .a ({temp_s1[68], temp_s0[68]}), .b ({temp_next_s1[68], temp_next_s0[68]}), .c ({y1_s1[68], y1_s0[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U736 ( .a ({temp_s1[69], temp_s0[69]}), .b ({temp_next_s1[69], temp_next_s0[69]}), .c ({y1_s1[69], y1_s0[69]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U737 ( .a ({temp_s1[6], temp_s0[6]}), .b ({temp_next_s1[6], temp_next_s0[6]}), .c ({y1_s1[6], y1_s0[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U738 ( .a ({temp_s1[70], temp_s0[70]}), .b ({temp_next_s1[70], temp_next_s0[70]}), .c ({y1_s1[70], y1_s0[70]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U739 ( .a ({temp_s1[71], temp_s0[71]}), .b ({temp_next_s1[71], temp_next_s0[71]}), .c ({y1_s1[71], y1_s0[71]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U740 ( .a ({temp_s1[72], temp_s0[72]}), .b ({temp_next_s1[72], temp_next_s0[72]}), .c ({y1_s1[72], y1_s0[72]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U741 ( .a ({temp_s1[73], temp_s0[73]}), .b ({temp_next_s1[73], temp_next_s0[73]}), .c ({y1_s1[73], y1_s0[73]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U742 ( .a ({temp_s1[74], temp_s0[74]}), .b ({temp_next_s1[74], temp_next_s0[74]}), .c ({y1_s1[74], y1_s0[74]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U743 ( .a ({temp_s1[75], temp_s0[75]}), .b ({temp_next_s1[75], temp_next_s0[75]}), .c ({y1_s1[75], y1_s0[75]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U744 ( .a ({temp_s1[76], temp_s0[76]}), .b ({temp_next_s1[76], temp_next_s0[76]}), .c ({y1_s1[76], y1_s0[76]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U745 ( .a ({temp_s1[77], temp_s0[77]}), .b ({temp_next_s1[77], temp_next_s0[77]}), .c ({y1_s1[77], y1_s0[77]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U746 ( .a ({temp_s1[78], temp_s0[78]}), .b ({temp_next_s1[78], temp_next_s0[78]}), .c ({y1_s1[78], y1_s0[78]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U747 ( .a ({temp_s1[79], temp_s0[79]}), .b ({temp_next_s1[79], temp_next_s0[79]}), .c ({y1_s1[79], y1_s0[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U748 ( .a ({temp_s1[7], temp_s0[7]}), .b ({temp_next_s1[7], temp_next_s0[7]}), .c ({y1_s1[7], y1_s0[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U749 ( .a ({temp_s1[80], temp_s0[80]}), .b ({temp_next_s1[80], temp_next_s0[80]}), .c ({y1_s1[80], y1_s0[80]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U750 ( .a ({temp_s1[81], temp_s0[81]}), .b ({temp_next_s1[81], temp_next_s0[81]}), .c ({y1_s1[81], y1_s0[81]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U751 ( .a ({temp_s1[82], temp_s0[82]}), .b ({temp_next_s1[82], temp_next_s0[82]}), .c ({y1_s1[82], y1_s0[82]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U752 ( .a ({temp_s1[83], temp_s0[83]}), .b ({temp_next_s1[83], temp_next_s0[83]}), .c ({y1_s1[83], y1_s0[83]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U753 ( .a ({temp_s1[84], temp_s0[84]}), .b ({temp_next_s1[84], temp_next_s0[84]}), .c ({y1_s1[84], y1_s0[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U754 ( .a ({temp_s1[85], temp_s0[85]}), .b ({temp_next_s1[85], temp_next_s0[85]}), .c ({y1_s1[85], y1_s0[85]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U755 ( .a ({temp_s1[86], temp_s0[86]}), .b ({temp_next_s1[86], temp_next_s0[86]}), .c ({y1_s1[86], y1_s0[86]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U756 ( .a ({temp_s1[87], temp_s0[87]}), .b ({temp_next_s1[87], temp_next_s0[87]}), .c ({y1_s1[87], y1_s0[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U757 ( .a ({temp_s1[88], temp_s0[88]}), .b ({temp_next_s1[88], temp_next_s0[88]}), .c ({y1_s1[88], y1_s0[88]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U758 ( .a ({temp_s1[89], temp_s0[89]}), .b ({temp_next_s1[89], temp_next_s0[89]}), .c ({y1_s1[89], y1_s0[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U759 ( .a ({temp_s1[8], temp_s0[8]}), .b ({temp_next_s1[8], temp_next_s0[8]}), .c ({y1_s1[8], y1_s0[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U760 ( .a ({temp_s1[90], temp_s0[90]}), .b ({temp_next_s1[90], temp_next_s0[90]}), .c ({y1_s1[90], y1_s0[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U761 ( .a ({temp_s1[91], temp_s0[91]}), .b ({temp_next_s1[91], temp_next_s0[91]}), .c ({y1_s1[91], y1_s0[91]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U762 ( .a ({temp_s1[92], temp_s0[92]}), .b ({temp_next_s1[92], temp_next_s0[92]}), .c ({y1_s1[92], y1_s0[92]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U763 ( .a ({temp_s1[93], temp_s0[93]}), .b ({temp_next_s1[93], temp_next_s0[93]}), .c ({y1_s1[93], y1_s0[93]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U764 ( .a ({temp_s1[94], temp_s0[94]}), .b ({temp_next_s1[94], temp_next_s0[94]}), .c ({y1_s1[94], y1_s0[94]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U765 ( .a ({temp_s1[95], temp_s0[95]}), .b ({temp_next_s1[95], temp_next_s0[95]}), .c ({y1_s1[95], y1_s0[95]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U766 ( .a ({temp_s1[96], temp_s0[96]}), .b ({temp_next_s1[96], temp_next_s0[96]}), .c ({y1_s1[96], y1_s0[96]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U767 ( .a ({temp_s1[97], temp_s0[97]}), .b ({temp_next_s1[97], temp_next_s0[97]}), .c ({y1_s1[97], y1_s0[97]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U768 ( .a ({temp_s1[98], temp_s0[98]}), .b ({temp_next_s1[98], temp_next_s0[98]}), .c ({y1_s1[98], y1_s0[98]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U769 ( .a ({temp_s1[99], temp_s0[99]}), .b ({temp_next_s1[99], temp_next_s0[99]}), .c ({y1_s1[99], y1_s0[99]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U770 ( .a ({temp_s1[9], temp_s0[9]}), .b ({temp_next_s1[9], temp_next_s0[9]}), .c ({y1_s1[9], y1_s0[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U96 ( .a ({new_AGEMA_signal_9364, mcs1_mcs_mat1_0_n128}), .b ({new_AGEMA_signal_9860, mcs1_mcs_mat1_0_n127}), .c ({temp_next_s1[93], temp_next_s0[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U95 ( .a ({new_AGEMA_signal_8623, mcs1_mcs_mat1_0_mcs_out[41]}), .b ({new_AGEMA_signal_9636, mcs1_mcs_mat1_0_mcs_out[45]}), .c ({new_AGEMA_signal_9860, mcs1_mcs_mat1_0_n127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U94 ( .a ({new_AGEMA_signal_7248, mcs1_mcs_mat1_0_mcs_out[33]}), .b ({new_AGEMA_signal_9084, mcs1_mcs_mat1_0_mcs_out[37]}), .c ({new_AGEMA_signal_9364, mcs1_mcs_mat1_0_n128}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U93 ( .a ({new_AGEMA_signal_9618, mcs1_mcs_mat1_0_n126}), .b ({new_AGEMA_signal_10864, mcs1_mcs_mat1_0_n125}), .c ({temp_next_s1[92], temp_next_s0[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U92 ( .a ({new_AGEMA_signal_8139, mcs1_mcs_mat1_0_mcs_out[40]}), .b ({new_AGEMA_signal_10625, mcs1_mcs_mat1_0_mcs_out[44]}), .c ({new_AGEMA_signal_10864, mcs1_mcs_mat1_0_n125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U91 ( .a ({new_AGEMA_signal_9391, mcs1_mcs_mat1_0_mcs_out[32]}), .b ({new_AGEMA_signal_8141, mcs1_mcs_mat1_0_mcs_out[36]}), .c ({new_AGEMA_signal_9618, mcs1_mcs_mat1_0_n126}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U90 ( .a ({new_AGEMA_signal_8580, mcs1_mcs_mat1_0_n124}), .b ({new_AGEMA_signal_10608, mcs1_mcs_mat1_0_n123}), .c ({temp_next_s1[63], temp_next_s0[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U89 ( .a ({new_AGEMA_signal_8145, mcs1_mcs_mat1_0_mcs_out[27]}), .b ({new_AGEMA_signal_10330, mcs1_mcs_mat1_0_mcs_out[31]}), .c ({new_AGEMA_signal_10608, mcs1_mcs_mat1_0_n123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U88 ( .a ({new_AGEMA_signal_8151, mcs1_mcs_mat1_0_mcs_out[19]}), .b ({new_AGEMA_signal_8148, mcs1_mcs_mat1_0_mcs_out[23]}), .c ({new_AGEMA_signal_8580, mcs1_mcs_mat1_0_n124}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U87 ( .a ({new_AGEMA_signal_9060, mcs1_mcs_mat1_0_n122}), .b ({new_AGEMA_signal_10312, mcs1_mcs_mat1_0_n121}), .c ({temp_next_s1[62], temp_next_s0[62]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U86 ( .a ({new_AGEMA_signal_8628, mcs1_mcs_mat1_0_mcs_out[26]}), .b ({new_AGEMA_signal_10087, mcs1_mcs_mat1_0_mcs_out[30]}), .c ({new_AGEMA_signal_10312, mcs1_mcs_mat1_0_n121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U85 ( .a ({new_AGEMA_signal_8632, mcs1_mcs_mat1_0_mcs_out[18]}), .b ({new_AGEMA_signal_8630, mcs1_mcs_mat1_0_mcs_out[22]}), .c ({new_AGEMA_signal_9060, mcs1_mcs_mat1_0_n122}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U84 ( .a ({new_AGEMA_signal_9365, mcs1_mcs_mat1_0_n120}), .b ({new_AGEMA_signal_10071, mcs1_mcs_mat1_0_n119}), .c ({temp_next_s1[61], temp_next_s0[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U83 ( .a ({new_AGEMA_signal_9086, mcs1_mcs_mat1_0_mcs_out[25]}), .b ({new_AGEMA_signal_9877, mcs1_mcs_mat1_0_mcs_out[29]}), .c ({new_AGEMA_signal_10071, mcs1_mcs_mat1_0_n119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U82 ( .a ({new_AGEMA_signal_9088, mcs1_mcs_mat1_0_mcs_out[17]}), .b ({new_AGEMA_signal_9087, mcs1_mcs_mat1_0_mcs_out[21]}), .c ({new_AGEMA_signal_9365, mcs1_mcs_mat1_0_n120}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U81 ( .a ({new_AGEMA_signal_8581, mcs1_mcs_mat1_0_n118}), .b ({new_AGEMA_signal_10610, mcs1_mcs_mat1_0_n117}), .c ({temp_next_s1[60], temp_next_s0[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U80 ( .a ({new_AGEMA_signal_8147, mcs1_mcs_mat1_0_mcs_out[24]}), .b ({new_AGEMA_signal_10331, mcs1_mcs_mat1_0_mcs_out[28]}), .c ({new_AGEMA_signal_10610, mcs1_mcs_mat1_0_n117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U79 ( .a ({new_AGEMA_signal_8153, mcs1_mcs_mat1_0_mcs_out[16]}), .b ({new_AGEMA_signal_8150, mcs1_mcs_mat1_0_mcs_out[20]}), .c ({new_AGEMA_signal_8581, mcs1_mcs_mat1_0_n118}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U78 ( .a ({new_AGEMA_signal_10611, mcs1_mcs_mat1_0_n116}), .b ({new_AGEMA_signal_9366, mcs1_mcs_mat1_0_n115}), .c ({temp_next_s1[31], temp_next_s0[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U77 ( .a ({new_AGEMA_signal_8158, mcs1_mcs_mat1_0_mcs_out[3]}), .b ({new_AGEMA_signal_9091, mcs1_mcs_mat1_0_mcs_out[7]}), .c ({new_AGEMA_signal_9366, mcs1_mcs_mat1_0_n115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U76 ( .a ({new_AGEMA_signal_7344, mcs1_mcs_mat1_0_mcs_out[11]}), .b ({new_AGEMA_signal_10332, mcs1_mcs_mat1_0_mcs_out[15]}), .c ({new_AGEMA_signal_10611, mcs1_mcs_mat1_0_n116}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U75 ( .a ({new_AGEMA_signal_9368, mcs1_mcs_mat1_0_n114}), .b ({new_AGEMA_signal_9367, mcs1_mcs_mat1_0_n113}), .c ({new_AGEMA_signal_9619, mcs_out[255]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U74 ( .a ({new_AGEMA_signal_9068, mcs1_mcs_mat1_0_mcs_out[123]}), .b ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_9367, mcs1_mcs_mat1_0_n113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U73 ( .a ({new_AGEMA_signal_8594, mcs1_mcs_mat1_0_mcs_out[115]}), .b ({new_AGEMA_signal_9070, mcs1_mcs_mat1_0_mcs_out[119]}), .c ({new_AGEMA_signal_9368, mcs1_mcs_mat1_0_n114}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U72 ( .a ({new_AGEMA_signal_9369, mcs1_mcs_mat1_0_n112}), .b ({new_AGEMA_signal_9620, mcs1_mcs_mat1_0_n111}), .c ({new_AGEMA_signal_9861, mcs_out[254]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U71 ( .a ({new_AGEMA_signal_7622, mcs1_mcs_mat1_0_mcs_out[122]}), .b ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_9620, mcs1_mcs_mat1_0_n111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U70 ( .a ({new_AGEMA_signal_8106, mcs1_mcs_mat1_0_mcs_out[114]}), .b ({new_AGEMA_signal_9071, mcs1_mcs_mat1_0_mcs_out[118]}), .c ({new_AGEMA_signal_9369, mcs1_mcs_mat1_0_n112}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U69 ( .a ({new_AGEMA_signal_10314, mcs1_mcs_mat1_0_n110}), .b ({new_AGEMA_signal_8582, mcs1_mcs_mat1_0_n109}), .c ({temp_next_s1[30], temp_next_s0[30]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U68 ( .a ({new_AGEMA_signal_8159, mcs1_mcs_mat1_0_mcs_out[2]}), .b ({new_AGEMA_signal_8157, mcs1_mcs_mat1_0_mcs_out[6]}), .c ({new_AGEMA_signal_8582, mcs1_mcs_mat1_0_n109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U67 ( .a ({new_AGEMA_signal_8635, mcs1_mcs_mat1_0_mcs_out[10]}), .b ({new_AGEMA_signal_10089, mcs1_mcs_mat1_0_mcs_out[14]}), .c ({new_AGEMA_signal_10314, mcs1_mcs_mat1_0_n110}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U66 ( .a ({new_AGEMA_signal_9061, mcs1_mcs_mat1_0_n108}), .b ({new_AGEMA_signal_9621, mcs1_mcs_mat1_0_n107}), .c ({new_AGEMA_signal_9862, mcs_out[253]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U65 ( .a ({new_AGEMA_signal_9069, mcs1_mcs_mat1_0_mcs_out[121]}), .b ({new_AGEMA_signal_9380, mcs1_mcs_mat1_0_mcs_out[125]}), .c ({new_AGEMA_signal_9621, mcs1_mcs_mat1_0_n107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U64 ( .a ({new_AGEMA_signal_7627, mcs1_mcs_mat1_0_mcs_out[113]}), .b ({new_AGEMA_signal_8593, mcs1_mcs_mat1_0_mcs_out[117]}), .c ({new_AGEMA_signal_9061, mcs1_mcs_mat1_0_n108}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U63 ( .a ({new_AGEMA_signal_9371, mcs1_mcs_mat1_0_n106}), .b ({new_AGEMA_signal_9370, mcs1_mcs_mat1_0_n105}), .c ({new_AGEMA_signal_9622, mcs_out[252]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U62 ( .a ({new_AGEMA_signal_8590, mcs1_mcs_mat1_0_mcs_out[120]}), .b ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_9370, mcs1_mcs_mat1_0_n105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U61 ( .a ({new_AGEMA_signal_9072, mcs1_mcs_mat1_0_mcs_out[112]}), .b ({new_AGEMA_signal_8105, mcs1_mcs_mat1_0_mcs_out[116]}), .c ({new_AGEMA_signal_9371, mcs1_mcs_mat1_0_n106}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U60 ( .a ({new_AGEMA_signal_9062, mcs1_mcs_mat1_0_n104}), .b ({new_AGEMA_signal_10613, mcs1_mcs_mat1_0_n103}), .c ({new_AGEMA_signal_10868, mcs_out[223]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U59 ( .a ({new_AGEMA_signal_10322, mcs1_mcs_mat1_0_mcs_out[111]}), .b ({new_AGEMA_signal_9074, mcs1_mcs_mat1_0_mcs_out[99]}), .c ({new_AGEMA_signal_10613, mcs1_mcs_mat1_0_n103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U58 ( .a ({new_AGEMA_signal_8601, mcs1_mcs_mat1_0_mcs_out[103]}), .b ({new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[107]}), .c ({new_AGEMA_signal_9062, mcs1_mcs_mat1_0_n104}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U57 ( .a ({new_AGEMA_signal_9063, mcs1_mcs_mat1_0_n102}), .b ({new_AGEMA_signal_10614, mcs1_mcs_mat1_0_n101}), .c ({new_AGEMA_signal_10869, mcs_out[222]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U56 ( .a ({new_AGEMA_signal_10323, mcs1_mcs_mat1_0_mcs_out[110]}), .b ({new_AGEMA_signal_8115, mcs1_mcs_mat1_0_mcs_out[98]}), .c ({new_AGEMA_signal_10614, mcs1_mcs_mat1_0_n101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U55 ( .a ({new_AGEMA_signal_7632, mcs1_mcs_mat1_0_mcs_out[102]}), .b ({new_AGEMA_signal_8598, mcs1_mcs_mat1_0_mcs_out[106]}), .c ({new_AGEMA_signal_9063, mcs1_mcs_mat1_0_n102}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U54 ( .a ({new_AGEMA_signal_9064, mcs1_mcs_mat1_0_n100}), .b ({new_AGEMA_signal_10615, mcs1_mcs_mat1_0_n99}), .c ({new_AGEMA_signal_10870, mcs_out[221]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U53 ( .a ({new_AGEMA_signal_10324, mcs1_mcs_mat1_0_mcs_out[109]}), .b ({new_AGEMA_signal_7323, mcs1_mcs_mat1_0_mcs_out[97]}), .c ({new_AGEMA_signal_10615, mcs1_mcs_mat1_0_n99}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U52 ( .a ({new_AGEMA_signal_8113, mcs1_mcs_mat1_0_mcs_out[101]}), .b ({new_AGEMA_signal_8599, mcs1_mcs_mat1_0_mcs_out[105]}), .c ({new_AGEMA_signal_9064, mcs1_mcs_mat1_0_n100}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U51 ( .a ({new_AGEMA_signal_9372, mcs1_mcs_mat1_0_n98}), .b ({new_AGEMA_signal_10616, mcs1_mcs_mat1_0_n97}), .c ({new_AGEMA_signal_10871, mcs_out[220]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U50 ( .a ({new_AGEMA_signal_10325, mcs1_mcs_mat1_0_mcs_out[108]}), .b ({new_AGEMA_signal_9628, mcs1_mcs_mat1_0_mcs_out[96]}), .c ({new_AGEMA_signal_10616, mcs1_mcs_mat1_0_n97}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U49 ( .a ({new_AGEMA_signal_8602, mcs1_mcs_mat1_0_mcs_out[100]}), .b ({new_AGEMA_signal_9073, mcs1_mcs_mat1_0_mcs_out[104]}), .c ({new_AGEMA_signal_9372, mcs1_mcs_mat1_0_n98}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U48 ( .a ({new_AGEMA_signal_8583, mcs1_mcs_mat1_0_n96}), .b ({new_AGEMA_signal_10315, mcs1_mcs_mat1_0_n95}), .c ({new_AGEMA_signal_10617, mcs_out[191]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U47 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_10079, mcs1_mcs_mat1_0_mcs_out[95]}), .c ({new_AGEMA_signal_10315, mcs1_mcs_mat1_0_n95}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U46 ( .a ({new_AGEMA_signal_8118, mcs1_mcs_mat1_0_mcs_out[83]}), .b ({new_AGEMA_signal_7637, mcs1_mcs_mat1_0_mcs_out[87]}), .c ({new_AGEMA_signal_8583, mcs1_mcs_mat1_0_n96}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U45 ( .a ({new_AGEMA_signal_8584, mcs1_mcs_mat1_0_n94}), .b ({new_AGEMA_signal_9863, mcs1_mcs_mat1_0_n93}), .c ({new_AGEMA_signal_10072, mcs_out[190]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U43 ( .a ({new_AGEMA_signal_8119, mcs1_mcs_mat1_0_mcs_out[82]}), .b ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_8584, mcs1_mcs_mat1_0_n94}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U42 ( .a ({new_AGEMA_signal_8585, mcs1_mcs_mat1_0_n92}), .b ({new_AGEMA_signal_9864, mcs1_mcs_mat1_0_n91}), .c ({new_AGEMA_signal_10073, mcs_out[189]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U41 ( .a ({new_AGEMA_signal_7326, mcs1_mcs_mat1_0_mcs_out[89]}), .b ({new_AGEMA_signal_9630, mcs1_mcs_mat1_0_mcs_out[93]}), .c ({new_AGEMA_signal_9864, mcs1_mcs_mat1_0_n91}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U40 ( .a ({new_AGEMA_signal_8120, mcs1_mcs_mat1_0_mcs_out[81]}), .b ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_8585, mcs1_mcs_mat1_0_n92}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U39 ( .a ({new_AGEMA_signal_9065, mcs1_mcs_mat1_0_n90}), .b ({new_AGEMA_signal_10618, mcs1_mcs_mat1_0_n89}), .c ({new_AGEMA_signal_10872, mcs_out[188]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U38 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_10326, mcs1_mcs_mat1_0_mcs_out[92]}), .c ({new_AGEMA_signal_10618, mcs1_mcs_mat1_0_n89}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U37 ( .a ({new_AGEMA_signal_8605, mcs1_mcs_mat1_0_mcs_out[80]}), .b ({new_AGEMA_signal_8117, mcs1_mcs_mat1_0_mcs_out[84]}), .c ({new_AGEMA_signal_9065, mcs1_mcs_mat1_0_n90}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U36 ( .a ({new_AGEMA_signal_10316, mcs1_mcs_mat1_0_n88}), .b ({new_AGEMA_signal_8586, mcs1_mcs_mat1_0_n87}), .c ({temp_next_s1[29], temp_next_s0[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U35 ( .a ({new_AGEMA_signal_7346, mcs1_mcs_mat1_0_mcs_out[5]}), .b ({new_AGEMA_signal_8155, mcs1_mcs_mat1_0_mcs_out[9]}), .c ({new_AGEMA_signal_8586, mcs1_mcs_mat1_0_n87}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U34 ( .a ({new_AGEMA_signal_10090, mcs1_mcs_mat1_0_mcs_out[13]}), .b ({new_AGEMA_signal_8638, mcs1_mcs_mat1_0_mcs_out[1]}), .c ({new_AGEMA_signal_10316, mcs1_mcs_mat1_0_n88}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U33 ( .a ({new_AGEMA_signal_9373, mcs1_mcs_mat1_0_n86}), .b ({new_AGEMA_signal_10317, mcs1_mcs_mat1_0_n85}), .c ({new_AGEMA_signal_10620, mcs_out[159]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U32 ( .a ({new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[75]}), .b ({new_AGEMA_signal_10081, mcs1_mcs_mat1_0_mcs_out[79]}), .c ({new_AGEMA_signal_10317, mcs1_mcs_mat1_0_n85}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U31 ( .a ({new_AGEMA_signal_9079, mcs1_mcs_mat1_0_mcs_out[67]}), .b ({new_AGEMA_signal_8610, mcs1_mcs_mat1_0_mcs_out[71]}), .c ({new_AGEMA_signal_9373, mcs1_mcs_mat1_0_n86}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U30 ( .a ({new_AGEMA_signal_9375, mcs1_mcs_mat1_0_n84}), .b ({new_AGEMA_signal_9374, mcs1_mcs_mat1_0_n83}), .c ({new_AGEMA_signal_9623, mcs_out[158]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U29 ( .a ({new_AGEMA_signal_9075, mcs1_mcs_mat1_0_mcs_out[74]}), .b ({new_AGEMA_signal_8606, mcs1_mcs_mat1_0_mcs_out[78]}), .c ({new_AGEMA_signal_9374, mcs1_mcs_mat1_0_n83}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U28 ( .a ({new_AGEMA_signal_8613, mcs1_mcs_mat1_0_mcs_out[66]}), .b ({new_AGEMA_signal_9077, mcs1_mcs_mat1_0_mcs_out[70]}), .c ({new_AGEMA_signal_9375, mcs1_mcs_mat1_0_n84}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U27 ( .a ({new_AGEMA_signal_9376, mcs1_mcs_mat1_0_n82}), .b ({new_AGEMA_signal_9865, mcs1_mcs_mat1_0_n81}), .c ({new_AGEMA_signal_10074, mcs_out[157]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U26 ( .a ({new_AGEMA_signal_8123, mcs1_mcs_mat1_0_mcs_out[73]}), .b ({new_AGEMA_signal_9632, mcs1_mcs_mat1_0_mcs_out[77]}), .c ({new_AGEMA_signal_9865, mcs1_mcs_mat1_0_n81}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U25 ( .a ({new_AGEMA_signal_7648, mcs1_mcs_mat1_0_mcs_out[65]}), .b ({new_AGEMA_signal_9078, mcs1_mcs_mat1_0_mcs_out[69]}), .c ({new_AGEMA_signal_9376, mcs1_mcs_mat1_0_n82}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U24 ( .a ({new_AGEMA_signal_9624, mcs1_mcs_mat1_0_n80}), .b ({new_AGEMA_signal_10621, mcs1_mcs_mat1_0_n79}), .c ({new_AGEMA_signal_10873, mcs_out[156]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U23 ( .a ({new_AGEMA_signal_9076, mcs1_mcs_mat1_0_mcs_out[72]}), .b ({new_AGEMA_signal_10327, mcs1_mcs_mat1_0_mcs_out[76]}), .c ({new_AGEMA_signal_10621, mcs1_mcs_mat1_0_n79}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U22 ( .a ({new_AGEMA_signal_9387, mcs1_mcs_mat1_0_mcs_out[64]}), .b ({new_AGEMA_signal_8612, mcs1_mcs_mat1_0_mcs_out[68]}), .c ({new_AGEMA_signal_9624, mcs1_mcs_mat1_0_n80}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U21 ( .a ({new_AGEMA_signal_9066, mcs1_mcs_mat1_0_n78}), .b ({new_AGEMA_signal_10318, mcs1_mcs_mat1_0_n77}), .c ({temp_next_s1[127], temp_next_s0[127]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U20 ( .a ({new_AGEMA_signal_8129, mcs1_mcs_mat1_0_mcs_out[59]}), .b ({new_AGEMA_signal_10083, mcs1_mcs_mat1_0_mcs_out[63]}), .c ({new_AGEMA_signal_10318, mcs1_mcs_mat1_0_n77}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U19 ( .a ({new_AGEMA_signal_7658, mcs1_mcs_mat1_0_mcs_out[51]}), .b ({new_AGEMA_signal_8617, mcs1_mcs_mat1_0_mcs_out[55]}), .c ({new_AGEMA_signal_9066, mcs1_mcs_mat1_0_n78}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U18 ( .a ({new_AGEMA_signal_9377, mcs1_mcs_mat1_0_n76}), .b ({new_AGEMA_signal_10075, mcs1_mcs_mat1_0_n75}), .c ({temp_next_s1[126], temp_next_s0[126]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U17 ( .a ({new_AGEMA_signal_7650, mcs1_mcs_mat1_0_mcs_out[58]}), .b ({new_AGEMA_signal_9872, mcs1_mcs_mat1_0_mcs_out[62]}), .c ({new_AGEMA_signal_10075, mcs1_mcs_mat1_0_n75}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U16 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_9081, mcs1_mcs_mat1_0_mcs_out[54]}), .c ({new_AGEMA_signal_9377, mcs1_mcs_mat1_0_n76}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U15 ( .a ({new_AGEMA_signal_9378, mcs1_mcs_mat1_0_n74}), .b ({new_AGEMA_signal_10076, mcs1_mcs_mat1_0_n73}), .c ({temp_next_s1[125], temp_next_s0[125]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U14 ( .a ({new_AGEMA_signal_8130, mcs1_mcs_mat1_0_mcs_out[57]}), .b ({new_AGEMA_signal_9873, mcs1_mcs_mat1_0_mcs_out[61]}), .c ({new_AGEMA_signal_10076, mcs1_mcs_mat1_0_n73}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U13 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_9082, mcs1_mcs_mat1_0_mcs_out[53]}), .c ({new_AGEMA_signal_9378, mcs1_mcs_mat1_0_n74}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U12 ( .a ({new_AGEMA_signal_9067, mcs1_mcs_mat1_0_n72}), .b ({new_AGEMA_signal_10623, mcs1_mcs_mat1_0_n71}), .c ({temp_next_s1[124], temp_next_s0[124]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U11 ( .a ({new_AGEMA_signal_8616, mcs1_mcs_mat1_0_mcs_out[56]}), .b ({new_AGEMA_signal_10328, mcs1_mcs_mat1_0_mcs_out[60]}), .c ({new_AGEMA_signal_10623, mcs1_mcs_mat1_0_n71}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U10 ( .a ({new_AGEMA_signal_8134, mcs1_mcs_mat1_0_mcs_out[48]}), .b ({new_AGEMA_signal_8619, mcs1_mcs_mat1_0_mcs_out[52]}), .c ({new_AGEMA_signal_9067, mcs1_mcs_mat1_0_n72}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U9 ( .a ({new_AGEMA_signal_9379, mcs1_mcs_mat1_0_n70}), .b ({new_AGEMA_signal_10321, mcs1_mcs_mat1_0_n69}), .c ({temp_next_s1[95], temp_next_s0[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U8 ( .a ({new_AGEMA_signal_8621, mcs1_mcs_mat1_0_mcs_out[43]}), .b ({new_AGEMA_signal_10085, mcs1_mcs_mat1_0_mcs_out[47]}), .c ({new_AGEMA_signal_10321, mcs1_mcs_mat1_0_n69}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U7 ( .a ({new_AGEMA_signal_8625, mcs1_mcs_mat1_0_mcs_out[35]}), .b ({new_AGEMA_signal_9083, mcs1_mcs_mat1_0_mcs_out[39]}), .c ({new_AGEMA_signal_9379, mcs1_mcs_mat1_0_n70}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U6 ( .a ({new_AGEMA_signal_8587, mcs1_mcs_mat1_0_n68}), .b ({new_AGEMA_signal_9625, mcs1_mcs_mat1_0_n67}), .c ({temp_next_s1[94], temp_next_s0[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U5 ( .a ({new_AGEMA_signal_8622, mcs1_mcs_mat1_0_mcs_out[42]}), .b ({new_AGEMA_signal_9389, mcs1_mcs_mat1_0_mcs_out[46]}), .c ({new_AGEMA_signal_9625, mcs1_mcs_mat1_0_n67}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U4 ( .a ({new_AGEMA_signal_8142, mcs1_mcs_mat1_0_mcs_out[34]}), .b ({new_AGEMA_signal_7662, mcs1_mcs_mat1_0_mcs_out[38]}), .c ({new_AGEMA_signal_8587, mcs1_mcs_mat1_0_n68}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U3 ( .a ({new_AGEMA_signal_10875, mcs1_mcs_mat1_0_n66}), .b ({new_AGEMA_signal_9867, mcs1_mcs_mat1_0_n65}), .c ({temp_next_s1[28], temp_next_s0[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U2 ( .a ({new_AGEMA_signal_9643, mcs1_mcs_mat1_0_mcs_out[4]}), .b ({new_AGEMA_signal_9090, mcs1_mcs_mat1_0_mcs_out[8]}), .c ({new_AGEMA_signal_9867, mcs1_mcs_mat1_0_n65}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_U1 ( .a ({new_AGEMA_signal_8639, mcs1_mcs_mat1_0_mcs_out[0]}), .b ({new_AGEMA_signal_10626, mcs1_mcs_mat1_0_mcs_out[12]}), .c ({new_AGEMA_signal_10875, mcs1_mcs_mat1_0_n66}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_8588, mcs1_mcs_mat1_0_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_9068, mcs1_mcs_mat1_0_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_8102, mcs1_mcs_mat1_0_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_6700, mcs1_mcs_mat1_0_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8588, mcs1_mcs_mat1_0_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_6952, mcs1_mcs_mat1_0_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_7312, mcs1_mcs_mat1_0_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_7622, mcs1_mcs_mat1_0_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_6953, mcs1_mcs_mat1_0_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_7233, shiftr_out[95]}), .c ({new_AGEMA_signal_7312, mcs1_mcs_mat1_0_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_8589, mcs1_mcs_mat1_0_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_7233, shiftr_out[95]}), .c ({new_AGEMA_signal_9069, mcs1_mcs_mat1_0_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_8102, mcs1_mcs_mat1_0_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_8589, mcs1_mcs_mat1_0_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_7623, mcs1_mcs_mat1_0_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_7313, mcs1_mcs_mat1_0_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_8102, mcs1_mcs_mat1_0_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_8103, mcs1_mcs_mat1_0_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_8590, mcs1_mcs_mat1_0_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_7623, mcs1_mcs_mat1_0_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_6953, mcs1_mcs_mat1_0_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_8103, mcs1_mcs_mat1_0_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[448]), .c ({new_AGEMA_signal_7623, mcs1_mcs_mat1_0_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[449]), .c ({new_AGEMA_signal_6953, mcs1_mcs_mat1_0_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7233, shiftr_out[95]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[450]), .c ({new_AGEMA_signal_7313, mcs1_mcs_mat1_0_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_8591, mcs1_mcs_mat1_0_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_6693, shiftr_out[62]}), .c ({new_AGEMA_signal_9070, mcs1_mcs_mat1_0_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_8104, mcs1_mcs_mat1_0_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7316, mcs1_mcs_mat1_0_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_8591, mcs1_mcs_mat1_0_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_8592, mcs1_mcs_mat1_0_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_7625, mcs1_mcs_mat1_0_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_9071, mcs1_mcs_mat1_0_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_8104, mcs1_mcs_mat1_0_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7305, shiftr_out[61]}), .c ({new_AGEMA_signal_8592, mcs1_mcs_mat1_0_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_8104, mcs1_mcs_mat1_0_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7624, mcs1_mcs_mat1_0_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_8593, mcs1_mcs_mat1_0_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_7626, mcs1_mcs_mat1_0_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_6954, mcs1_mcs_mat1_0_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_8104, mcs1_mcs_mat1_0_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_7315, mcs1_mcs_mat1_0_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_7625, mcs1_mcs_mat1_0_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_8105, mcs1_mcs_mat1_0_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_6701, mcs1_mcs_mat1_0_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7316, mcs1_mcs_mat1_0_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_7625, mcs1_mcs_mat1_0_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_6954, mcs1_mcs_mat1_0_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_7315, mcs1_mcs_mat1_0_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7305, shiftr_out[61]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[451]), .c ({new_AGEMA_signal_7626, mcs1_mcs_mat1_0_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[452]), .c ({new_AGEMA_signal_6954, mcs1_mcs_mat1_0_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[453]), .c ({new_AGEMA_signal_7316, mcs1_mcs_mat1_0_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_8107, mcs1_mcs_mat1_0_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_6955, mcs1_mcs_mat1_0_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_8594, mcs1_mcs_mat1_0_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_7317, mcs1_mcs_mat1_0_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_7318, mcs1_mcs_mat1_0_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_7627, mcs1_mcs_mat1_0_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_8108, mcs1_mcs_mat1_0_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_8595, mcs1_mcs_mat1_0_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_9072, mcs1_mcs_mat1_0_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_8107, mcs1_mcs_mat1_0_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_8595, mcs1_mcs_mat1_0_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_6702, mcs1_mcs_mat1_0_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_7629, mcs1_mcs_mat1_0_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_8107, mcs1_mcs_mat1_0_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_6956, mcs1_mcs_mat1_0_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_7628, mcs1_mcs_mat1_0_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8108, mcs1_mcs_mat1_0_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7311, shiftr_out[29]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[454]), .c ({new_AGEMA_signal_7629, mcs1_mcs_mat1_0_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[455]), .c ({new_AGEMA_signal_6956, mcs1_mcs_mat1_0_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[456]), .c ({new_AGEMA_signal_7318, mcs1_mcs_mat1_0_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({new_AGEMA_signal_10077, mcs1_mcs_mat1_0_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_10322, mcs1_mcs_mat1_0_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({new_AGEMA_signal_10078, mcs1_mcs_mat1_0_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_10323, mcs1_mcs_mat1_0_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_9381, mcs1_mcs_mat1_0_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_10077, mcs1_mcs_mat1_0_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_10324, mcs1_mcs_mat1_0_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_8596, mcs1_mcs_mat1_0_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_9868, mcs1_mcs_mat1_0_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_10077, mcs1_mcs_mat1_0_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_9626, mcs1_mcs_mat1_0_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_10078, mcs1_mcs_mat1_0_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_10325, mcs1_mcs_mat1_0_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_9869, mcs1_mcs_mat1_0_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_10078, mcs1_mcs_mat1_0_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_9381, mcs1_mcs_mat1_0_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_9627, mcs1_mcs_mat1_0_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_9869, mcs1_mcs_mat1_0_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[457]), .c ({new_AGEMA_signal_9627, mcs1_mcs_mat1_0_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[458]), .c ({new_AGEMA_signal_8596, mcs1_mcs_mat1_0_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[459]), .c ({new_AGEMA_signal_9381, mcs1_mcs_mat1_0_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_8111, mcs1_mcs_mat1_0_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_8110, mcs1_mcs_mat1_0_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_8110, mcs1_mcs_mat1_0_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_7319, mcs1_mcs_mat1_0_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_8598, mcs1_mcs_mat1_0_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_6957, mcs1_mcs_mat1_0_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7233, shiftr_out[95]}), .c ({new_AGEMA_signal_7319, mcs1_mcs_mat1_0_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_8110, mcs1_mcs_mat1_0_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8599, mcs1_mcs_mat1_0_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_7631, mcs1_mcs_mat1_0_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_6703, mcs1_mcs_mat1_0_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_8110, mcs1_mcs_mat1_0_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_8600, mcs1_mcs_mat1_0_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_9073, mcs1_mcs_mat1_0_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_8111, mcs1_mcs_mat1_0_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_7631, mcs1_mcs_mat1_0_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_8600, mcs1_mcs_mat1_0_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_7630, mcs1_mcs_mat1_0_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_6619, shiftr_out[92]}), .c ({new_AGEMA_signal_8111, mcs1_mcs_mat1_0_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_6957, mcs1_mcs_mat1_0_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7320, mcs1_mcs_mat1_0_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_7630, mcs1_mcs_mat1_0_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[460]), .c ({new_AGEMA_signal_7631, mcs1_mcs_mat1_0_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[461]), .c ({new_AGEMA_signal_6957, mcs1_mcs_mat1_0_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7233, shiftr_out[95]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[462]), .c ({new_AGEMA_signal_7320, mcs1_mcs_mat1_0_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_7321, mcs1_mcs_mat1_0_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_8112, mcs1_mcs_mat1_0_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_8601, mcs1_mcs_mat1_0_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_7635, mcs1_mcs_mat1_0_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_8112, mcs1_mcs_mat1_0_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_7633, mcs1_mcs_mat1_0_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_7322, mcs1_mcs_mat1_0_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_8113, mcs1_mcs_mat1_0_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_7634, mcs1_mcs_mat1_0_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_8114, mcs1_mcs_mat1_0_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_8602, mcs1_mcs_mat1_0_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_6704, mcs1_mcs_mat1_0_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7635, mcs1_mcs_mat1_0_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_8114, mcs1_mcs_mat1_0_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_6958, mcs1_mcs_mat1_0_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_7305, shiftr_out[61]}), .c ({new_AGEMA_signal_7634, mcs1_mcs_mat1_0_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7305, shiftr_out[61]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[463]), .c ({new_AGEMA_signal_7635, mcs1_mcs_mat1_0_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[464]), .c ({new_AGEMA_signal_6958, mcs1_mcs_mat1_0_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[465]), .c ({new_AGEMA_signal_7322, mcs1_mcs_mat1_0_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_9382, mcs1_mcs_mat1_0_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_7324, mcs1_mcs_mat1_0_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_9628, mcs1_mcs_mat1_0_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_9074, mcs1_mcs_mat1_0_mcs_out[99]}), .b ({new_AGEMA_signal_6699, shiftr_out[30]}), .c ({new_AGEMA_signal_9382, mcs1_mcs_mat1_0_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_8603, mcs1_mcs_mat1_0_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_7311, shiftr_out[29]}), .c ({new_AGEMA_signal_9074, mcs1_mcs_mat1_0_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_8115, mcs1_mcs_mat1_0_mcs_out[98]}), .b ({new_AGEMA_signal_6960, mcs1_mcs_mat1_0_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_8603, mcs1_mcs_mat1_0_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_6959, mcs1_mcs_mat1_0_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_7636, mcs1_mcs_mat1_0_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_8115, mcs1_mcs_mat1_0_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7311, shiftr_out[29]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[466]), .c ({new_AGEMA_signal_7636, mcs1_mcs_mat1_0_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[467]), .c ({new_AGEMA_signal_6960, mcs1_mcs_mat1_0_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[468]), .c ({new_AGEMA_signal_7324, mcs1_mcs_mat1_0_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_9870, mcs1_mcs_mat1_0_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_10079, mcs1_mcs_mat1_0_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_9384, mcs1_mcs_mat1_0_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_9385, mcs1_mcs_mat1_0_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_9630, mcs1_mcs_mat1_0_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_10080, mcs1_mcs_mat1_0_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_8604, mcs1_mcs_mat1_0_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_10326, mcs1_mcs_mat1_0_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_9870, mcs1_mcs_mat1_0_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_10080, mcs1_mcs_mat1_0_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_8116, mcs1_mcs_mat1_0_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_9631, mcs1_mcs_mat1_0_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_9870, mcs1_mcs_mat1_0_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[469]), .c ({new_AGEMA_signal_9631, mcs1_mcs_mat1_0_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[470]), .c ({new_AGEMA_signal_8604, mcs1_mcs_mat1_0_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[471]), .c ({new_AGEMA_signal_9385, mcs1_mcs_mat1_0_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_7640, mcs1_mcs_mat1_0_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_7641, mcs1_mcs_mat1_0_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_8118, mcs1_mcs_mat1_0_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_7638, mcs1_mcs_mat1_0_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_6706, mcs1_mcs_mat1_0_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_8119, mcs1_mcs_mat1_0_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_7327, mcs1_mcs_mat1_0_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_7638, mcs1_mcs_mat1_0_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_7639, mcs1_mcs_mat1_0_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_8120, mcs1_mcs_mat1_0_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_6961, mcs1_mcs_mat1_0_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_7327, mcs1_mcs_mat1_0_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_7639, mcs1_mcs_mat1_0_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_8121, mcs1_mcs_mat1_0_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_6699, shiftr_out[30]}), .c ({new_AGEMA_signal_8605, mcs1_mcs_mat1_0_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_7640, mcs1_mcs_mat1_0_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_6961, mcs1_mcs_mat1_0_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_8121, mcs1_mcs_mat1_0_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7311, shiftr_out[29]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[472]), .c ({new_AGEMA_signal_7641, mcs1_mcs_mat1_0_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[473]), .c ({new_AGEMA_signal_6961, mcs1_mcs_mat1_0_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[474]), .c ({new_AGEMA_signal_7327, mcs1_mcs_mat1_0_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_9871, mcs1_mcs_mat1_0_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_10081, mcs1_mcs_mat1_0_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_9386, mcs1_mcs_mat1_0_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_9632, mcs1_mcs_mat1_0_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_10082, mcs1_mcs_mat1_0_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_8607, mcs1_mcs_mat1_0_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_10327, mcs1_mcs_mat1_0_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_9871, mcs1_mcs_mat1_0_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7615, shiftr_out[124]}), .c ({new_AGEMA_signal_10082, mcs1_mcs_mat1_0_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_8122, mcs1_mcs_mat1_0_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_9633, mcs1_mcs_mat1_0_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_9871, mcs1_mcs_mat1_0_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[475]), .c ({new_AGEMA_signal_9633, mcs1_mcs_mat1_0_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[476]), .c ({new_AGEMA_signal_8607, mcs1_mcs_mat1_0_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[477]), .c ({new_AGEMA_signal_9386, mcs1_mcs_mat1_0_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_8608, mcs1_mcs_mat1_0_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_9075, mcs1_mcs_mat1_0_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_8124, mcs1_mcs_mat1_0_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7643, mcs1_mcs_mat1_0_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_8608, mcs1_mcs_mat1_0_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_7246, mcs1_mcs_mat1_0_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_7643, mcs1_mcs_mat1_0_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_7246, mcs1_mcs_mat1_0_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_8123, mcs1_mcs_mat1_0_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_6962, mcs1_mcs_mat1_0_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_6963, mcs1_mcs_mat1_0_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_7246, mcs1_mcs_mat1_0_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_7328, mcs1_mcs_mat1_0_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_6619, shiftr_out[92]}), .c ({new_AGEMA_signal_7643, mcs1_mcs_mat1_0_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_8609, mcs1_mcs_mat1_0_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_6962, mcs1_mcs_mat1_0_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_9076, mcs1_mcs_mat1_0_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_8124, mcs1_mcs_mat1_0_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7328, mcs1_mcs_mat1_0_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_8609, mcs1_mcs_mat1_0_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_7233, shiftr_out[95]}), .b ({new_AGEMA_signal_7644, mcs1_mcs_mat1_0_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_8124, mcs1_mcs_mat1_0_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[478]), .c ({new_AGEMA_signal_7644, mcs1_mcs_mat1_0_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[479]), .c ({new_AGEMA_signal_6963, mcs1_mcs_mat1_0_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7233, shiftr_out[95]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[480]), .c ({new_AGEMA_signal_7328, mcs1_mcs_mat1_0_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_8125, mcs1_mcs_mat1_0_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_7329, mcs1_mcs_mat1_0_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_8610, mcs1_mcs_mat1_0_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_7646, mcs1_mcs_mat1_0_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_8611, mcs1_mcs_mat1_0_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9077, mcs1_mcs_mat1_0_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_8125, mcs1_mcs_mat1_0_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_8611, mcs1_mcs_mat1_0_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9078, mcs1_mcs_mat1_0_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_7329, mcs1_mcs_mat1_0_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_8126, mcs1_mcs_mat1_0_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_8611, mcs1_mcs_mat1_0_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({new_AGEMA_signal_6964, mcs1_mcs_mat1_0_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_7329, mcs1_mcs_mat1_0_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_7645, mcs1_mcs_mat1_0_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_7305, shiftr_out[61]}), .c ({new_AGEMA_signal_8125, mcs1_mcs_mat1_0_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_7330, mcs1_mcs_mat1_0_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6708, mcs1_mcs_mat1_0_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_7645, mcs1_mcs_mat1_0_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_8126, mcs1_mcs_mat1_0_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_7646, mcs1_mcs_mat1_0_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_8612, mcs1_mcs_mat1_0_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_7330, mcs1_mcs_mat1_0_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_7646, mcs1_mcs_mat1_0_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({new_AGEMA_signal_7647, mcs1_mcs_mat1_0_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_8126, mcs1_mcs_mat1_0_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7305, shiftr_out[61]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[481]), .c ({new_AGEMA_signal_7647, mcs1_mcs_mat1_0_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[482]), .c ({new_AGEMA_signal_6964, mcs1_mcs_mat1_0_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[483]), .c ({new_AGEMA_signal_7330, mcs1_mcs_mat1_0_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_8614, mcs1_mcs_mat1_0_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_9079, mcs1_mcs_mat1_0_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({new_AGEMA_signal_8127, mcs1_mcs_mat1_0_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_8613, mcs1_mcs_mat1_0_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_9080, mcs1_mcs_mat1_0_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_7331, mcs1_mcs_mat1_0_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_9387, mcs1_mcs_mat1_0_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_8614, mcs1_mcs_mat1_0_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .c ({new_AGEMA_signal_9080, mcs1_mcs_mat1_0_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_6965, mcs1_mcs_mat1_0_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_8127, mcs1_mcs_mat1_0_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_8614, mcs1_mcs_mat1_0_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_6709, mcs1_mcs_mat1_0_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7649, mcs1_mcs_mat1_0_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_8127, mcs1_mcs_mat1_0_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7311, shiftr_out[29]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[484]), .c ({new_AGEMA_signal_7649, mcs1_mcs_mat1_0_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[485]), .c ({new_AGEMA_signal_6965, mcs1_mcs_mat1_0_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[486]), .c ({new_AGEMA_signal_7331, mcs1_mcs_mat1_0_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_9874, mcs1_mcs_mat1_0_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_9388, mcs1_mcs_mat1_0_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_10083, mcs1_mcs_mat1_0_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_8615, mcs1_mcs_mat1_0_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_9634, mcs1_mcs_mat1_0_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_9872, mcs1_mcs_mat1_0_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({new_AGEMA_signal_9635, mcs1_mcs_mat1_0_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_9873, mcs1_mcs_mat1_0_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[487]), .c ({new_AGEMA_signal_9635, mcs1_mcs_mat1_0_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[488]), .c ({new_AGEMA_signal_8615, mcs1_mcs_mat1_0_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[489]), .c ({new_AGEMA_signal_9388, mcs1_mcs_mat1_0_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_6967, mcs1_mcs_mat1_0_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_7332, mcs1_mcs_mat1_0_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_7650, mcs1_mcs_mat1_0_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_6968, mcs1_mcs_mat1_0_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_7651, mcs1_mcs_mat1_0_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_8130, mcs1_mcs_mat1_0_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_8131, mcs1_mcs_mat1_0_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_7652, mcs1_mcs_mat1_0_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_8616, mcs1_mcs_mat1_0_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_7653, mcs1_mcs_mat1_0_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_8131, mcs1_mcs_mat1_0_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[490]), .c ({new_AGEMA_signal_7653, mcs1_mcs_mat1_0_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[491]), .c ({new_AGEMA_signal_6968, mcs1_mcs_mat1_0_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7233, shiftr_out[95]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[492]), .c ({new_AGEMA_signal_7332, mcs1_mcs_mat1_0_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_7655, mcs1_mcs_mat1_0_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8132, mcs1_mcs_mat1_0_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_8617, mcs1_mcs_mat1_0_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_8618, mcs1_mcs_mat1_0_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_7654, mcs1_mcs_mat1_0_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_9081, mcs1_mcs_mat1_0_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_7333, mcs1_mcs_mat1_0_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_7654, mcs1_mcs_mat1_0_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({new_AGEMA_signal_8618, mcs1_mcs_mat1_0_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_9082, mcs1_mcs_mat1_0_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_6711, mcs1_mcs_mat1_0_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_8132, mcs1_mcs_mat1_0_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_8618, mcs1_mcs_mat1_0_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_6969, mcs1_mcs_mat1_0_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_7657, mcs1_mcs_mat1_0_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_8132, mcs1_mcs_mat1_0_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_7656, mcs1_mcs_mat1_0_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_8133, mcs1_mcs_mat1_0_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_8619, mcs1_mcs_mat1_0_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_7655, mcs1_mcs_mat1_0_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_6969, mcs1_mcs_mat1_0_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_8133, mcs1_mcs_mat1_0_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_7333, mcs1_mcs_mat1_0_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_7655, mcs1_mcs_mat1_0_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7305, shiftr_out[61]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[493]), .c ({new_AGEMA_signal_7657, mcs1_mcs_mat1_0_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[494]), .c ({new_AGEMA_signal_6969, mcs1_mcs_mat1_0_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[495]), .c ({new_AGEMA_signal_7333, mcs1_mcs_mat1_0_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_9390, mcs1_mcs_mat1_0_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_9636, mcs1_mcs_mat1_0_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_10329, mcs1_mcs_mat1_0_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_8620, mcs1_mcs_mat1_0_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_10625, mcs1_mcs_mat1_0_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_10085, mcs1_mcs_mat1_0_mcs_out[47]}), .b ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_10329, mcs1_mcs_mat1_0_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_9875, mcs1_mcs_mat1_0_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_7615, shiftr_out[124]}), .c ({new_AGEMA_signal_10085, mcs1_mcs_mat1_0_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_8135, mcs1_mcs_mat1_0_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_9637, mcs1_mcs_mat1_0_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_9875, mcs1_mcs_mat1_0_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[496]), .c ({new_AGEMA_signal_9637, mcs1_mcs_mat1_0_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[497]), .c ({new_AGEMA_signal_8620, mcs1_mcs_mat1_0_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[498]), .c ({new_AGEMA_signal_9390, mcs1_mcs_mat1_0_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_8136, mcs1_mcs_mat1_0_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_7334, mcs1_mcs_mat1_0_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_8621, mcs1_mcs_mat1_0_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_7659, mcs1_mcs_mat1_0_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_6970, mcs1_mcs_mat1_0_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_8136, mcs1_mcs_mat1_0_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_8137, mcs1_mcs_mat1_0_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_7661, mcs1_mcs_mat1_0_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_8622, mcs1_mcs_mat1_0_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_8138, mcs1_mcs_mat1_0_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_6712, mcs1_mcs_mat1_0_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_8623, mcs1_mcs_mat1_0_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_7659, mcs1_mcs_mat1_0_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7335, mcs1_mcs_mat1_0_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8138, mcs1_mcs_mat1_0_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_7660, mcs1_mcs_mat1_0_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_7335, mcs1_mcs_mat1_0_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8139, mcs1_mcs_mat1_0_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[499]), .c ({new_AGEMA_signal_7661, mcs1_mcs_mat1_0_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[500]), .c ({new_AGEMA_signal_6970, mcs1_mcs_mat1_0_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7233, shiftr_out[95]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[501]), .c ({new_AGEMA_signal_7335, mcs1_mcs_mat1_0_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_8624, mcs1_mcs_mat1_0_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_6713, mcs1_mcs_mat1_0_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9083, mcs1_mcs_mat1_0_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_7337, mcs1_mcs_mat1_0_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_7336, mcs1_mcs_mat1_0_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_7662, mcs1_mcs_mat1_0_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({new_AGEMA_signal_8624, mcs1_mcs_mat1_0_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_9084, mcs1_mcs_mat1_0_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_7663, mcs1_mcs_mat1_0_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_8140, mcs1_mcs_mat1_0_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_8624, mcs1_mcs_mat1_0_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_7664, mcs1_mcs_mat1_0_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7338, mcs1_mcs_mat1_0_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_8140, mcs1_mcs_mat1_0_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_7664, mcs1_mcs_mat1_0_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7337, mcs1_mcs_mat1_0_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_8141, mcs1_mcs_mat1_0_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_7247, mcs1_mcs_mat1_0_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_7337, mcs1_mcs_mat1_0_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({new_AGEMA_signal_6971, mcs1_mcs_mat1_0_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_7247, mcs1_mcs_mat1_0_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7305, shiftr_out[61]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[502]), .c ({new_AGEMA_signal_7664, mcs1_mcs_mat1_0_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[503]), .c ({new_AGEMA_signal_6971, mcs1_mcs_mat1_0_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[504]), .c ({new_AGEMA_signal_7338, mcs1_mcs_mat1_0_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_7665, mcs1_mcs_mat1_0_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7339, mcs1_mcs_mat1_0_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_8142, mcs1_mcs_mat1_0_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_6972, mcs1_mcs_mat1_0_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_7248, mcs1_mcs_mat1_0_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_9085, mcs1_mcs_mat1_0_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_7666, mcs1_mcs_mat1_0_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_9391, mcs1_mcs_mat1_0_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7311, shiftr_out[29]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[505]), .c ({new_AGEMA_signal_7666, mcs1_mcs_mat1_0_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[506]), .c ({new_AGEMA_signal_6972, mcs1_mcs_mat1_0_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[507]), .c ({new_AGEMA_signal_7339, mcs1_mcs_mat1_0_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_10086, mcs1_mcs_mat1_0_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_9876, mcs1_mcs_mat1_0_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_10330, mcs1_mcs_mat1_0_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_8627, mcs1_mcs_mat1_0_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_9877, mcs1_mcs_mat1_0_mcs_out[29]}), .c ({new_AGEMA_signal_10086, mcs1_mcs_mat1_0_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_8626, mcs1_mcs_mat1_0_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_9876, mcs1_mcs_mat1_0_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_10087, mcs1_mcs_mat1_0_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_9640, mcs1_mcs_mat1_0_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7615, shiftr_out[124]}), .c ({new_AGEMA_signal_9876, mcs1_mcs_mat1_0_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_10088, mcs1_mcs_mat1_0_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_9638, mcs1_mcs_mat1_0_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_10331, mcs1_mcs_mat1_0_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_9878, mcs1_mcs_mat1_0_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_9639, mcs1_mcs_mat1_0_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_10088, mcs1_mcs_mat1_0_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_9392, mcs1_mcs_mat1_0_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_9639, mcs1_mcs_mat1_0_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_9640, mcs1_mcs_mat1_0_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8627, mcs1_mcs_mat1_0_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_9878, mcs1_mcs_mat1_0_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[508]), .c ({new_AGEMA_signal_9640, mcs1_mcs_mat1_0_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[509]), .c ({new_AGEMA_signal_8627, mcs1_mcs_mat1_0_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[510]), .c ({new_AGEMA_signal_9392, mcs1_mcs_mat1_0_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_7667, mcs1_mcs_mat1_0_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_8145, mcs1_mcs_mat1_0_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_7340, mcs1_mcs_mat1_0_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_6973, mcs1_mcs_mat1_0_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_7667, mcs1_mcs_mat1_0_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_8146, mcs1_mcs_mat1_0_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_8628, mcs1_mcs_mat1_0_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_7669, mcs1_mcs_mat1_0_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_6973, mcs1_mcs_mat1_0_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_8146, mcs1_mcs_mat1_0_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_8629, mcs1_mcs_mat1_0_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_6619, shiftr_out[92]}), .c ({new_AGEMA_signal_9086, mcs1_mcs_mat1_0_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_7669, mcs1_mcs_mat1_0_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8147, mcs1_mcs_mat1_0_mcs_out[24]}), .c ({new_AGEMA_signal_8629, mcs1_mcs_mat1_0_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_7668, mcs1_mcs_mat1_0_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_7233, shiftr_out[95]}), .c ({new_AGEMA_signal_8147, mcs1_mcs_mat1_0_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_7340, mcs1_mcs_mat1_0_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_6715, mcs1_mcs_mat1_0_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_7668, mcs1_mcs_mat1_0_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[511]), .c ({new_AGEMA_signal_7669, mcs1_mcs_mat1_0_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[512]), .c ({new_AGEMA_signal_6973, mcs1_mcs_mat1_0_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7233, shiftr_out[95]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[513]), .c ({new_AGEMA_signal_7340, mcs1_mcs_mat1_0_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_7670, mcs1_mcs_mat1_0_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_6693, shiftr_out[62]}), .c ({new_AGEMA_signal_8148, mcs1_mcs_mat1_0_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_7341, mcs1_mcs_mat1_0_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_6974, mcs1_mcs_mat1_0_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_7670, mcs1_mcs_mat1_0_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_8149, mcs1_mcs_mat1_0_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_7305, shiftr_out[61]}), .c ({new_AGEMA_signal_8630, mcs1_mcs_mat1_0_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_7672, mcs1_mcs_mat1_0_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_6974, mcs1_mcs_mat1_0_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_8149, mcs1_mcs_mat1_0_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_8631, mcs1_mcs_mat1_0_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_6625, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_9087, mcs1_mcs_mat1_0_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_7672, mcs1_mcs_mat1_0_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8150, mcs1_mcs_mat1_0_mcs_out[20]}), .c ({new_AGEMA_signal_8631, mcs1_mcs_mat1_0_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_7671, mcs1_mcs_mat1_0_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_8150, mcs1_mcs_mat1_0_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_7341, mcs1_mcs_mat1_0_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_6716, mcs1_mcs_mat1_0_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_7671, mcs1_mcs_mat1_0_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7305, shiftr_out[61]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[514]), .c ({new_AGEMA_signal_7672, mcs1_mcs_mat1_0_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[515]), .c ({new_AGEMA_signal_6974, mcs1_mcs_mat1_0_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[516]), .c ({new_AGEMA_signal_7341, mcs1_mcs_mat1_0_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_7673, mcs1_mcs_mat1_0_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_7676, mcs1_mcs_mat1_0_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_8151, mcs1_mcs_mat1_0_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_8152, mcs1_mcs_mat1_0_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_6717, mcs1_mcs_mat1_0_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_8632, mcs1_mcs_mat1_0_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_8633, mcs1_mcs_mat1_0_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_6975, mcs1_mcs_mat1_0_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_9088, mcs1_mcs_mat1_0_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_6631, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_8152, mcs1_mcs_mat1_0_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_8633, mcs1_mcs_mat1_0_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_7674, mcs1_mcs_mat1_0_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_7311, shiftr_out[29]}), .c ({new_AGEMA_signal_8152, mcs1_mcs_mat1_0_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_7342, mcs1_mcs_mat1_0_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_7343, mcs1_mcs_mat1_0_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_7674, mcs1_mcs_mat1_0_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_7675, mcs1_mcs_mat1_0_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_6975, mcs1_mcs_mat1_0_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_8153, mcs1_mcs_mat1_0_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7311, shiftr_out[29]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[517]), .c ({new_AGEMA_signal_7676, mcs1_mcs_mat1_0_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[518]), .c ({new_AGEMA_signal_6975, mcs1_mcs_mat1_0_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[519]), .c ({new_AGEMA_signal_7343, mcs1_mcs_mat1_0_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_10091, mcs1_mcs_mat1_0_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_9089, mcs1_mcs_mat1_0_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_10332, mcs1_mcs_mat1_0_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_9881, mcs1_mcs_mat1_0_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_9879, mcs1_mcs_mat1_0_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_10089, mcs1_mcs_mat1_0_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_9642, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_8634, mcs1_mcs_mat1_0_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_9879, mcs1_mcs_mat1_0_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_9089, mcs1_mcs_mat1_0_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_9880, mcs1_mcs_mat1_0_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_10090, mcs1_mcs_mat1_0_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_9641, mcs1_mcs_mat1_0_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_9642, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_9880, mcs1_mcs_mat1_0_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_8154, mcs1_mcs_mat1_0_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_8634, mcs1_mcs_mat1_0_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_9089, mcs1_mcs_mat1_0_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_10333, mcs1_mcs_mat1_0_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_10626, mcs1_mcs_mat1_0_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_10091, mcs1_mcs_mat1_0_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_9642, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_10333, mcs1_mcs_mat1_0_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_9881, mcs1_mcs_mat1_0_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_10091, mcs1_mcs_mat1_0_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_9641, mcs1_mcs_mat1_0_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_9881, mcs1_mcs_mat1_0_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_7615, shiftr_out[124]}), .b ({new_AGEMA_signal_9393, mcs1_mcs_mat1_0_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_9641, mcs1_mcs_mat1_0_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9357, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[520]), .c ({new_AGEMA_signal_9642, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8095, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[521]), .c ({new_AGEMA_signal_8634, mcs1_mcs_mat1_0_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9053, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[522]), .c ({new_AGEMA_signal_9393, mcs1_mcs_mat1_0_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_7249, mcs1_mcs_mat1_0_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_7233, shiftr_out[95]}), .c ({new_AGEMA_signal_7344, mcs1_mcs_mat1_0_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_8156, mcs1_mcs_mat1_0_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_8635, mcs1_mcs_mat1_0_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_7677, mcs1_mcs_mat1_0_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_8155, mcs1_mcs_mat1_0_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_7345, mcs1_mcs_mat1_0_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_7249, mcs1_mcs_mat1_0_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_7677, mcs1_mcs_mat1_0_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_6718, mcs1_mcs_mat1_0_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_6976, mcs1_mcs_mat1_0_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_7249, mcs1_mcs_mat1_0_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_8636, mcs1_mcs_mat1_0_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_6619, shiftr_out[92]}), .c ({new_AGEMA_signal_9090, mcs1_mcs_mat1_0_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_6718, mcs1_mcs_mat1_0_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8156, mcs1_mcs_mat1_0_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_8636, mcs1_mcs_mat1_0_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_7678, mcs1_mcs_mat1_0_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_7345, mcs1_mcs_mat1_0_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_8156, mcs1_mcs_mat1_0_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7299, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[523]), .c ({new_AGEMA_signal_7678, mcs1_mcs_mat1_0_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6687, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[524]), .c ({new_AGEMA_signal_6976, mcs1_mcs_mat1_0_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7233, shiftr_out[95]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[525]), .c ({new_AGEMA_signal_7345, mcs1_mcs_mat1_0_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_9394, mcs1_mcs_mat1_0_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_7347, mcs1_mcs_mat1_0_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_9643, mcs1_mcs_mat1_0_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_9091, mcs1_mcs_mat1_0_mcs_out[7]}), .b ({new_AGEMA_signal_6693, shiftr_out[62]}), .c ({new_AGEMA_signal_9394, mcs1_mcs_mat1_0_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_8637, mcs1_mcs_mat1_0_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_7305, shiftr_out[61]}), .c ({new_AGEMA_signal_9091, mcs1_mcs_mat1_0_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_8157, mcs1_mcs_mat1_0_mcs_out[6]}), .b ({new_AGEMA_signal_6978, mcs1_mcs_mat1_0_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_8637, mcs1_mcs_mat1_0_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_6977, mcs1_mcs_mat1_0_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_7679, mcs1_mcs_mat1_0_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_8157, mcs1_mcs_mat1_0_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7305, shiftr_out[61]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[526]), .c ({new_AGEMA_signal_7679, mcs1_mcs_mat1_0_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6693, shiftr_out[62]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[527]), .c ({new_AGEMA_signal_6978, mcs1_mcs_mat1_0_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7239, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[528]), .c ({new_AGEMA_signal_7347, mcs1_mcs_mat1_0_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_7348, mcs1_mcs_mat1_0_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_7680, mcs1_mcs_mat1_0_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_8159, mcs1_mcs_mat1_0_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_7311, shiftr_out[29]}), .b ({new_AGEMA_signal_7349, mcs1_mcs_mat1_0_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_7680, mcs1_mcs_mat1_0_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_8160, mcs1_mcs_mat1_0_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_6979, mcs1_mcs_mat1_0_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_8638, mcs1_mcs_mat1_0_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_8161, mcs1_mcs_mat1_0_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_7682, mcs1_mcs_mat1_0_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_8639, mcs1_mcs_mat1_0_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_7683, mcs1_mcs_mat1_0_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_6720, mcs1_mcs_mat1_0_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8161, mcs1_mcs_mat1_0_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7311, shiftr_out[29]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[529]), .c ({new_AGEMA_signal_7683, mcs1_mcs_mat1_0_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6699, shiftr_out[30]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[530]), .c ({new_AGEMA_signal_6979, mcs1_mcs_mat1_0_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7245, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[531]), .c ({new_AGEMA_signal_7349, mcs1_mcs_mat1_0_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U96 ( .a ({new_AGEMA_signal_9395, mcs1_mcs_mat1_1_n128}), .b ({new_AGEMA_signal_9092, mcs1_mcs_mat1_1_n127}), .c ({temp_next_s1[89], temp_next_s0[89]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U95 ( .a ({new_AGEMA_signal_8682, mcs1_mcs_mat1_1_mcs_out[41]}), .b ({new_AGEMA_signal_7719, mcs1_mcs_mat1_1_mcs_out[45]}), .c ({new_AGEMA_signal_9092, mcs1_mcs_mat1_1_n127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U94 ( .a ({new_AGEMA_signal_9125, mcs1_mcs_mat1_1_mcs_out[33]}), .b ({new_AGEMA_signal_9124, mcs1_mcs_mat1_1_mcs_out[37]}), .c ({new_AGEMA_signal_9395, mcs1_mcs_mat1_1_n128}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U93 ( .a ({new_AGEMA_signal_10876, mcs1_mcs_mat1_1_n126}), .b ({new_AGEMA_signal_9645, mcs1_mcs_mat1_1_n125}), .c ({temp_next_s1[88], temp_next_s0[88]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U92 ( .a ({new_AGEMA_signal_8199, mcs1_mcs_mat1_1_mcs_out[40]}), .b ({new_AGEMA_signal_9415, mcs1_mcs_mat1_1_mcs_out[44]}), .c ({new_AGEMA_signal_9645, mcs1_mcs_mat1_1_n125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U91 ( .a ({new_AGEMA_signal_10640, mcs1_mcs_mat1_1_mcs_out[32]}), .b ({new_AGEMA_signal_8201, mcs1_mcs_mat1_1_mcs_out[36]}), .c ({new_AGEMA_signal_10876, mcs1_mcs_mat1_1_n126}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U90 ( .a ({new_AGEMA_signal_10092, mcs1_mcs_mat1_1_n124}), .b ({new_AGEMA_signal_9396, mcs1_mcs_mat1_1_n123}), .c ({temp_next_s1[59], temp_next_s0[59]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U89 ( .a ({new_AGEMA_signal_8206, mcs1_mcs_mat1_1_mcs_out[27]}), .b ({new_AGEMA_signal_9126, mcs1_mcs_mat1_1_mcs_out[31]}), .c ({new_AGEMA_signal_9396, mcs1_mcs_mat1_1_n123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U88 ( .a ({new_AGEMA_signal_9899, mcs1_mcs_mat1_1_mcs_out[19]}), .b ({new_AGEMA_signal_8209, mcs1_mcs_mat1_1_mcs_out[23]}), .c ({new_AGEMA_signal_10092, mcs1_mcs_mat1_1_n124}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U87 ( .a ({new_AGEMA_signal_10335, mcs1_mcs_mat1_1_n122}), .b ({new_AGEMA_signal_9093, mcs1_mcs_mat1_1_n121}), .c ({temp_next_s1[58], temp_next_s0[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U86 ( .a ({new_AGEMA_signal_8688, mcs1_mcs_mat1_1_mcs_out[26]}), .b ({new_AGEMA_signal_8686, mcs1_mcs_mat1_1_mcs_out[30]}), .c ({new_AGEMA_signal_9093, mcs1_mcs_mat1_1_n121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U85 ( .a ({new_AGEMA_signal_10113, mcs1_mcs_mat1_1_mcs_out[18]}), .b ({new_AGEMA_signal_8690, mcs1_mcs_mat1_1_mcs_out[22]}), .c ({new_AGEMA_signal_10335, mcs1_mcs_mat1_1_n122}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U84 ( .a ({new_AGEMA_signal_10628, mcs1_mcs_mat1_1_n120}), .b ({new_AGEMA_signal_9397, mcs1_mcs_mat1_1_n119}), .c ({temp_next_s1[57], temp_next_s0[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U83 ( .a ({new_AGEMA_signal_9128, mcs1_mcs_mat1_1_mcs_out[25]}), .b ({new_AGEMA_signal_8204, mcs1_mcs_mat1_1_mcs_out[29]}), .c ({new_AGEMA_signal_9397, mcs1_mcs_mat1_1_n119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U82 ( .a ({new_AGEMA_signal_10357, mcs1_mcs_mat1_1_mcs_out[17]}), .b ({new_AGEMA_signal_9129, mcs1_mcs_mat1_1_mcs_out[21]}), .c ({new_AGEMA_signal_10628, mcs1_mcs_mat1_1_n120}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U81 ( .a ({new_AGEMA_signal_10093, mcs1_mcs_mat1_1_n118}), .b ({new_AGEMA_signal_9398, mcs1_mcs_mat1_1_n117}), .c ({temp_next_s1[56], temp_next_s0[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U80 ( .a ({new_AGEMA_signal_8208, mcs1_mcs_mat1_1_mcs_out[24]}), .b ({new_AGEMA_signal_9127, mcs1_mcs_mat1_1_mcs_out[28]}), .c ({new_AGEMA_signal_9398, mcs1_mcs_mat1_1_n117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U79 ( .a ({new_AGEMA_signal_9901, mcs1_mcs_mat1_1_mcs_out[16]}), .b ({new_AGEMA_signal_8211, mcs1_mcs_mat1_1_mcs_out[20]}), .c ({new_AGEMA_signal_10093, mcs1_mcs_mat1_1_n118}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U78 ( .a ({new_AGEMA_signal_9399, mcs1_mcs_mat1_1_n116}), .b ({new_AGEMA_signal_10094, mcs1_mcs_mat1_1_n115}), .c ({temp_next_s1[27], temp_next_s0[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U77 ( .a ({new_AGEMA_signal_9902, mcs1_mcs_mat1_1_mcs_out[3]}), .b ({new_AGEMA_signal_9133, mcs1_mcs_mat1_1_mcs_out[7]}), .c ({new_AGEMA_signal_10094, mcs1_mcs_mat1_1_n115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U76 ( .a ({new_AGEMA_signal_7384, mcs1_mcs_mat1_1_mcs_out[11]}), .b ({new_AGEMA_signal_9130, mcs1_mcs_mat1_1_mcs_out[15]}), .c ({new_AGEMA_signal_9399, mcs1_mcs_mat1_1_n116}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U75 ( .a ({new_AGEMA_signal_10338, mcs1_mcs_mat1_1_n114}), .b ({new_AGEMA_signal_9400, mcs1_mcs_mat1_1_n113}), .c ({new_AGEMA_signal_10629, mcs_out[251]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U74 ( .a ({new_AGEMA_signal_9104, mcs1_mcs_mat1_1_mcs_out[123]}), .b ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_9400, mcs1_mcs_mat1_1_n113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U73 ( .a ({new_AGEMA_signal_10106, mcs1_mcs_mat1_1_mcs_out[115]}), .b ({new_AGEMA_signal_9106, mcs1_mcs_mat1_1_mcs_out[119]}), .c ({new_AGEMA_signal_10338, mcs1_mcs_mat1_1_n114}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U72 ( .a ({new_AGEMA_signal_10095, mcs1_mcs_mat1_1_n112}), .b ({new_AGEMA_signal_8162, mcs1_mcs_mat1_1_n111}), .c ({new_AGEMA_signal_10339, mcs_out[250]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U71 ( .a ({new_AGEMA_signal_7684, mcs1_mcs_mat1_1_mcs_out[122]}), .b ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_8162, mcs1_mcs_mat1_1_n111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U70 ( .a ({new_AGEMA_signal_9887, mcs1_mcs_mat1_1_mcs_out[114]}), .b ({new_AGEMA_signal_9107, mcs1_mcs_mat1_1_mcs_out[118]}), .c ({new_AGEMA_signal_10095, mcs1_mcs_mat1_1_n112}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U69 ( .a ({new_AGEMA_signal_9094, mcs1_mcs_mat1_1_n110}), .b ({new_AGEMA_signal_10096, mcs1_mcs_mat1_1_n109}), .c ({temp_next_s1[26], temp_next_s0[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U68 ( .a ({new_AGEMA_signal_9903, mcs1_mcs_mat1_1_mcs_out[2]}), .b ({new_AGEMA_signal_8218, mcs1_mcs_mat1_1_mcs_out[6]}), .c ({new_AGEMA_signal_10096, mcs1_mcs_mat1_1_n109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U67 ( .a ({new_AGEMA_signal_8696, mcs1_mcs_mat1_1_mcs_out[10]}), .b ({new_AGEMA_signal_8693, mcs1_mcs_mat1_1_mcs_out[14]}), .c ({new_AGEMA_signal_9094, mcs1_mcs_mat1_1_n110}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U66 ( .a ({new_AGEMA_signal_9882, mcs1_mcs_mat1_1_n108}), .b ({new_AGEMA_signal_9401, mcs1_mcs_mat1_1_n107}), .c ({new_AGEMA_signal_10097, mcs_out[249]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U65 ( .a ({new_AGEMA_signal_9105, mcs1_mcs_mat1_1_mcs_out[121]}), .b ({new_AGEMA_signal_7350, mcs1_mcs_mat1_1_mcs_out[125]}), .c ({new_AGEMA_signal_9401, mcs1_mcs_mat1_1_n107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U64 ( .a ({new_AGEMA_signal_9649, mcs1_mcs_mat1_1_mcs_out[113]}), .b ({new_AGEMA_signal_8649, mcs1_mcs_mat1_1_mcs_out[117]}), .c ({new_AGEMA_signal_9882, mcs1_mcs_mat1_1_n108}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U63 ( .a ({new_AGEMA_signal_10630, mcs1_mcs_mat1_1_n106}), .b ({new_AGEMA_signal_9095, mcs1_mcs_mat1_1_n105}), .c ({new_AGEMA_signal_10878, mcs_out[248]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U62 ( .a ({new_AGEMA_signal_8646, mcs1_mcs_mat1_1_mcs_out[120]}), .b ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_9095, mcs1_mcs_mat1_1_n105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U61 ( .a ({new_AGEMA_signal_10352, mcs1_mcs_mat1_1_mcs_out[112]}), .b ({new_AGEMA_signal_8168, mcs1_mcs_mat1_1_mcs_out[116]}), .c ({new_AGEMA_signal_10630, mcs1_mcs_mat1_1_n106}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U60 ( .a ({new_AGEMA_signal_9096, mcs1_mcs_mat1_1_n104}), .b ({new_AGEMA_signal_10631, mcs1_mcs_mat1_1_n103}), .c ({new_AGEMA_signal_10879, mcs_out[219]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U59 ( .a ({new_AGEMA_signal_9108, mcs1_mcs_mat1_1_mcs_out[111]}), .b ({new_AGEMA_signal_10353, mcs1_mcs_mat1_1_mcs_out[99]}), .c ({new_AGEMA_signal_10631, mcs1_mcs_mat1_1_n103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U58 ( .a ({new_AGEMA_signal_8658, mcs1_mcs_mat1_1_mcs_out[103]}), .b ({new_AGEMA_signal_8654, mcs1_mcs_mat1_1_mcs_out[107]}), .c ({new_AGEMA_signal_9096, mcs1_mcs_mat1_1_n104}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U57 ( .a ({new_AGEMA_signal_9097, mcs1_mcs_mat1_1_n102}), .b ({new_AGEMA_signal_10098, mcs1_mcs_mat1_1_n101}), .c ({new_AGEMA_signal_10341, mcs_out[218]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U56 ( .a ({new_AGEMA_signal_9109, mcs1_mcs_mat1_1_mcs_out[110]}), .b ({new_AGEMA_signal_9890, mcs1_mcs_mat1_1_mcs_out[98]}), .c ({new_AGEMA_signal_10098, mcs1_mcs_mat1_1_n101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U55 ( .a ({new_AGEMA_signal_7693, mcs1_mcs_mat1_1_mcs_out[102]}), .b ({new_AGEMA_signal_8655, mcs1_mcs_mat1_1_mcs_out[106]}), .c ({new_AGEMA_signal_9097, mcs1_mcs_mat1_1_n102}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U54 ( .a ({new_AGEMA_signal_9098, mcs1_mcs_mat1_1_n100}), .b ({new_AGEMA_signal_9646, mcs1_mcs_mat1_1_n99}), .c ({new_AGEMA_signal_9883, mcs_out[217]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U53 ( .a ({new_AGEMA_signal_9110, mcs1_mcs_mat1_1_mcs_out[109]}), .b ({new_AGEMA_signal_9411, mcs1_mcs_mat1_1_mcs_out[97]}), .c ({new_AGEMA_signal_9646, mcs1_mcs_mat1_1_n99}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U52 ( .a ({new_AGEMA_signal_8175, mcs1_mcs_mat1_1_mcs_out[101]}), .b ({new_AGEMA_signal_8656, mcs1_mcs_mat1_1_mcs_out[105]}), .c ({new_AGEMA_signal_9098, mcs1_mcs_mat1_1_n100}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U51 ( .a ({new_AGEMA_signal_9402, mcs1_mcs_mat1_1_n98}), .b ({new_AGEMA_signal_11047, mcs1_mcs_mat1_1_n97}), .c ({new_AGEMA_signal_11098, mcs_out[216]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U50 ( .a ({new_AGEMA_signal_9111, mcs1_mcs_mat1_1_mcs_out[108]}), .b ({new_AGEMA_signal_10882, mcs1_mcs_mat1_1_mcs_out[96]}), .c ({new_AGEMA_signal_11047, mcs1_mcs_mat1_1_n97}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U49 ( .a ({new_AGEMA_signal_8659, mcs1_mcs_mat1_1_mcs_out[100]}), .b ({new_AGEMA_signal_9112, mcs1_mcs_mat1_1_mcs_out[104]}), .c ({new_AGEMA_signal_9402, mcs1_mcs_mat1_1_n98}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U48 ( .a ({new_AGEMA_signal_10099, mcs1_mcs_mat1_1_n96}), .b ({new_AGEMA_signal_9099, mcs1_mcs_mat1_1_n95}), .c ({new_AGEMA_signal_10342, mcs_out[187]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U47 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_8662, mcs1_mcs_mat1_1_mcs_out[95]}), .c ({new_AGEMA_signal_9099, mcs1_mcs_mat1_1_n95}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U46 ( .a ({new_AGEMA_signal_9891, mcs1_mcs_mat1_1_mcs_out[83]}), .b ({new_AGEMA_signal_7700, mcs1_mcs_mat1_1_mcs_out[87]}), .c ({new_AGEMA_signal_10099, mcs1_mcs_mat1_1_n96}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U45 ( .a ({new_AGEMA_signal_10100, mcs1_mcs_mat1_1_n94}), .b ({new_AGEMA_signal_8163, mcs1_mcs_mat1_1_n93}), .c ({new_AGEMA_signal_10343, mcs_out[186]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U43 ( .a ({new_AGEMA_signal_9892, mcs1_mcs_mat1_1_mcs_out[82]}), .b ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_10100, mcs1_mcs_mat1_1_n94}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U42 ( .a ({new_AGEMA_signal_10101, mcs1_mcs_mat1_1_n92}), .b ({new_AGEMA_signal_8164, mcs1_mcs_mat1_1_n91}), .c ({new_AGEMA_signal_10344, mcs_out[185]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U41 ( .a ({new_AGEMA_signal_7365, mcs1_mcs_mat1_1_mcs_out[89]}), .b ({new_AGEMA_signal_7698, mcs1_mcs_mat1_1_mcs_out[93]}), .c ({new_AGEMA_signal_8164, mcs1_mcs_mat1_1_n91}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U40 ( .a ({new_AGEMA_signal_9893, mcs1_mcs_mat1_1_mcs_out[81]}), .b ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_10101, mcs1_mcs_mat1_1_n92}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U39 ( .a ({new_AGEMA_signal_10345, mcs1_mcs_mat1_1_n90}), .b ({new_AGEMA_signal_9403, mcs1_mcs_mat1_1_n89}), .c ({new_AGEMA_signal_10632, mcs_out[184]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U38 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_9113, mcs1_mcs_mat1_1_mcs_out[92]}), .c ({new_AGEMA_signal_9403, mcs1_mcs_mat1_1_n89}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U37 ( .a ({new_AGEMA_signal_10109, mcs1_mcs_mat1_1_mcs_out[80]}), .b ({new_AGEMA_signal_8179, mcs1_mcs_mat1_1_mcs_out[84]}), .c ({new_AGEMA_signal_10345, mcs1_mcs_mat1_1_n90}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U36 ( .a ({new_AGEMA_signal_10346, mcs1_mcs_mat1_1_n88}), .b ({new_AGEMA_signal_8640, mcs1_mcs_mat1_1_n87}), .c ({temp_next_s1[25], temp_next_s0[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U35 ( .a ({new_AGEMA_signal_7386, mcs1_mcs_mat1_1_mcs_out[5]}), .b ({new_AGEMA_signal_8216, mcs1_mcs_mat1_1_mcs_out[9]}), .c ({new_AGEMA_signal_8640, mcs1_mcs_mat1_1_n87}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U34 ( .a ({new_AGEMA_signal_8694, mcs1_mcs_mat1_1_mcs_out[13]}), .b ({new_AGEMA_signal_10115, mcs1_mcs_mat1_1_mcs_out[1]}), .c ({new_AGEMA_signal_10346, mcs1_mcs_mat1_1_n88}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U33 ( .a ({new_AGEMA_signal_10634, mcs1_mcs_mat1_1_n86}), .b ({new_AGEMA_signal_9100, mcs1_mcs_mat1_1_n85}), .c ({new_AGEMA_signal_10880, mcs_out[155]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U32 ( .a ({new_AGEMA_signal_7703, mcs1_mcs_mat1_1_mcs_out[75]}), .b ({new_AGEMA_signal_8665, mcs1_mcs_mat1_1_mcs_out[79]}), .c ({new_AGEMA_signal_9100, mcs1_mcs_mat1_1_n85}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U31 ( .a ({new_AGEMA_signal_10354, mcs1_mcs_mat1_1_mcs_out[67]}), .b ({new_AGEMA_signal_8669, mcs1_mcs_mat1_1_mcs_out[71]}), .c ({new_AGEMA_signal_10634, mcs1_mcs_mat1_1_n86}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U30 ( .a ({new_AGEMA_signal_10347, mcs1_mcs_mat1_1_n84}), .b ({new_AGEMA_signal_9404, mcs1_mcs_mat1_1_n83}), .c ({new_AGEMA_signal_10635, mcs_out[154]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U29 ( .a ({new_AGEMA_signal_9115, mcs1_mcs_mat1_1_mcs_out[74]}), .b ({new_AGEMA_signal_6987, mcs1_mcs_mat1_1_mcs_out[78]}), .c ({new_AGEMA_signal_9404, mcs1_mcs_mat1_1_n83}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U28 ( .a ({new_AGEMA_signal_10110, mcs1_mcs_mat1_1_mcs_out[66]}), .b ({new_AGEMA_signal_9117, mcs1_mcs_mat1_1_mcs_out[70]}), .c ({new_AGEMA_signal_10347, mcs1_mcs_mat1_1_n84}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U27 ( .a ({new_AGEMA_signal_9884, mcs1_mcs_mat1_1_n82}), .b ({new_AGEMA_signal_8641, mcs1_mcs_mat1_1_n81}), .c ({new_AGEMA_signal_10102, mcs_out[153]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U26 ( .a ({new_AGEMA_signal_8182, mcs1_mcs_mat1_1_mcs_out[73]}), .b ({new_AGEMA_signal_7701, mcs1_mcs_mat1_1_mcs_out[77]}), .c ({new_AGEMA_signal_8641, mcs1_mcs_mat1_1_n81}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U25 ( .a ({new_AGEMA_signal_9657, mcs1_mcs_mat1_1_mcs_out[65]}), .b ({new_AGEMA_signal_9118, mcs1_mcs_mat1_1_mcs_out[69]}), .c ({new_AGEMA_signal_9884, mcs1_mcs_mat1_1_n82}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U24 ( .a ({new_AGEMA_signal_10881, mcs1_mcs_mat1_1_n80}), .b ({new_AGEMA_signal_9405, mcs1_mcs_mat1_1_n79}), .c ({new_AGEMA_signal_11048, mcs_out[152]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U23 ( .a ({new_AGEMA_signal_9116, mcs1_mcs_mat1_1_mcs_out[72]}), .b ({new_AGEMA_signal_9114, mcs1_mcs_mat1_1_mcs_out[76]}), .c ({new_AGEMA_signal_9405, mcs1_mcs_mat1_1_n79}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U22 ( .a ({new_AGEMA_signal_10639, mcs1_mcs_mat1_1_mcs_out[64]}), .b ({new_AGEMA_signal_8671, mcs1_mcs_mat1_1_mcs_out[68]}), .c ({new_AGEMA_signal_10881, mcs1_mcs_mat1_1_n80}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U21 ( .a ({new_AGEMA_signal_9885, mcs1_mcs_mat1_1_n78}), .b ({new_AGEMA_signal_9101, mcs1_mcs_mat1_1_n77}), .c ({temp_next_s1[123], temp_next_s0[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U20 ( .a ({new_AGEMA_signal_8190, mcs1_mcs_mat1_1_mcs_out[59]}), .b ({new_AGEMA_signal_8673, mcs1_mcs_mat1_1_mcs_out[63]}), .c ({new_AGEMA_signal_9101, mcs1_mcs_mat1_1_n77}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U19 ( .a ({new_AGEMA_signal_9659, mcs1_mcs_mat1_1_mcs_out[51]}), .b ({new_AGEMA_signal_8676, mcs1_mcs_mat1_1_mcs_out[55]}), .c ({new_AGEMA_signal_9885, mcs1_mcs_mat1_1_n78}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U18 ( .a ({new_AGEMA_signal_9406, mcs1_mcs_mat1_1_n76}), .b ({new_AGEMA_signal_8642, mcs1_mcs_mat1_1_n75}), .c ({temp_next_s1[122], temp_next_s0[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U17 ( .a ({new_AGEMA_signal_7711, mcs1_mcs_mat1_1_mcs_out[58]}), .b ({new_AGEMA_signal_8187, mcs1_mcs_mat1_1_mcs_out[62]}), .c ({new_AGEMA_signal_8642, mcs1_mcs_mat1_1_n75}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U16 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_9120, mcs1_mcs_mat1_1_mcs_out[54]}), .c ({new_AGEMA_signal_9406, mcs1_mcs_mat1_1_n76}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U15 ( .a ({new_AGEMA_signal_9407, mcs1_mcs_mat1_1_n74}), .b ({new_AGEMA_signal_8643, mcs1_mcs_mat1_1_n73}), .c ({temp_next_s1[121], temp_next_s0[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U14 ( .a ({new_AGEMA_signal_8191, mcs1_mcs_mat1_1_mcs_out[57]}), .b ({new_AGEMA_signal_8188, mcs1_mcs_mat1_1_mcs_out[61]}), .c ({new_AGEMA_signal_8643, mcs1_mcs_mat1_1_n73}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U13 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_9121, mcs1_mcs_mat1_1_mcs_out[53]}), .c ({new_AGEMA_signal_9407, mcs1_mcs_mat1_1_n74}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U12 ( .a ({new_AGEMA_signal_10104, mcs1_mcs_mat1_1_n72}), .b ({new_AGEMA_signal_9408, mcs1_mcs_mat1_1_n71}), .c ({temp_next_s1[120], temp_next_s0[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U11 ( .a ({new_AGEMA_signal_8675, mcs1_mcs_mat1_1_mcs_out[56]}), .b ({new_AGEMA_signal_9119, mcs1_mcs_mat1_1_mcs_out[60]}), .c ({new_AGEMA_signal_9408, mcs1_mcs_mat1_1_n71}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U10 ( .a ({new_AGEMA_signal_9896, mcs1_mcs_mat1_1_mcs_out[48]}), .b ({new_AGEMA_signal_8678, mcs1_mcs_mat1_1_mcs_out[52]}), .c ({new_AGEMA_signal_10104, mcs1_mcs_mat1_1_n72}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U9 ( .a ({new_AGEMA_signal_10349, mcs1_mcs_mat1_1_n70}), .b ({new_AGEMA_signal_9102, mcs1_mcs_mat1_1_n69}), .c ({temp_next_s1[91], temp_next_s0[91]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U8 ( .a ({new_AGEMA_signal_8680, mcs1_mcs_mat1_1_mcs_out[43]}), .b ({new_AGEMA_signal_8679, mcs1_mcs_mat1_1_mcs_out[47]}), .c ({new_AGEMA_signal_9102, mcs1_mcs_mat1_1_n69}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U7 ( .a ({new_AGEMA_signal_10112, mcs1_mcs_mat1_1_mcs_out[35]}), .b ({new_AGEMA_signal_9123, mcs1_mcs_mat1_1_mcs_out[39]}), .c ({new_AGEMA_signal_10349, mcs1_mcs_mat1_1_n70}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U6 ( .a ({new_AGEMA_signal_10105, mcs1_mcs_mat1_1_n68}), .b ({new_AGEMA_signal_9103, mcs1_mcs_mat1_1_n67}), .c ({temp_next_s1[90], temp_next_s0[90]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U5 ( .a ({new_AGEMA_signal_8681, mcs1_mcs_mat1_1_mcs_out[42]}), .b ({new_AGEMA_signal_7373, mcs1_mcs_mat1_1_mcs_out[46]}), .c ({new_AGEMA_signal_9103, mcs1_mcs_mat1_1_n67}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U4 ( .a ({new_AGEMA_signal_9897, mcs1_mcs_mat1_1_mcs_out[34]}), .b ({new_AGEMA_signal_7724, mcs1_mcs_mat1_1_mcs_out[38]}), .c ({new_AGEMA_signal_10105, mcs1_mcs_mat1_1_n68}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U3 ( .a ({new_AGEMA_signal_10351, mcs1_mcs_mat1_1_n66}), .b ({new_AGEMA_signal_9886, mcs1_mcs_mat1_1_n65}), .c ({temp_next_s1[24], temp_next_s0[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U2 ( .a ({new_AGEMA_signal_9666, mcs1_mcs_mat1_1_mcs_out[4]}), .b ({new_AGEMA_signal_9132, mcs1_mcs_mat1_1_mcs_out[8]}), .c ({new_AGEMA_signal_9886, mcs1_mcs_mat1_1_n65}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_U1 ( .a ({new_AGEMA_signal_10116, mcs1_mcs_mat1_1_mcs_out[0]}), .b ({new_AGEMA_signal_9419, mcs1_mcs_mat1_1_mcs_out[12]}), .c ({new_AGEMA_signal_10351, mcs1_mcs_mat1_1_n66}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_8644, mcs1_mcs_mat1_1_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_9104, mcs1_mcs_mat1_1_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_8165, mcs1_mcs_mat1_1_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_6721, mcs1_mcs_mat1_1_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8644, mcs1_mcs_mat1_1_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_6980, mcs1_mcs_mat1_1_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_7351, mcs1_mcs_mat1_1_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_7684, mcs1_mcs_mat1_1_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_6981, mcs1_mcs_mat1_1_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_7232, shiftr_out[91]}), .c ({new_AGEMA_signal_7351, mcs1_mcs_mat1_1_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_8645, mcs1_mcs_mat1_1_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_7232, shiftr_out[91]}), .c ({new_AGEMA_signal_9105, mcs1_mcs_mat1_1_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_8165, mcs1_mcs_mat1_1_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_8645, mcs1_mcs_mat1_1_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_7685, mcs1_mcs_mat1_1_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_7352, mcs1_mcs_mat1_1_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_8165, mcs1_mcs_mat1_1_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_8166, mcs1_mcs_mat1_1_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_8646, mcs1_mcs_mat1_1_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_7685, mcs1_mcs_mat1_1_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_6981, mcs1_mcs_mat1_1_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_8166, mcs1_mcs_mat1_1_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[532]), .c ({new_AGEMA_signal_7685, mcs1_mcs_mat1_1_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[533]), .c ({new_AGEMA_signal_6981, mcs1_mcs_mat1_1_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7232, shiftr_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[534]), .c ({new_AGEMA_signal_7352, mcs1_mcs_mat1_1_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_8647, mcs1_mcs_mat1_1_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_6692, shiftr_out[58]}), .c ({new_AGEMA_signal_9106, mcs1_mcs_mat1_1_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_8167, mcs1_mcs_mat1_1_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7355, mcs1_mcs_mat1_1_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_8647, mcs1_mcs_mat1_1_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_8648, mcs1_mcs_mat1_1_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_7687, mcs1_mcs_mat1_1_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_9107, mcs1_mcs_mat1_1_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_8167, mcs1_mcs_mat1_1_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7304, shiftr_out[57]}), .c ({new_AGEMA_signal_8648, mcs1_mcs_mat1_1_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_8167, mcs1_mcs_mat1_1_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7686, mcs1_mcs_mat1_1_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_8649, mcs1_mcs_mat1_1_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_7688, mcs1_mcs_mat1_1_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_6982, mcs1_mcs_mat1_1_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_8167, mcs1_mcs_mat1_1_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_7354, mcs1_mcs_mat1_1_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_7687, mcs1_mcs_mat1_1_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_8168, mcs1_mcs_mat1_1_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_6722, mcs1_mcs_mat1_1_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7355, mcs1_mcs_mat1_1_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_7687, mcs1_mcs_mat1_1_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_6982, mcs1_mcs_mat1_1_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_7354, mcs1_mcs_mat1_1_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7304, shiftr_out[57]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[535]), .c ({new_AGEMA_signal_7688, mcs1_mcs_mat1_1_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[536]), .c ({new_AGEMA_signal_6982, mcs1_mcs_mat1_1_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[537]), .c ({new_AGEMA_signal_7355, mcs1_mcs_mat1_1_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_9888, mcs1_mcs_mat1_1_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_8650, mcs1_mcs_mat1_1_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_10106, mcs1_mcs_mat1_1_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_9409, mcs1_mcs_mat1_1_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_9410, mcs1_mcs_mat1_1_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_9649, mcs1_mcs_mat1_1_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_9889, mcs1_mcs_mat1_1_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_10107, mcs1_mcs_mat1_1_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_10352, mcs1_mcs_mat1_1_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_9888, mcs1_mcs_mat1_1_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_10107, mcs1_mcs_mat1_1_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_8169, mcs1_mcs_mat1_1_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9651, mcs1_mcs_mat1_1_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_9888, mcs1_mcs_mat1_1_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_8651, mcs1_mcs_mat1_1_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_9650, mcs1_mcs_mat1_1_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_9889, mcs1_mcs_mat1_1_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9363, shiftr_out[25]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[538]), .c ({new_AGEMA_signal_9651, mcs1_mcs_mat1_1_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[539]), .c ({new_AGEMA_signal_8651, mcs1_mcs_mat1_1_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[540]), .c ({new_AGEMA_signal_9410, mcs1_mcs_mat1_1_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({new_AGEMA_signal_8652, mcs1_mcs_mat1_1_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9108, mcs1_mcs_mat1_1_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({new_AGEMA_signal_8653, mcs1_mcs_mat1_1_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9109, mcs1_mcs_mat1_1_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_7356, mcs1_mcs_mat1_1_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_8652, mcs1_mcs_mat1_1_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9110, mcs1_mcs_mat1_1_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_6983, mcs1_mcs_mat1_1_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_8170, mcs1_mcs_mat1_1_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_8652, mcs1_mcs_mat1_1_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_7689, mcs1_mcs_mat1_1_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8653, mcs1_mcs_mat1_1_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9111, mcs1_mcs_mat1_1_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_8171, mcs1_mcs_mat1_1_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_8653, mcs1_mcs_mat1_1_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_7356, mcs1_mcs_mat1_1_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_7690, mcs1_mcs_mat1_1_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_8171, mcs1_mcs_mat1_1_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[541]), .c ({new_AGEMA_signal_7690, mcs1_mcs_mat1_1_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[542]), .c ({new_AGEMA_signal_6983, mcs1_mcs_mat1_1_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[543]), .c ({new_AGEMA_signal_7356, mcs1_mcs_mat1_1_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_8173, mcs1_mcs_mat1_1_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_8172, mcs1_mcs_mat1_1_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8654, mcs1_mcs_mat1_1_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_8172, mcs1_mcs_mat1_1_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_7357, mcs1_mcs_mat1_1_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_8655, mcs1_mcs_mat1_1_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_6984, mcs1_mcs_mat1_1_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7232, shiftr_out[91]}), .c ({new_AGEMA_signal_7357, mcs1_mcs_mat1_1_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_8172, mcs1_mcs_mat1_1_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8656, mcs1_mcs_mat1_1_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_7692, mcs1_mcs_mat1_1_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_6724, mcs1_mcs_mat1_1_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_8172, mcs1_mcs_mat1_1_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_8657, mcs1_mcs_mat1_1_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_9112, mcs1_mcs_mat1_1_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_8173, mcs1_mcs_mat1_1_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_7692, mcs1_mcs_mat1_1_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_8657, mcs1_mcs_mat1_1_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_7691, mcs1_mcs_mat1_1_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_6618, shiftr_out[88]}), .c ({new_AGEMA_signal_8173, mcs1_mcs_mat1_1_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_6984, mcs1_mcs_mat1_1_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7358, mcs1_mcs_mat1_1_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_7691, mcs1_mcs_mat1_1_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[544]), .c ({new_AGEMA_signal_7692, mcs1_mcs_mat1_1_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[545]), .c ({new_AGEMA_signal_6984, mcs1_mcs_mat1_1_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7232, shiftr_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[546]), .c ({new_AGEMA_signal_7358, mcs1_mcs_mat1_1_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_7359, mcs1_mcs_mat1_1_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_8174, mcs1_mcs_mat1_1_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_8658, mcs1_mcs_mat1_1_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_7696, mcs1_mcs_mat1_1_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_8174, mcs1_mcs_mat1_1_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_7694, mcs1_mcs_mat1_1_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_7360, mcs1_mcs_mat1_1_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_8175, mcs1_mcs_mat1_1_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_7695, mcs1_mcs_mat1_1_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_8176, mcs1_mcs_mat1_1_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_8659, mcs1_mcs_mat1_1_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_6725, mcs1_mcs_mat1_1_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7696, mcs1_mcs_mat1_1_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_8176, mcs1_mcs_mat1_1_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_6985, mcs1_mcs_mat1_1_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_7304, shiftr_out[57]}), .c ({new_AGEMA_signal_7695, mcs1_mcs_mat1_1_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7304, shiftr_out[57]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[547]), .c ({new_AGEMA_signal_7696, mcs1_mcs_mat1_1_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[548]), .c ({new_AGEMA_signal_6985, mcs1_mcs_mat1_1_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[549]), .c ({new_AGEMA_signal_7360, mcs1_mcs_mat1_1_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_10638, mcs1_mcs_mat1_1_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_9412, mcs1_mcs_mat1_1_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_10882, mcs1_mcs_mat1_1_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_10353, mcs1_mcs_mat1_1_mcs_out[99]}), .b ({new_AGEMA_signal_8101, shiftr_out[26]}), .c ({new_AGEMA_signal_10638, mcs1_mcs_mat1_1_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_10108, mcs1_mcs_mat1_1_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_9363, shiftr_out[25]}), .c ({new_AGEMA_signal_10353, mcs1_mcs_mat1_1_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_9890, mcs1_mcs_mat1_1_mcs_out[98]}), .b ({new_AGEMA_signal_8661, mcs1_mcs_mat1_1_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_10108, mcs1_mcs_mat1_1_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_8660, mcs1_mcs_mat1_1_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_9652, mcs1_mcs_mat1_1_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_9890, mcs1_mcs_mat1_1_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9363, shiftr_out[25]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[550]), .c ({new_AGEMA_signal_9652, mcs1_mcs_mat1_1_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[551]), .c ({new_AGEMA_signal_8661, mcs1_mcs_mat1_1_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[552]), .c ({new_AGEMA_signal_9412, mcs1_mcs_mat1_1_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_8178, mcs1_mcs_mat1_1_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_8662, mcs1_mcs_mat1_1_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_7362, mcs1_mcs_mat1_1_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_7363, mcs1_mcs_mat1_1_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_7698, mcs1_mcs_mat1_1_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_8663, mcs1_mcs_mat1_1_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_6986, mcs1_mcs_mat1_1_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_9113, mcs1_mcs_mat1_1_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_8178, mcs1_mcs_mat1_1_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_8663, mcs1_mcs_mat1_1_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_6726, mcs1_mcs_mat1_1_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7699, mcs1_mcs_mat1_1_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_8178, mcs1_mcs_mat1_1_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[553]), .c ({new_AGEMA_signal_7699, mcs1_mcs_mat1_1_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[554]), .c ({new_AGEMA_signal_6986, mcs1_mcs_mat1_1_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[555]), .c ({new_AGEMA_signal_7363, mcs1_mcs_mat1_1_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_9655, mcs1_mcs_mat1_1_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_9656, mcs1_mcs_mat1_1_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_9891, mcs1_mcs_mat1_1_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_9653, mcs1_mcs_mat1_1_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_8180, mcs1_mcs_mat1_1_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_9892, mcs1_mcs_mat1_1_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_9413, mcs1_mcs_mat1_1_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_9653, mcs1_mcs_mat1_1_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_9654, mcs1_mcs_mat1_1_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_9893, mcs1_mcs_mat1_1_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_8664, mcs1_mcs_mat1_1_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_9413, mcs1_mcs_mat1_1_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_9654, mcs1_mcs_mat1_1_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_9894, mcs1_mcs_mat1_1_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_8101, shiftr_out[26]}), .c ({new_AGEMA_signal_10109, mcs1_mcs_mat1_1_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_9655, mcs1_mcs_mat1_1_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_8664, mcs1_mcs_mat1_1_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_9894, mcs1_mcs_mat1_1_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9363, shiftr_out[25]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[556]), .c ({new_AGEMA_signal_9656, mcs1_mcs_mat1_1_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[557]), .c ({new_AGEMA_signal_8664, mcs1_mcs_mat1_1_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[558]), .c ({new_AGEMA_signal_9413, mcs1_mcs_mat1_1_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_8181, mcs1_mcs_mat1_1_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_8665, mcs1_mcs_mat1_1_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_7366, mcs1_mcs_mat1_1_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_7701, mcs1_mcs_mat1_1_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_8666, mcs1_mcs_mat1_1_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_6988, mcs1_mcs_mat1_1_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_9114, mcs1_mcs_mat1_1_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_8181, mcs1_mcs_mat1_1_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_6613, shiftr_out[120]}), .c ({new_AGEMA_signal_8666, mcs1_mcs_mat1_1_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_6727, mcs1_mcs_mat1_1_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7702, mcs1_mcs_mat1_1_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_8181, mcs1_mcs_mat1_1_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[559]), .c ({new_AGEMA_signal_7702, mcs1_mcs_mat1_1_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[560]), .c ({new_AGEMA_signal_6988, mcs1_mcs_mat1_1_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[561]), .c ({new_AGEMA_signal_7366, mcs1_mcs_mat1_1_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_8667, mcs1_mcs_mat1_1_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_9115, mcs1_mcs_mat1_1_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_8183, mcs1_mcs_mat1_1_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7704, mcs1_mcs_mat1_1_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_8667, mcs1_mcs_mat1_1_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_7250, mcs1_mcs_mat1_1_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_7703, mcs1_mcs_mat1_1_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_7704, mcs1_mcs_mat1_1_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_7250, mcs1_mcs_mat1_1_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_8182, mcs1_mcs_mat1_1_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_6989, mcs1_mcs_mat1_1_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_6990, mcs1_mcs_mat1_1_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_7250, mcs1_mcs_mat1_1_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_7367, mcs1_mcs_mat1_1_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_6618, shiftr_out[88]}), .c ({new_AGEMA_signal_7704, mcs1_mcs_mat1_1_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_8668, mcs1_mcs_mat1_1_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_6989, mcs1_mcs_mat1_1_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_9116, mcs1_mcs_mat1_1_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_8183, mcs1_mcs_mat1_1_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7367, mcs1_mcs_mat1_1_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_8668, mcs1_mcs_mat1_1_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_7232, shiftr_out[91]}), .b ({new_AGEMA_signal_7705, mcs1_mcs_mat1_1_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_8183, mcs1_mcs_mat1_1_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[562]), .c ({new_AGEMA_signal_7705, mcs1_mcs_mat1_1_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[563]), .c ({new_AGEMA_signal_6990, mcs1_mcs_mat1_1_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7232, shiftr_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[564]), .c ({new_AGEMA_signal_7367, mcs1_mcs_mat1_1_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_8184, mcs1_mcs_mat1_1_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_7368, mcs1_mcs_mat1_1_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_8669, mcs1_mcs_mat1_1_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_7707, mcs1_mcs_mat1_1_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_8670, mcs1_mcs_mat1_1_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9117, mcs1_mcs_mat1_1_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_8184, mcs1_mcs_mat1_1_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_8670, mcs1_mcs_mat1_1_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9118, mcs1_mcs_mat1_1_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_7368, mcs1_mcs_mat1_1_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_8185, mcs1_mcs_mat1_1_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_8670, mcs1_mcs_mat1_1_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({new_AGEMA_signal_6991, mcs1_mcs_mat1_1_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_7368, mcs1_mcs_mat1_1_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_7706, mcs1_mcs_mat1_1_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_7304, shiftr_out[57]}), .c ({new_AGEMA_signal_8184, mcs1_mcs_mat1_1_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_7369, mcs1_mcs_mat1_1_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6729, mcs1_mcs_mat1_1_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_7706, mcs1_mcs_mat1_1_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_8185, mcs1_mcs_mat1_1_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_7707, mcs1_mcs_mat1_1_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_8671, mcs1_mcs_mat1_1_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_7369, mcs1_mcs_mat1_1_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_7707, mcs1_mcs_mat1_1_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({new_AGEMA_signal_7708, mcs1_mcs_mat1_1_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_8185, mcs1_mcs_mat1_1_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7304, shiftr_out[57]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[565]), .c ({new_AGEMA_signal_7708, mcs1_mcs_mat1_1_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[566]), .c ({new_AGEMA_signal_6991, mcs1_mcs_mat1_1_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[567]), .c ({new_AGEMA_signal_7369, mcs1_mcs_mat1_1_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_10111, mcs1_mcs_mat1_1_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_10354, mcs1_mcs_mat1_1_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({new_AGEMA_signal_9895, mcs1_mcs_mat1_1_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_10110, mcs1_mcs_mat1_1_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_10355, mcs1_mcs_mat1_1_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_9414, mcs1_mcs_mat1_1_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_10639, mcs1_mcs_mat1_1_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_10111, mcs1_mcs_mat1_1_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .c ({new_AGEMA_signal_10355, mcs1_mcs_mat1_1_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_8672, mcs1_mcs_mat1_1_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_9895, mcs1_mcs_mat1_1_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_10111, mcs1_mcs_mat1_1_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_8186, mcs1_mcs_mat1_1_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_9658, mcs1_mcs_mat1_1_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_9895, mcs1_mcs_mat1_1_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9363, shiftr_out[25]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[568]), .c ({new_AGEMA_signal_9658, mcs1_mcs_mat1_1_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[569]), .c ({new_AGEMA_signal_8672, mcs1_mcs_mat1_1_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[570]), .c ({new_AGEMA_signal_9414, mcs1_mcs_mat1_1_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_8189, mcs1_mcs_mat1_1_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7370, mcs1_mcs_mat1_1_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_8673, mcs1_mcs_mat1_1_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_6992, mcs1_mcs_mat1_1_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_7709, mcs1_mcs_mat1_1_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8187, mcs1_mcs_mat1_1_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({new_AGEMA_signal_7710, mcs1_mcs_mat1_1_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_8188, mcs1_mcs_mat1_1_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[571]), .c ({new_AGEMA_signal_7710, mcs1_mcs_mat1_1_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[572]), .c ({new_AGEMA_signal_6992, mcs1_mcs_mat1_1_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[573]), .c ({new_AGEMA_signal_7370, mcs1_mcs_mat1_1_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_6994, mcs1_mcs_mat1_1_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_7371, mcs1_mcs_mat1_1_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_7711, mcs1_mcs_mat1_1_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_6995, mcs1_mcs_mat1_1_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_7712, mcs1_mcs_mat1_1_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_8191, mcs1_mcs_mat1_1_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_8192, mcs1_mcs_mat1_1_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_7713, mcs1_mcs_mat1_1_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_8675, mcs1_mcs_mat1_1_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_7714, mcs1_mcs_mat1_1_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_8192, mcs1_mcs_mat1_1_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[574]), .c ({new_AGEMA_signal_7714, mcs1_mcs_mat1_1_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[575]), .c ({new_AGEMA_signal_6995, mcs1_mcs_mat1_1_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7232, shiftr_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[576]), .c ({new_AGEMA_signal_7371, mcs1_mcs_mat1_1_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_7716, mcs1_mcs_mat1_1_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8193, mcs1_mcs_mat1_1_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_8676, mcs1_mcs_mat1_1_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_8677, mcs1_mcs_mat1_1_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_7715, mcs1_mcs_mat1_1_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_9120, mcs1_mcs_mat1_1_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_7372, mcs1_mcs_mat1_1_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_7715, mcs1_mcs_mat1_1_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({new_AGEMA_signal_8677, mcs1_mcs_mat1_1_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_9121, mcs1_mcs_mat1_1_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_6732, mcs1_mcs_mat1_1_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_8193, mcs1_mcs_mat1_1_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_8677, mcs1_mcs_mat1_1_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_6996, mcs1_mcs_mat1_1_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_7718, mcs1_mcs_mat1_1_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_8193, mcs1_mcs_mat1_1_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_7717, mcs1_mcs_mat1_1_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_8194, mcs1_mcs_mat1_1_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_8678, mcs1_mcs_mat1_1_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_7716, mcs1_mcs_mat1_1_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_6996, mcs1_mcs_mat1_1_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_8194, mcs1_mcs_mat1_1_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_7372, mcs1_mcs_mat1_1_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_7716, mcs1_mcs_mat1_1_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7304, shiftr_out[57]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[577]), .c ({new_AGEMA_signal_7718, mcs1_mcs_mat1_1_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[578]), .c ({new_AGEMA_signal_6996, mcs1_mcs_mat1_1_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[579]), .c ({new_AGEMA_signal_7372, mcs1_mcs_mat1_1_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_7374, mcs1_mcs_mat1_1_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_7719, mcs1_mcs_mat1_1_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_9122, mcs1_mcs_mat1_1_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_6997, mcs1_mcs_mat1_1_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_9415, mcs1_mcs_mat1_1_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_8679, mcs1_mcs_mat1_1_mcs_out[47]}), .b ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_9122, mcs1_mcs_mat1_1_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_8195, mcs1_mcs_mat1_1_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_6613, shiftr_out[120]}), .c ({new_AGEMA_signal_8679, mcs1_mcs_mat1_1_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_6733, mcs1_mcs_mat1_1_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_7720, mcs1_mcs_mat1_1_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_8195, mcs1_mcs_mat1_1_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[580]), .c ({new_AGEMA_signal_7720, mcs1_mcs_mat1_1_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[581]), .c ({new_AGEMA_signal_6997, mcs1_mcs_mat1_1_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[582]), .c ({new_AGEMA_signal_7374, mcs1_mcs_mat1_1_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_8196, mcs1_mcs_mat1_1_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_7375, mcs1_mcs_mat1_1_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_8680, mcs1_mcs_mat1_1_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_7721, mcs1_mcs_mat1_1_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_6998, mcs1_mcs_mat1_1_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_8196, mcs1_mcs_mat1_1_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_8197, mcs1_mcs_mat1_1_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_7723, mcs1_mcs_mat1_1_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_8681, mcs1_mcs_mat1_1_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_8198, mcs1_mcs_mat1_1_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_6734, mcs1_mcs_mat1_1_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_8682, mcs1_mcs_mat1_1_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_7721, mcs1_mcs_mat1_1_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7376, mcs1_mcs_mat1_1_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8198, mcs1_mcs_mat1_1_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_7722, mcs1_mcs_mat1_1_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_7376, mcs1_mcs_mat1_1_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8199, mcs1_mcs_mat1_1_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[583]), .c ({new_AGEMA_signal_7723, mcs1_mcs_mat1_1_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[584]), .c ({new_AGEMA_signal_6998, mcs1_mcs_mat1_1_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7232, shiftr_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[585]), .c ({new_AGEMA_signal_7376, mcs1_mcs_mat1_1_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_8683, mcs1_mcs_mat1_1_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_6735, mcs1_mcs_mat1_1_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9123, mcs1_mcs_mat1_1_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_7378, mcs1_mcs_mat1_1_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_7377, mcs1_mcs_mat1_1_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_7724, mcs1_mcs_mat1_1_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({new_AGEMA_signal_8683, mcs1_mcs_mat1_1_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_9124, mcs1_mcs_mat1_1_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_7725, mcs1_mcs_mat1_1_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_8200, mcs1_mcs_mat1_1_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_8683, mcs1_mcs_mat1_1_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_7726, mcs1_mcs_mat1_1_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7379, mcs1_mcs_mat1_1_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_8200, mcs1_mcs_mat1_1_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_7726, mcs1_mcs_mat1_1_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7378, mcs1_mcs_mat1_1_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_8201, mcs1_mcs_mat1_1_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_7251, mcs1_mcs_mat1_1_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_7378, mcs1_mcs_mat1_1_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({new_AGEMA_signal_6999, mcs1_mcs_mat1_1_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_7251, mcs1_mcs_mat1_1_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7304, shiftr_out[57]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[586]), .c ({new_AGEMA_signal_7726, mcs1_mcs_mat1_1_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[587]), .c ({new_AGEMA_signal_6999, mcs1_mcs_mat1_1_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[588]), .c ({new_AGEMA_signal_7379, mcs1_mcs_mat1_1_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_9660, mcs1_mcs_mat1_1_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_9416, mcs1_mcs_mat1_1_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_9897, mcs1_mcs_mat1_1_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_8684, mcs1_mcs_mat1_1_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_9125, mcs1_mcs_mat1_1_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_10356, mcs1_mcs_mat1_1_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_9661, mcs1_mcs_mat1_1_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_10640, mcs1_mcs_mat1_1_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9363, shiftr_out[25]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[589]), .c ({new_AGEMA_signal_9661, mcs1_mcs_mat1_1_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[590]), .c ({new_AGEMA_signal_8684, mcs1_mcs_mat1_1_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[591]), .c ({new_AGEMA_signal_9416, mcs1_mcs_mat1_1_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_8685, mcs1_mcs_mat1_1_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_8203, mcs1_mcs_mat1_1_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_9126, mcs1_mcs_mat1_1_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_7001, mcs1_mcs_mat1_1_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_8204, mcs1_mcs_mat1_1_mcs_out[29]}), .c ({new_AGEMA_signal_8685, mcs1_mcs_mat1_1_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_7000, mcs1_mcs_mat1_1_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_8203, mcs1_mcs_mat1_1_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_8686, mcs1_mcs_mat1_1_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_7729, mcs1_mcs_mat1_1_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_6613, shiftr_out[120]}), .c ({new_AGEMA_signal_8203, mcs1_mcs_mat1_1_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_8687, mcs1_mcs_mat1_1_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_7727, mcs1_mcs_mat1_1_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_9127, mcs1_mcs_mat1_1_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_8205, mcs1_mcs_mat1_1_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_7728, mcs1_mcs_mat1_1_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_8687, mcs1_mcs_mat1_1_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_7380, mcs1_mcs_mat1_1_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_7728, mcs1_mcs_mat1_1_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_7729, mcs1_mcs_mat1_1_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7001, mcs1_mcs_mat1_1_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_8205, mcs1_mcs_mat1_1_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[592]), .c ({new_AGEMA_signal_7729, mcs1_mcs_mat1_1_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[593]), .c ({new_AGEMA_signal_7001, mcs1_mcs_mat1_1_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[594]), .c ({new_AGEMA_signal_7380, mcs1_mcs_mat1_1_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_7730, mcs1_mcs_mat1_1_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_8206, mcs1_mcs_mat1_1_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_7381, mcs1_mcs_mat1_1_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7002, mcs1_mcs_mat1_1_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_7730, mcs1_mcs_mat1_1_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_8207, mcs1_mcs_mat1_1_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_8688, mcs1_mcs_mat1_1_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_7732, mcs1_mcs_mat1_1_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_7002, mcs1_mcs_mat1_1_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_8207, mcs1_mcs_mat1_1_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_8689, mcs1_mcs_mat1_1_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_6618, shiftr_out[88]}), .c ({new_AGEMA_signal_9128, mcs1_mcs_mat1_1_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_7732, mcs1_mcs_mat1_1_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8208, mcs1_mcs_mat1_1_mcs_out[24]}), .c ({new_AGEMA_signal_8689, mcs1_mcs_mat1_1_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_7731, mcs1_mcs_mat1_1_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_7232, shiftr_out[91]}), .c ({new_AGEMA_signal_8208, mcs1_mcs_mat1_1_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_7381, mcs1_mcs_mat1_1_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_6737, mcs1_mcs_mat1_1_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_7731, mcs1_mcs_mat1_1_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[595]), .c ({new_AGEMA_signal_7732, mcs1_mcs_mat1_1_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[596]), .c ({new_AGEMA_signal_7002, mcs1_mcs_mat1_1_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7232, shiftr_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[597]), .c ({new_AGEMA_signal_7381, mcs1_mcs_mat1_1_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_7733, mcs1_mcs_mat1_1_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_6692, shiftr_out[58]}), .c ({new_AGEMA_signal_8209, mcs1_mcs_mat1_1_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_7382, mcs1_mcs_mat1_1_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7003, mcs1_mcs_mat1_1_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_7733, mcs1_mcs_mat1_1_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_8210, mcs1_mcs_mat1_1_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_7304, shiftr_out[57]}), .c ({new_AGEMA_signal_8690, mcs1_mcs_mat1_1_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_7735, mcs1_mcs_mat1_1_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_7003, mcs1_mcs_mat1_1_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_8210, mcs1_mcs_mat1_1_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_8691, mcs1_mcs_mat1_1_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_6624, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_9129, mcs1_mcs_mat1_1_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_7735, mcs1_mcs_mat1_1_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8211, mcs1_mcs_mat1_1_mcs_out[20]}), .c ({new_AGEMA_signal_8691, mcs1_mcs_mat1_1_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_7734, mcs1_mcs_mat1_1_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_8211, mcs1_mcs_mat1_1_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_7382, mcs1_mcs_mat1_1_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_6738, mcs1_mcs_mat1_1_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_7734, mcs1_mcs_mat1_1_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7304, shiftr_out[57]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[598]), .c ({new_AGEMA_signal_7735, mcs1_mcs_mat1_1_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[599]), .c ({new_AGEMA_signal_7003, mcs1_mcs_mat1_1_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[600]), .c ({new_AGEMA_signal_7382, mcs1_mcs_mat1_1_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_9662, mcs1_mcs_mat1_1_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_9665, mcs1_mcs_mat1_1_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_9899, mcs1_mcs_mat1_1_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_9900, mcs1_mcs_mat1_1_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_8212, mcs1_mcs_mat1_1_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_10113, mcs1_mcs_mat1_1_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_10114, mcs1_mcs_mat1_1_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_8692, mcs1_mcs_mat1_1_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_10357, mcs1_mcs_mat1_1_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_7621, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_9900, mcs1_mcs_mat1_1_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_10114, mcs1_mcs_mat1_1_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_9663, mcs1_mcs_mat1_1_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_9363, shiftr_out[25]}), .c ({new_AGEMA_signal_9900, mcs1_mcs_mat1_1_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_9417, mcs1_mcs_mat1_1_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_9418, mcs1_mcs_mat1_1_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_9663, mcs1_mcs_mat1_1_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_9664, mcs1_mcs_mat1_1_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_8692, mcs1_mcs_mat1_1_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_9901, mcs1_mcs_mat1_1_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9363, shiftr_out[25]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[601]), .c ({new_AGEMA_signal_9665, mcs1_mcs_mat1_1_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[602]), .c ({new_AGEMA_signal_8692, mcs1_mcs_mat1_1_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[603]), .c ({new_AGEMA_signal_9418, mcs1_mcs_mat1_1_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_8695, mcs1_mcs_mat1_1_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_7252, mcs1_mcs_mat1_1_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_9130, mcs1_mcs_mat1_1_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_8215, mcs1_mcs_mat1_1_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_8213, mcs1_mcs_mat1_1_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_8693, mcs1_mcs_mat1_1_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_7737, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_7004, mcs1_mcs_mat1_1_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8213, mcs1_mcs_mat1_1_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_7252, mcs1_mcs_mat1_1_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_8214, mcs1_mcs_mat1_1_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_8694, mcs1_mcs_mat1_1_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_7736, mcs1_mcs_mat1_1_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_7737, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_8214, mcs1_mcs_mat1_1_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_6739, mcs1_mcs_mat1_1_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_7004, mcs1_mcs_mat1_1_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_7252, mcs1_mcs_mat1_1_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_9131, mcs1_mcs_mat1_1_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_9419, mcs1_mcs_mat1_1_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_8695, mcs1_mcs_mat1_1_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_7737, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_9131, mcs1_mcs_mat1_1_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_8215, mcs1_mcs_mat1_1_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_8695, mcs1_mcs_mat1_1_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_7736, mcs1_mcs_mat1_1_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_8215, mcs1_mcs_mat1_1_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_6613, shiftr_out[120]}), .b ({new_AGEMA_signal_7383, mcs1_mcs_mat1_1_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_7736, mcs1_mcs_mat1_1_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7293, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[604]), .c ({new_AGEMA_signal_7737, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6681, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[605]), .c ({new_AGEMA_signal_7004, mcs1_mcs_mat1_1_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7227, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[606]), .c ({new_AGEMA_signal_7383, mcs1_mcs_mat1_1_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_7253, mcs1_mcs_mat1_1_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_7232, shiftr_out[91]}), .c ({new_AGEMA_signal_7384, mcs1_mcs_mat1_1_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_8217, mcs1_mcs_mat1_1_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_8696, mcs1_mcs_mat1_1_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_7738, mcs1_mcs_mat1_1_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_8216, mcs1_mcs_mat1_1_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_7385, mcs1_mcs_mat1_1_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_7253, mcs1_mcs_mat1_1_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_7738, mcs1_mcs_mat1_1_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_6740, mcs1_mcs_mat1_1_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_7005, mcs1_mcs_mat1_1_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_7253, mcs1_mcs_mat1_1_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_8697, mcs1_mcs_mat1_1_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_6618, shiftr_out[88]}), .c ({new_AGEMA_signal_9132, mcs1_mcs_mat1_1_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_6740, mcs1_mcs_mat1_1_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8217, mcs1_mcs_mat1_1_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_8697, mcs1_mcs_mat1_1_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_7739, mcs1_mcs_mat1_1_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_7385, mcs1_mcs_mat1_1_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_8217, mcs1_mcs_mat1_1_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7298, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[607]), .c ({new_AGEMA_signal_7739, mcs1_mcs_mat1_1_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6686, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[608]), .c ({new_AGEMA_signal_7005, mcs1_mcs_mat1_1_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7232, shiftr_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[609]), .c ({new_AGEMA_signal_7385, mcs1_mcs_mat1_1_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_9420, mcs1_mcs_mat1_1_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_7387, mcs1_mcs_mat1_1_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_9666, mcs1_mcs_mat1_1_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_9133, mcs1_mcs_mat1_1_mcs_out[7]}), .b ({new_AGEMA_signal_6692, shiftr_out[58]}), .c ({new_AGEMA_signal_9420, mcs1_mcs_mat1_1_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_8698, mcs1_mcs_mat1_1_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_7304, shiftr_out[57]}), .c ({new_AGEMA_signal_9133, mcs1_mcs_mat1_1_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_8218, mcs1_mcs_mat1_1_mcs_out[6]}), .b ({new_AGEMA_signal_7007, mcs1_mcs_mat1_1_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_8698, mcs1_mcs_mat1_1_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_7006, mcs1_mcs_mat1_1_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_7740, mcs1_mcs_mat1_1_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_8218, mcs1_mcs_mat1_1_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7304, shiftr_out[57]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[610]), .c ({new_AGEMA_signal_7740, mcs1_mcs_mat1_1_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6692, shiftr_out[58]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[611]), .c ({new_AGEMA_signal_7007, mcs1_mcs_mat1_1_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7238, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[612]), .c ({new_AGEMA_signal_7387, mcs1_mcs_mat1_1_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_9421, mcs1_mcs_mat1_1_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_9667, mcs1_mcs_mat1_1_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_9903, mcs1_mcs_mat1_1_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_9363, shiftr_out[25]}), .b ({new_AGEMA_signal_9422, mcs1_mcs_mat1_1_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_9667, mcs1_mcs_mat1_1_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_9904, mcs1_mcs_mat1_1_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_8699, mcs1_mcs_mat1_1_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_10115, mcs1_mcs_mat1_1_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_9905, mcs1_mcs_mat1_1_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_9669, mcs1_mcs_mat1_1_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_10116, mcs1_mcs_mat1_1_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_9670, mcs1_mcs_mat1_1_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_8219, mcs1_mcs_mat1_1_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_9905, mcs1_mcs_mat1_1_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9363, shiftr_out[25]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[613]), .c ({new_AGEMA_signal_9670, mcs1_mcs_mat1_1_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8101, shiftr_out[26]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[614]), .c ({new_AGEMA_signal_8699, mcs1_mcs_mat1_1_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9059, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[615]), .c ({new_AGEMA_signal_9422, mcs1_mcs_mat1_1_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U96 ( .a ({new_AGEMA_signal_10641, mcs1_mcs_mat1_2_n128}), .b ({new_AGEMA_signal_9134, mcs1_mcs_mat1_2_n127}), .c ({temp_next_s1[85], temp_next_s0[85]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U95 ( .a ({new_AGEMA_signal_8735, mcs1_mcs_mat1_2_mcs_out[41]}), .b ({new_AGEMA_signal_7772, mcs1_mcs_mat1_2_mcs_out[45]}), .c ({new_AGEMA_signal_9134, mcs1_mcs_mat1_2_n127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U94 ( .a ({new_AGEMA_signal_7255, mcs1_mcs_mat1_2_mcs_out[33]}), .b ({new_AGEMA_signal_10380, mcs1_mcs_mat1_2_mcs_out[37]}), .c ({new_AGEMA_signal_10641, mcs1_mcs_mat1_2_n128}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U93 ( .a ({new_AGEMA_signal_10117, mcs1_mcs_mat1_2_n126}), .b ({new_AGEMA_signal_9671, mcs1_mcs_mat1_2_n125}), .c ({temp_next_s1[84], temp_next_s0[84]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U92 ( .a ({new_AGEMA_signal_8257, mcs1_mcs_mat1_2_mcs_out[40]}), .b ({new_AGEMA_signal_9447, mcs1_mcs_mat1_2_mcs_out[44]}), .c ({new_AGEMA_signal_9671, mcs1_mcs_mat1_2_n125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U91 ( .a ({new_AGEMA_signal_9451, mcs1_mcs_mat1_2_mcs_out[32]}), .b ({new_AGEMA_signal_9922, mcs1_mcs_mat1_2_mcs_out[36]}), .c ({new_AGEMA_signal_10117, mcs1_mcs_mat1_2_n126}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U90 ( .a ({new_AGEMA_signal_10118, mcs1_mcs_mat1_2_n124}), .b ({new_AGEMA_signal_9423, mcs1_mcs_mat1_2_n123}), .c ({temp_next_s1[55], temp_next_s0[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U89 ( .a ({new_AGEMA_signal_8264, mcs1_mcs_mat1_2_mcs_out[27]}), .b ({new_AGEMA_signal_9164, mcs1_mcs_mat1_2_mcs_out[31]}), .c ({new_AGEMA_signal_9423, mcs1_mcs_mat1_2_n123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U88 ( .a ({new_AGEMA_signal_8268, mcs1_mcs_mat1_2_mcs_out[19]}), .b ({new_AGEMA_signal_9923, mcs1_mcs_mat1_2_mcs_out[23]}), .c ({new_AGEMA_signal_10118, mcs1_mcs_mat1_2_n124}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U87 ( .a ({new_AGEMA_signal_10360, mcs1_mcs_mat1_2_n122}), .b ({new_AGEMA_signal_9135, mcs1_mcs_mat1_2_n121}), .c ({temp_next_s1[54], temp_next_s0[54]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U86 ( .a ({new_AGEMA_signal_8741, mcs1_mcs_mat1_2_mcs_out[26]}), .b ({new_AGEMA_signal_8739, mcs1_mcs_mat1_2_mcs_out[30]}), .c ({new_AGEMA_signal_9135, mcs1_mcs_mat1_2_n121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U85 ( .a ({new_AGEMA_signal_8744, mcs1_mcs_mat1_2_mcs_out[18]}), .b ({new_AGEMA_signal_10139, mcs1_mcs_mat1_2_mcs_out[22]}), .c ({new_AGEMA_signal_10360, mcs1_mcs_mat1_2_n122}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U84 ( .a ({new_AGEMA_signal_10643, mcs1_mcs_mat1_2_n120}), .b ({new_AGEMA_signal_9424, mcs1_mcs_mat1_2_n119}), .c ({temp_next_s1[53], temp_next_s0[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U83 ( .a ({new_AGEMA_signal_9166, mcs1_mcs_mat1_2_mcs_out[25]}), .b ({new_AGEMA_signal_8262, mcs1_mcs_mat1_2_mcs_out[29]}), .c ({new_AGEMA_signal_9424, mcs1_mcs_mat1_2_n119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U82 ( .a ({new_AGEMA_signal_9167, mcs1_mcs_mat1_2_mcs_out[17]}), .b ({new_AGEMA_signal_10381, mcs1_mcs_mat1_2_mcs_out[21]}), .c ({new_AGEMA_signal_10643, mcs1_mcs_mat1_2_n120}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U81 ( .a ({new_AGEMA_signal_10119, mcs1_mcs_mat1_2_n118}), .b ({new_AGEMA_signal_9425, mcs1_mcs_mat1_2_n117}), .c ({temp_next_s1[52], temp_next_s0[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U80 ( .a ({new_AGEMA_signal_8266, mcs1_mcs_mat1_2_mcs_out[24]}), .b ({new_AGEMA_signal_9165, mcs1_mcs_mat1_2_mcs_out[28]}), .c ({new_AGEMA_signal_9425, mcs1_mcs_mat1_2_n117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U79 ( .a ({new_AGEMA_signal_8270, mcs1_mcs_mat1_2_mcs_out[16]}), .b ({new_AGEMA_signal_9925, mcs1_mcs_mat1_2_mcs_out[20]}), .c ({new_AGEMA_signal_10119, mcs1_mcs_mat1_2_n118}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U78 ( .a ({new_AGEMA_signal_9426, mcs1_mcs_mat1_2_n116}), .b ({new_AGEMA_signal_10644, mcs1_mcs_mat1_2_n115}), .c ({temp_next_s1[23], temp_next_s0[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U77 ( .a ({new_AGEMA_signal_8277, mcs1_mcs_mat1_2_mcs_out[3]}), .b ({new_AGEMA_signal_10382, mcs1_mcs_mat1_2_mcs_out[7]}), .c ({new_AGEMA_signal_10644, mcs1_mcs_mat1_2_n115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U76 ( .a ({new_AGEMA_signal_7419, mcs1_mcs_mat1_2_mcs_out[11]}), .b ({new_AGEMA_signal_9168, mcs1_mcs_mat1_2_mcs_out[15]}), .c ({new_AGEMA_signal_9426, mcs1_mcs_mat1_2_n116}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U75 ( .a ({new_AGEMA_signal_10645, mcs1_mcs_mat1_2_n114}), .b ({new_AGEMA_signal_9427, mcs1_mcs_mat1_2_n113}), .c ({new_AGEMA_signal_10886, mcs_out[247]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U74 ( .a ({new_AGEMA_signal_9145, mcs1_mcs_mat1_2_mcs_out[123]}), .b ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_9427, mcs1_mcs_mat1_2_n113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U73 ( .a ({new_AGEMA_signal_8708, mcs1_mcs_mat1_2_mcs_out[115]}), .b ({new_AGEMA_signal_10373, mcs1_mcs_mat1_2_mcs_out[119]}), .c ({new_AGEMA_signal_10645, mcs1_mcs_mat1_2_n114}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U72 ( .a ({new_AGEMA_signal_10646, mcs1_mcs_mat1_2_n112}), .b ({new_AGEMA_signal_8220, mcs1_mcs_mat1_2_n111}), .c ({new_AGEMA_signal_10887, mcs_out[246]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U71 ( .a ({new_AGEMA_signal_7741, mcs1_mcs_mat1_2_mcs_out[122]}), .b ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_8220, mcs1_mcs_mat1_2_n111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U70 ( .a ({new_AGEMA_signal_8226, mcs1_mcs_mat1_2_mcs_out[114]}), .b ({new_AGEMA_signal_10374, mcs1_mcs_mat1_2_mcs_out[118]}), .c ({new_AGEMA_signal_10646, mcs1_mcs_mat1_2_n112}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U69 ( .a ({new_AGEMA_signal_9136, mcs1_mcs_mat1_2_n110}), .b ({new_AGEMA_signal_10120, mcs1_mcs_mat1_2_n109}), .c ({temp_next_s1[22], temp_next_s0[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U68 ( .a ({new_AGEMA_signal_8278, mcs1_mcs_mat1_2_mcs_out[2]}), .b ({new_AGEMA_signal_9926, mcs1_mcs_mat1_2_mcs_out[6]}), .c ({new_AGEMA_signal_10120, mcs1_mcs_mat1_2_n109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U67 ( .a ({new_AGEMA_signal_8749, mcs1_mcs_mat1_2_mcs_out[10]}), .b ({new_AGEMA_signal_8746, mcs1_mcs_mat1_2_mcs_out[14]}), .c ({new_AGEMA_signal_9136, mcs1_mcs_mat1_2_n110}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U66 ( .a ({new_AGEMA_signal_10363, mcs1_mcs_mat1_2_n108}), .b ({new_AGEMA_signal_9428, mcs1_mcs_mat1_2_n107}), .c ({new_AGEMA_signal_10647, mcs_out[245]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U65 ( .a ({new_AGEMA_signal_9146, mcs1_mcs_mat1_2_mcs_out[121]}), .b ({new_AGEMA_signal_7388, mcs1_mcs_mat1_2_mcs_out[125]}), .c ({new_AGEMA_signal_9428, mcs1_mcs_mat1_2_n107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U64 ( .a ({new_AGEMA_signal_7743, mcs1_mcs_mat1_2_mcs_out[113]}), .b ({new_AGEMA_signal_10129, mcs1_mcs_mat1_2_mcs_out[117]}), .c ({new_AGEMA_signal_10363, mcs1_mcs_mat1_2_n108}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U63 ( .a ({new_AGEMA_signal_10121, mcs1_mcs_mat1_2_n106}), .b ({new_AGEMA_signal_9137, mcs1_mcs_mat1_2_n105}), .c ({new_AGEMA_signal_10364, mcs_out[244]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U62 ( .a ({new_AGEMA_signal_8706, mcs1_mcs_mat1_2_mcs_out[120]}), .b ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_9137, mcs1_mcs_mat1_2_n105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U61 ( .a ({new_AGEMA_signal_9147, mcs1_mcs_mat1_2_mcs_out[112]}), .b ({new_AGEMA_signal_9912, mcs1_mcs_mat1_2_mcs_out[116]}), .c ({new_AGEMA_signal_10121, mcs1_mcs_mat1_2_n106}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U60 ( .a ({new_AGEMA_signal_10365, mcs1_mcs_mat1_2_n104}), .b ({new_AGEMA_signal_9429, mcs1_mcs_mat1_2_n103}), .c ({new_AGEMA_signal_10648, mcs_out[215]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U59 ( .a ({new_AGEMA_signal_9148, mcs1_mcs_mat1_2_mcs_out[111]}), .b ({new_AGEMA_signal_9153, mcs1_mcs_mat1_2_mcs_out[99]}), .c ({new_AGEMA_signal_9429, mcs1_mcs_mat1_2_n103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U58 ( .a ({new_AGEMA_signal_10130, mcs1_mcs_mat1_2_mcs_out[103]}), .b ({new_AGEMA_signal_8712, mcs1_mcs_mat1_2_mcs_out[107]}), .c ({new_AGEMA_signal_10365, mcs1_mcs_mat1_2_n104}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U57 ( .a ({new_AGEMA_signal_9906, mcs1_mcs_mat1_2_n102}), .b ({new_AGEMA_signal_9430, mcs1_mcs_mat1_2_n101}), .c ({new_AGEMA_signal_10122, mcs_out[214]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U56 ( .a ({new_AGEMA_signal_9149, mcs1_mcs_mat1_2_mcs_out[110]}), .b ({new_AGEMA_signal_8234, mcs1_mcs_mat1_2_mcs_out[98]}), .c ({new_AGEMA_signal_9430, mcs1_mcs_mat1_2_n101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U55 ( .a ({new_AGEMA_signal_9678, mcs1_mcs_mat1_2_mcs_out[102]}), .b ({new_AGEMA_signal_8713, mcs1_mcs_mat1_2_mcs_out[106]}), .c ({new_AGEMA_signal_9906, mcs1_mcs_mat1_2_n102}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U54 ( .a ({new_AGEMA_signal_10123, mcs1_mcs_mat1_2_n100}), .b ({new_AGEMA_signal_9431, mcs1_mcs_mat1_2_n99}), .c ({new_AGEMA_signal_10366, mcs_out[213]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U53 ( .a ({new_AGEMA_signal_9150, mcs1_mcs_mat1_2_mcs_out[109]}), .b ({new_AGEMA_signal_7396, mcs1_mcs_mat1_2_mcs_out[97]}), .c ({new_AGEMA_signal_9431, mcs1_mcs_mat1_2_n99}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U52 ( .a ({new_AGEMA_signal_9914, mcs1_mcs_mat1_2_mcs_out[101]}), .b ({new_AGEMA_signal_8714, mcs1_mcs_mat1_2_mcs_out[105]}), .c ({new_AGEMA_signal_10123, mcs1_mcs_mat1_2_n100}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U51 ( .a ({new_AGEMA_signal_10367, mcs1_mcs_mat1_2_n98}), .b ({new_AGEMA_signal_9907, mcs1_mcs_mat1_2_n97}), .c ({new_AGEMA_signal_10649, mcs_out[212]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U50 ( .a ({new_AGEMA_signal_9151, mcs1_mcs_mat1_2_mcs_out[108]}), .b ({new_AGEMA_signal_9682, mcs1_mcs_mat1_2_mcs_out[96]}), .c ({new_AGEMA_signal_9907, mcs1_mcs_mat1_2_n97}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U49 ( .a ({new_AGEMA_signal_10131, mcs1_mcs_mat1_2_mcs_out[100]}), .b ({new_AGEMA_signal_9152, mcs1_mcs_mat1_2_mcs_out[104]}), .c ({new_AGEMA_signal_10367, mcs1_mcs_mat1_2_n98}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U48 ( .a ({new_AGEMA_signal_9908, mcs1_mcs_mat1_2_n96}), .b ({new_AGEMA_signal_9138, mcs1_mcs_mat1_2_n95}), .c ({new_AGEMA_signal_10124, mcs_out[183]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U47 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_8718, mcs1_mcs_mat1_2_mcs_out[95]}), .c ({new_AGEMA_signal_9138, mcs1_mcs_mat1_2_n95}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U46 ( .a ({new_AGEMA_signal_8236, mcs1_mcs_mat1_2_mcs_out[83]}), .b ({new_AGEMA_signal_9683, mcs1_mcs_mat1_2_mcs_out[87]}), .c ({new_AGEMA_signal_9908, mcs1_mcs_mat1_2_n96}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U45 ( .a ({new_AGEMA_signal_8700, mcs1_mcs_mat1_2_n94}), .b ({new_AGEMA_signal_8221, mcs1_mcs_mat1_2_n93}), .c ({new_AGEMA_signal_9139, mcs_out[182]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U43 ( .a ({new_AGEMA_signal_8237, mcs1_mcs_mat1_2_mcs_out[82]}), .b ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_8700, mcs1_mcs_mat1_2_n94}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U42 ( .a ({new_AGEMA_signal_9432, mcs1_mcs_mat1_2_n92}), .b ({new_AGEMA_signal_8222, mcs1_mcs_mat1_2_n91}), .c ({new_AGEMA_signal_9672, mcs_out[181]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U41 ( .a ({new_AGEMA_signal_7402, mcs1_mcs_mat1_2_mcs_out[89]}), .b ({new_AGEMA_signal_7752, mcs1_mcs_mat1_2_mcs_out[93]}), .c ({new_AGEMA_signal_8222, mcs1_mcs_mat1_2_n91}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U40 ( .a ({new_AGEMA_signal_8238, mcs1_mcs_mat1_2_mcs_out[81]}), .b ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_9432, mcs1_mcs_mat1_2_n92}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U39 ( .a ({new_AGEMA_signal_10125, mcs1_mcs_mat1_2_n90}), .b ({new_AGEMA_signal_9433, mcs1_mcs_mat1_2_n89}), .c ({new_AGEMA_signal_10368, mcs_out[180]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U38 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_9154, mcs1_mcs_mat1_2_mcs_out[92]}), .c ({new_AGEMA_signal_9433, mcs1_mcs_mat1_2_n89}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U37 ( .a ({new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[80]}), .b ({new_AGEMA_signal_9916, mcs1_mcs_mat1_2_mcs_out[84]}), .c ({new_AGEMA_signal_10125, mcs1_mcs_mat1_2_n90}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U36 ( .a ({new_AGEMA_signal_9140, mcs1_mcs_mat1_2_n88}), .b ({new_AGEMA_signal_9673, mcs1_mcs_mat1_2_n87}), .c ({temp_next_s1[21], temp_next_s0[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U35 ( .a ({new_AGEMA_signal_9454, mcs1_mcs_mat1_2_mcs_out[5]}), .b ({new_AGEMA_signal_8274, mcs1_mcs_mat1_2_mcs_out[9]}), .c ({new_AGEMA_signal_9673, mcs1_mcs_mat1_2_n87}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U34 ( .a ({new_AGEMA_signal_8747, mcs1_mcs_mat1_2_mcs_out[13]}), .b ({new_AGEMA_signal_8753, mcs1_mcs_mat1_2_mcs_out[1]}), .c ({new_AGEMA_signal_9140, mcs1_mcs_mat1_2_n88}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U33 ( .a ({new_AGEMA_signal_10369, mcs1_mcs_mat1_2_n86}), .b ({new_AGEMA_signal_9141, mcs1_mcs_mat1_2_n85}), .c ({new_AGEMA_signal_10650, mcs_out[151]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U32 ( .a ({new_AGEMA_signal_7760, mcs1_mcs_mat1_2_mcs_out[75]}), .b ({new_AGEMA_signal_8721, mcs1_mcs_mat1_2_mcs_out[79]}), .c ({new_AGEMA_signal_9141, mcs1_mcs_mat1_2_n85}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U31 ( .a ({new_AGEMA_signal_9158, mcs1_mcs_mat1_2_mcs_out[67]}), .b ({new_AGEMA_signal_10132, mcs1_mcs_mat1_2_mcs_out[71]}), .c ({new_AGEMA_signal_10369, mcs1_mcs_mat1_2_n86}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U30 ( .a ({new_AGEMA_signal_10651, mcs1_mcs_mat1_2_n84}), .b ({new_AGEMA_signal_9434, mcs1_mcs_mat1_2_n83}), .c ({new_AGEMA_signal_10888, mcs_out[150]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U29 ( .a ({new_AGEMA_signal_9156, mcs1_mcs_mat1_2_mcs_out[74]}), .b ({new_AGEMA_signal_7018, mcs1_mcs_mat1_2_mcs_out[78]}), .c ({new_AGEMA_signal_9434, mcs1_mcs_mat1_2_n83}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U28 ( .a ({new_AGEMA_signal_8726, mcs1_mcs_mat1_2_mcs_out[66]}), .b ({new_AGEMA_signal_10375, mcs1_mcs_mat1_2_mcs_out[70]}), .c ({new_AGEMA_signal_10651, mcs1_mcs_mat1_2_n84}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U27 ( .a ({new_AGEMA_signal_10652, mcs1_mcs_mat1_2_n82}), .b ({new_AGEMA_signal_8701, mcs1_mcs_mat1_2_n81}), .c ({new_AGEMA_signal_10889, mcs_out[149]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U26 ( .a ({new_AGEMA_signal_8241, mcs1_mcs_mat1_2_mcs_out[73]}), .b ({new_AGEMA_signal_7758, mcs1_mcs_mat1_2_mcs_out[77]}), .c ({new_AGEMA_signal_8701, mcs1_mcs_mat1_2_n81}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U25 ( .a ({new_AGEMA_signal_7763, mcs1_mcs_mat1_2_mcs_out[65]}), .b ({new_AGEMA_signal_10376, mcs1_mcs_mat1_2_mcs_out[69]}), .c ({new_AGEMA_signal_10652, mcs1_mcs_mat1_2_n82}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U24 ( .a ({new_AGEMA_signal_10370, mcs1_mcs_mat1_2_n80}), .b ({new_AGEMA_signal_9435, mcs1_mcs_mat1_2_n79}), .c ({new_AGEMA_signal_10653, mcs_out[148]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U23 ( .a ({new_AGEMA_signal_9157, mcs1_mcs_mat1_2_mcs_out[72]}), .b ({new_AGEMA_signal_9155, mcs1_mcs_mat1_2_mcs_out[76]}), .c ({new_AGEMA_signal_9435, mcs1_mcs_mat1_2_n79}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U22 ( .a ({new_AGEMA_signal_9445, mcs1_mcs_mat1_2_mcs_out[64]}), .b ({new_AGEMA_signal_10134, mcs1_mcs_mat1_2_mcs_out[68]}), .c ({new_AGEMA_signal_10370, mcs1_mcs_mat1_2_n80}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U21 ( .a ({new_AGEMA_signal_10371, mcs1_mcs_mat1_2_n78}), .b ({new_AGEMA_signal_9142, mcs1_mcs_mat1_2_n77}), .c ({temp_next_s1[119], temp_next_s0[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U20 ( .a ({new_AGEMA_signal_8248, mcs1_mcs_mat1_2_mcs_out[59]}), .b ({new_AGEMA_signal_8728, mcs1_mcs_mat1_2_mcs_out[63]}), .c ({new_AGEMA_signal_9142, mcs1_mcs_mat1_2_n77}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U19 ( .a ({new_AGEMA_signal_7771, mcs1_mcs_mat1_2_mcs_out[51]}), .b ({new_AGEMA_signal_10135, mcs1_mcs_mat1_2_mcs_out[55]}), .c ({new_AGEMA_signal_10371, mcs1_mcs_mat1_2_n78}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U18 ( .a ({new_AGEMA_signal_10655, mcs1_mcs_mat1_2_n76}), .b ({new_AGEMA_signal_8702, mcs1_mcs_mat1_2_n75}), .c ({temp_next_s1[118], temp_next_s0[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U17 ( .a ({new_AGEMA_signal_7767, mcs1_mcs_mat1_2_mcs_out[58]}), .b ({new_AGEMA_signal_8245, mcs1_mcs_mat1_2_mcs_out[62]}), .c ({new_AGEMA_signal_8702, mcs1_mcs_mat1_2_n75}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U16 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_10377, mcs1_mcs_mat1_2_mcs_out[54]}), .c ({new_AGEMA_signal_10655, mcs1_mcs_mat1_2_n76}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U15 ( .a ({new_AGEMA_signal_10656, mcs1_mcs_mat1_2_n74}), .b ({new_AGEMA_signal_8703, mcs1_mcs_mat1_2_n73}), .c ({temp_next_s1[117], temp_next_s0[117]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U14 ( .a ({new_AGEMA_signal_8249, mcs1_mcs_mat1_2_mcs_out[57]}), .b ({new_AGEMA_signal_8246, mcs1_mcs_mat1_2_mcs_out[61]}), .c ({new_AGEMA_signal_8703, mcs1_mcs_mat1_2_n73}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U13 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_10378, mcs1_mcs_mat1_2_mcs_out[53]}), .c ({new_AGEMA_signal_10656, mcs1_mcs_mat1_2_n74}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U12 ( .a ({new_AGEMA_signal_10372, mcs1_mcs_mat1_2_n72}), .b ({new_AGEMA_signal_9436, mcs1_mcs_mat1_2_n71}), .c ({temp_next_s1[116], temp_next_s0[116]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U11 ( .a ({new_AGEMA_signal_8730, mcs1_mcs_mat1_2_mcs_out[56]}), .b ({new_AGEMA_signal_9160, mcs1_mcs_mat1_2_mcs_out[60]}), .c ({new_AGEMA_signal_9436, mcs1_mcs_mat1_2_n71}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U10 ( .a ({new_AGEMA_signal_8252, mcs1_mcs_mat1_2_mcs_out[48]}), .b ({new_AGEMA_signal_10137, mcs1_mcs_mat1_2_mcs_out[52]}), .c ({new_AGEMA_signal_10372, mcs1_mcs_mat1_2_n72}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U9 ( .a ({new_AGEMA_signal_10658, mcs1_mcs_mat1_2_n70}), .b ({new_AGEMA_signal_9143, mcs1_mcs_mat1_2_n69}), .c ({temp_next_s1[87], temp_next_s0[87]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U8 ( .a ({new_AGEMA_signal_8733, mcs1_mcs_mat1_2_mcs_out[43]}), .b ({new_AGEMA_signal_8732, mcs1_mcs_mat1_2_mcs_out[47]}), .c ({new_AGEMA_signal_9143, mcs1_mcs_mat1_2_n69}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U7 ( .a ({new_AGEMA_signal_8737, mcs1_mcs_mat1_2_mcs_out[35]}), .b ({new_AGEMA_signal_10379, mcs1_mcs_mat1_2_mcs_out[39]}), .c ({new_AGEMA_signal_10658, mcs1_mcs_mat1_2_n70}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U6 ( .a ({new_AGEMA_signal_9910, mcs1_mcs_mat1_2_n68}), .b ({new_AGEMA_signal_9144, mcs1_mcs_mat1_2_n67}), .c ({temp_next_s1[86], temp_next_s0[86]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U5 ( .a ({new_AGEMA_signal_8734, mcs1_mcs_mat1_2_mcs_out[42]}), .b ({new_AGEMA_signal_7409, mcs1_mcs_mat1_2_mcs_out[46]}), .c ({new_AGEMA_signal_9144, mcs1_mcs_mat1_2_n67}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U4 ( .a ({new_AGEMA_signal_8259, mcs1_mcs_mat1_2_mcs_out[34]}), .b ({new_AGEMA_signal_9691, mcs1_mcs_mat1_2_mcs_out[38]}), .c ({new_AGEMA_signal_9910, mcs1_mcs_mat1_2_n68}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U3 ( .a ({new_AGEMA_signal_9674, mcs1_mcs_mat1_2_n66}), .b ({new_AGEMA_signal_11049, mcs1_mcs_mat1_2_n65}), .c ({temp_next_s1[20], temp_next_s0[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U2 ( .a ({new_AGEMA_signal_10893, mcs1_mcs_mat1_2_mcs_out[4]}), .b ({new_AGEMA_signal_9170, mcs1_mcs_mat1_2_mcs_out[8]}), .c ({new_AGEMA_signal_11049, mcs1_mcs_mat1_2_n65}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_U1 ( .a ({new_AGEMA_signal_8754, mcs1_mcs_mat1_2_mcs_out[0]}), .b ({new_AGEMA_signal_9453, mcs1_mcs_mat1_2_mcs_out[12]}), .c ({new_AGEMA_signal_9674, mcs1_mcs_mat1_2_n66}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_8704, mcs1_mcs_mat1_2_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_9145, mcs1_mcs_mat1_2_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_8223, mcs1_mcs_mat1_2_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_6742, mcs1_mcs_mat1_2_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8704, mcs1_mcs_mat1_2_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_7008, mcs1_mcs_mat1_2_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_7389, mcs1_mcs_mat1_2_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_7741, mcs1_mcs_mat1_2_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_7009, mcs1_mcs_mat1_2_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_7231, shiftr_out[87]}), .c ({new_AGEMA_signal_7389, mcs1_mcs_mat1_2_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_8705, mcs1_mcs_mat1_2_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_7231, shiftr_out[87]}), .c ({new_AGEMA_signal_9146, mcs1_mcs_mat1_2_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_8223, mcs1_mcs_mat1_2_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_8705, mcs1_mcs_mat1_2_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_7742, mcs1_mcs_mat1_2_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_7390, mcs1_mcs_mat1_2_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_8223, mcs1_mcs_mat1_2_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_8224, mcs1_mcs_mat1_2_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_8706, mcs1_mcs_mat1_2_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_7742, mcs1_mcs_mat1_2_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_7009, mcs1_mcs_mat1_2_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_8224, mcs1_mcs_mat1_2_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[616]), .c ({new_AGEMA_signal_7742, mcs1_mcs_mat1_2_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[617]), .c ({new_AGEMA_signal_7009, mcs1_mcs_mat1_2_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7231, shiftr_out[87]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[618]), .c ({new_AGEMA_signal_7390, mcs1_mcs_mat1_2_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_10127, mcs1_mcs_mat1_2_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_8099, shiftr_out[54]}), .c ({new_AGEMA_signal_10373, mcs1_mcs_mat1_2_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_9911, mcs1_mcs_mat1_2_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9439, mcs1_mcs_mat1_2_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_10127, mcs1_mcs_mat1_2_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_10128, mcs1_mcs_mat1_2_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_9676, mcs1_mcs_mat1_2_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_10374, mcs1_mcs_mat1_2_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_9911, mcs1_mcs_mat1_2_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9361, shiftr_out[53]}), .c ({new_AGEMA_signal_10128, mcs1_mcs_mat1_2_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_9911, mcs1_mcs_mat1_2_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9675, mcs1_mcs_mat1_2_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_10129, mcs1_mcs_mat1_2_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_9677, mcs1_mcs_mat1_2_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_8707, mcs1_mcs_mat1_2_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_9911, mcs1_mcs_mat1_2_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_9438, mcs1_mcs_mat1_2_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_9676, mcs1_mcs_mat1_2_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_9912, mcs1_mcs_mat1_2_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_8225, mcs1_mcs_mat1_2_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_9439, mcs1_mcs_mat1_2_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_9676, mcs1_mcs_mat1_2_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_8707, mcs1_mcs_mat1_2_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_9438, mcs1_mcs_mat1_2_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9361, shiftr_out[53]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[619]), .c ({new_AGEMA_signal_9677, mcs1_mcs_mat1_2_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[620]), .c ({new_AGEMA_signal_8707, mcs1_mcs_mat1_2_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[621]), .c ({new_AGEMA_signal_9439, mcs1_mcs_mat1_2_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_8227, mcs1_mcs_mat1_2_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_7010, mcs1_mcs_mat1_2_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_8708, mcs1_mcs_mat1_2_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_7391, mcs1_mcs_mat1_2_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_7392, mcs1_mcs_mat1_2_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_7743, mcs1_mcs_mat1_2_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_8228, mcs1_mcs_mat1_2_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_8709, mcs1_mcs_mat1_2_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_9147, mcs1_mcs_mat1_2_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_8227, mcs1_mcs_mat1_2_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_8709, mcs1_mcs_mat1_2_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_6743, mcs1_mcs_mat1_2_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_7745, mcs1_mcs_mat1_2_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_8227, mcs1_mcs_mat1_2_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_7011, mcs1_mcs_mat1_2_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_7744, mcs1_mcs_mat1_2_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8228, mcs1_mcs_mat1_2_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7310, shiftr_out[21]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[622]), .c ({new_AGEMA_signal_7745, mcs1_mcs_mat1_2_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[623]), .c ({new_AGEMA_signal_7011, mcs1_mcs_mat1_2_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[624]), .c ({new_AGEMA_signal_7392, mcs1_mcs_mat1_2_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({new_AGEMA_signal_8710, mcs1_mcs_mat1_2_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9148, mcs1_mcs_mat1_2_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({new_AGEMA_signal_8711, mcs1_mcs_mat1_2_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9149, mcs1_mcs_mat1_2_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_7393, mcs1_mcs_mat1_2_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_8710, mcs1_mcs_mat1_2_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9150, mcs1_mcs_mat1_2_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_7012, mcs1_mcs_mat1_2_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_8229, mcs1_mcs_mat1_2_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_8710, mcs1_mcs_mat1_2_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_7746, mcs1_mcs_mat1_2_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8711, mcs1_mcs_mat1_2_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9151, mcs1_mcs_mat1_2_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_8230, mcs1_mcs_mat1_2_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_8711, mcs1_mcs_mat1_2_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_7393, mcs1_mcs_mat1_2_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_7747, mcs1_mcs_mat1_2_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_8230, mcs1_mcs_mat1_2_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[625]), .c ({new_AGEMA_signal_7747, mcs1_mcs_mat1_2_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[626]), .c ({new_AGEMA_signal_7012, mcs1_mcs_mat1_2_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[627]), .c ({new_AGEMA_signal_7393, mcs1_mcs_mat1_2_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_8232, mcs1_mcs_mat1_2_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_8231, mcs1_mcs_mat1_2_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8712, mcs1_mcs_mat1_2_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_8231, mcs1_mcs_mat1_2_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_7394, mcs1_mcs_mat1_2_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_8713, mcs1_mcs_mat1_2_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_7013, mcs1_mcs_mat1_2_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7231, shiftr_out[87]}), .c ({new_AGEMA_signal_7394, mcs1_mcs_mat1_2_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_8231, mcs1_mcs_mat1_2_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8714, mcs1_mcs_mat1_2_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_7749, mcs1_mcs_mat1_2_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_6745, mcs1_mcs_mat1_2_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_8231, mcs1_mcs_mat1_2_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_8715, mcs1_mcs_mat1_2_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_9152, mcs1_mcs_mat1_2_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_8232, mcs1_mcs_mat1_2_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_7749, mcs1_mcs_mat1_2_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_8715, mcs1_mcs_mat1_2_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_7748, mcs1_mcs_mat1_2_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_6617, shiftr_out[84]}), .c ({new_AGEMA_signal_8232, mcs1_mcs_mat1_2_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_7013, mcs1_mcs_mat1_2_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7395, mcs1_mcs_mat1_2_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_7748, mcs1_mcs_mat1_2_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[628]), .c ({new_AGEMA_signal_7749, mcs1_mcs_mat1_2_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[629]), .c ({new_AGEMA_signal_7013, mcs1_mcs_mat1_2_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7231, shiftr_out[87]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[630]), .c ({new_AGEMA_signal_7395, mcs1_mcs_mat1_2_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_9440, mcs1_mcs_mat1_2_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_9913, mcs1_mcs_mat1_2_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_10130, mcs1_mcs_mat1_2_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_9681, mcs1_mcs_mat1_2_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_9913, mcs1_mcs_mat1_2_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_9679, mcs1_mcs_mat1_2_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_9441, mcs1_mcs_mat1_2_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_9914, mcs1_mcs_mat1_2_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_9680, mcs1_mcs_mat1_2_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_9915, mcs1_mcs_mat1_2_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_10131, mcs1_mcs_mat1_2_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_8233, mcs1_mcs_mat1_2_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_9681, mcs1_mcs_mat1_2_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_9915, mcs1_mcs_mat1_2_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_8716, mcs1_mcs_mat1_2_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_9361, shiftr_out[53]}), .c ({new_AGEMA_signal_9680, mcs1_mcs_mat1_2_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9361, shiftr_out[53]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[631]), .c ({new_AGEMA_signal_9681, mcs1_mcs_mat1_2_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[632]), .c ({new_AGEMA_signal_8716, mcs1_mcs_mat1_2_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[633]), .c ({new_AGEMA_signal_9441, mcs1_mcs_mat1_2_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_9442, mcs1_mcs_mat1_2_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_7397, mcs1_mcs_mat1_2_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_9682, mcs1_mcs_mat1_2_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_9153, mcs1_mcs_mat1_2_mcs_out[99]}), .b ({new_AGEMA_signal_6698, shiftr_out[22]}), .c ({new_AGEMA_signal_9442, mcs1_mcs_mat1_2_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_8717, mcs1_mcs_mat1_2_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_7310, shiftr_out[21]}), .c ({new_AGEMA_signal_9153, mcs1_mcs_mat1_2_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_8234, mcs1_mcs_mat1_2_mcs_out[98]}), .b ({new_AGEMA_signal_7015, mcs1_mcs_mat1_2_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_8717, mcs1_mcs_mat1_2_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_7014, mcs1_mcs_mat1_2_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_7750, mcs1_mcs_mat1_2_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_8234, mcs1_mcs_mat1_2_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7310, shiftr_out[21]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[634]), .c ({new_AGEMA_signal_7750, mcs1_mcs_mat1_2_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[635]), .c ({new_AGEMA_signal_7015, mcs1_mcs_mat1_2_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[636]), .c ({new_AGEMA_signal_7397, mcs1_mcs_mat1_2_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_8235, mcs1_mcs_mat1_2_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_8718, mcs1_mcs_mat1_2_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_7399, mcs1_mcs_mat1_2_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_7400, mcs1_mcs_mat1_2_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_7752, mcs1_mcs_mat1_2_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_8719, mcs1_mcs_mat1_2_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_7016, mcs1_mcs_mat1_2_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_9154, mcs1_mcs_mat1_2_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_8235, mcs1_mcs_mat1_2_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_8719, mcs1_mcs_mat1_2_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_6747, mcs1_mcs_mat1_2_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7753, mcs1_mcs_mat1_2_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_8235, mcs1_mcs_mat1_2_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[637]), .c ({new_AGEMA_signal_7753, mcs1_mcs_mat1_2_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[638]), .c ({new_AGEMA_signal_7016, mcs1_mcs_mat1_2_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[639]), .c ({new_AGEMA_signal_7400, mcs1_mcs_mat1_2_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_7756, mcs1_mcs_mat1_2_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_7757, mcs1_mcs_mat1_2_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_8236, mcs1_mcs_mat1_2_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_7754, mcs1_mcs_mat1_2_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_6748, mcs1_mcs_mat1_2_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_8237, mcs1_mcs_mat1_2_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_7403, mcs1_mcs_mat1_2_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_7754, mcs1_mcs_mat1_2_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_7755, mcs1_mcs_mat1_2_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_8238, mcs1_mcs_mat1_2_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_7017, mcs1_mcs_mat1_2_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_7403, mcs1_mcs_mat1_2_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_7755, mcs1_mcs_mat1_2_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_8239, mcs1_mcs_mat1_2_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_6698, shiftr_out[22]}), .c ({new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_7756, mcs1_mcs_mat1_2_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_7017, mcs1_mcs_mat1_2_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_8239, mcs1_mcs_mat1_2_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7310, shiftr_out[21]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[640]), .c ({new_AGEMA_signal_7757, mcs1_mcs_mat1_2_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[641]), .c ({new_AGEMA_signal_7017, mcs1_mcs_mat1_2_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[642]), .c ({new_AGEMA_signal_7403, mcs1_mcs_mat1_2_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_8240, mcs1_mcs_mat1_2_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_8721, mcs1_mcs_mat1_2_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_7404, mcs1_mcs_mat1_2_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_7758, mcs1_mcs_mat1_2_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_8722, mcs1_mcs_mat1_2_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_7019, mcs1_mcs_mat1_2_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_9155, mcs1_mcs_mat1_2_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_8240, mcs1_mcs_mat1_2_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_6612, shiftr_out[116]}), .c ({new_AGEMA_signal_8722, mcs1_mcs_mat1_2_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_6749, mcs1_mcs_mat1_2_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7759, mcs1_mcs_mat1_2_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_8240, mcs1_mcs_mat1_2_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[643]), .c ({new_AGEMA_signal_7759, mcs1_mcs_mat1_2_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[644]), .c ({new_AGEMA_signal_7019, mcs1_mcs_mat1_2_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[645]), .c ({new_AGEMA_signal_7404, mcs1_mcs_mat1_2_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_8723, mcs1_mcs_mat1_2_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_9156, mcs1_mcs_mat1_2_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_8242, mcs1_mcs_mat1_2_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7761, mcs1_mcs_mat1_2_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_8723, mcs1_mcs_mat1_2_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_7254, mcs1_mcs_mat1_2_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_7760, mcs1_mcs_mat1_2_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_7761, mcs1_mcs_mat1_2_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_7254, mcs1_mcs_mat1_2_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_8241, mcs1_mcs_mat1_2_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_7020, mcs1_mcs_mat1_2_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_7021, mcs1_mcs_mat1_2_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_7254, mcs1_mcs_mat1_2_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_7405, mcs1_mcs_mat1_2_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_6617, shiftr_out[84]}), .c ({new_AGEMA_signal_7761, mcs1_mcs_mat1_2_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_8724, mcs1_mcs_mat1_2_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_7020, mcs1_mcs_mat1_2_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_9157, mcs1_mcs_mat1_2_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_8242, mcs1_mcs_mat1_2_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7405, mcs1_mcs_mat1_2_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_8724, mcs1_mcs_mat1_2_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_7231, shiftr_out[87]}), .b ({new_AGEMA_signal_7762, mcs1_mcs_mat1_2_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_8242, mcs1_mcs_mat1_2_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[646]), .c ({new_AGEMA_signal_7762, mcs1_mcs_mat1_2_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[647]), .c ({new_AGEMA_signal_7021, mcs1_mcs_mat1_2_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7231, shiftr_out[87]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[648]), .c ({new_AGEMA_signal_7405, mcs1_mcs_mat1_2_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_9917, mcs1_mcs_mat1_2_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_9443, mcs1_mcs_mat1_2_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_10132, mcs1_mcs_mat1_2_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_9685, mcs1_mcs_mat1_2_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_10133, mcs1_mcs_mat1_2_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_10375, mcs1_mcs_mat1_2_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_9917, mcs1_mcs_mat1_2_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_10133, mcs1_mcs_mat1_2_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_10376, mcs1_mcs_mat1_2_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_9443, mcs1_mcs_mat1_2_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_9918, mcs1_mcs_mat1_2_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_10133, mcs1_mcs_mat1_2_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({new_AGEMA_signal_8725, mcs1_mcs_mat1_2_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_9443, mcs1_mcs_mat1_2_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_9684, mcs1_mcs_mat1_2_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_9361, shiftr_out[53]}), .c ({new_AGEMA_signal_9917, mcs1_mcs_mat1_2_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_9444, mcs1_mcs_mat1_2_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8243, mcs1_mcs_mat1_2_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_9684, mcs1_mcs_mat1_2_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_9918, mcs1_mcs_mat1_2_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_9685, mcs1_mcs_mat1_2_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_10134, mcs1_mcs_mat1_2_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_9444, mcs1_mcs_mat1_2_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_9685, mcs1_mcs_mat1_2_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({new_AGEMA_signal_9686, mcs1_mcs_mat1_2_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_9918, mcs1_mcs_mat1_2_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9361, shiftr_out[53]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[649]), .c ({new_AGEMA_signal_9686, mcs1_mcs_mat1_2_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[650]), .c ({new_AGEMA_signal_8725, mcs1_mcs_mat1_2_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[651]), .c ({new_AGEMA_signal_9444, mcs1_mcs_mat1_2_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_8727, mcs1_mcs_mat1_2_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_9158, mcs1_mcs_mat1_2_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({new_AGEMA_signal_8244, mcs1_mcs_mat1_2_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_8726, mcs1_mcs_mat1_2_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_9159, mcs1_mcs_mat1_2_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_7406, mcs1_mcs_mat1_2_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_9445, mcs1_mcs_mat1_2_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_8727, mcs1_mcs_mat1_2_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .c ({new_AGEMA_signal_9159, mcs1_mcs_mat1_2_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_7022, mcs1_mcs_mat1_2_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_8244, mcs1_mcs_mat1_2_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_8727, mcs1_mcs_mat1_2_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_6751, mcs1_mcs_mat1_2_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7764, mcs1_mcs_mat1_2_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_8244, mcs1_mcs_mat1_2_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7310, shiftr_out[21]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[652]), .c ({new_AGEMA_signal_7764, mcs1_mcs_mat1_2_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[653]), .c ({new_AGEMA_signal_7022, mcs1_mcs_mat1_2_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[654]), .c ({new_AGEMA_signal_7406, mcs1_mcs_mat1_2_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_8247, mcs1_mcs_mat1_2_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7407, mcs1_mcs_mat1_2_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_8728, mcs1_mcs_mat1_2_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_7023, mcs1_mcs_mat1_2_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_7765, mcs1_mcs_mat1_2_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8245, mcs1_mcs_mat1_2_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({new_AGEMA_signal_7766, mcs1_mcs_mat1_2_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_8246, mcs1_mcs_mat1_2_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[655]), .c ({new_AGEMA_signal_7766, mcs1_mcs_mat1_2_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[656]), .c ({new_AGEMA_signal_7023, mcs1_mcs_mat1_2_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[657]), .c ({new_AGEMA_signal_7407, mcs1_mcs_mat1_2_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_7025, mcs1_mcs_mat1_2_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_7408, mcs1_mcs_mat1_2_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_7767, mcs1_mcs_mat1_2_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_7026, mcs1_mcs_mat1_2_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_7768, mcs1_mcs_mat1_2_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_8249, mcs1_mcs_mat1_2_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_8250, mcs1_mcs_mat1_2_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_7769, mcs1_mcs_mat1_2_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_8730, mcs1_mcs_mat1_2_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_7770, mcs1_mcs_mat1_2_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_8250, mcs1_mcs_mat1_2_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[658]), .c ({new_AGEMA_signal_7770, mcs1_mcs_mat1_2_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[659]), .c ({new_AGEMA_signal_7026, mcs1_mcs_mat1_2_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7231, shiftr_out[87]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[660]), .c ({new_AGEMA_signal_7408, mcs1_mcs_mat1_2_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_9688, mcs1_mcs_mat1_2_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_9919, mcs1_mcs_mat1_2_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_10135, mcs1_mcs_mat1_2_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_10136, mcs1_mcs_mat1_2_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_9687, mcs1_mcs_mat1_2_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_10377, mcs1_mcs_mat1_2_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_9446, mcs1_mcs_mat1_2_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_9687, mcs1_mcs_mat1_2_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({new_AGEMA_signal_10136, mcs1_mcs_mat1_2_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_10378, mcs1_mcs_mat1_2_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_8251, mcs1_mcs_mat1_2_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_9919, mcs1_mcs_mat1_2_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_10136, mcs1_mcs_mat1_2_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_8731, mcs1_mcs_mat1_2_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_9690, mcs1_mcs_mat1_2_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_9919, mcs1_mcs_mat1_2_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_9689, mcs1_mcs_mat1_2_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_9920, mcs1_mcs_mat1_2_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_10137, mcs1_mcs_mat1_2_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_9688, mcs1_mcs_mat1_2_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8731, mcs1_mcs_mat1_2_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_9920, mcs1_mcs_mat1_2_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_9446, mcs1_mcs_mat1_2_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_9688, mcs1_mcs_mat1_2_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9361, shiftr_out[53]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[661]), .c ({new_AGEMA_signal_9690, mcs1_mcs_mat1_2_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[662]), .c ({new_AGEMA_signal_8731, mcs1_mcs_mat1_2_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[663]), .c ({new_AGEMA_signal_9446, mcs1_mcs_mat1_2_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_7410, mcs1_mcs_mat1_2_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_7772, mcs1_mcs_mat1_2_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_9161, mcs1_mcs_mat1_2_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_7027, mcs1_mcs_mat1_2_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_9447, mcs1_mcs_mat1_2_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_8732, mcs1_mcs_mat1_2_mcs_out[47]}), .b ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_9161, mcs1_mcs_mat1_2_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_8253, mcs1_mcs_mat1_2_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_6612, shiftr_out[116]}), .c ({new_AGEMA_signal_8732, mcs1_mcs_mat1_2_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_6754, mcs1_mcs_mat1_2_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_7773, mcs1_mcs_mat1_2_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_8253, mcs1_mcs_mat1_2_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[664]), .c ({new_AGEMA_signal_7773, mcs1_mcs_mat1_2_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[665]), .c ({new_AGEMA_signal_7027, mcs1_mcs_mat1_2_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[666]), .c ({new_AGEMA_signal_7410, mcs1_mcs_mat1_2_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_8254, mcs1_mcs_mat1_2_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_7411, mcs1_mcs_mat1_2_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_8733, mcs1_mcs_mat1_2_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_7774, mcs1_mcs_mat1_2_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7028, mcs1_mcs_mat1_2_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_8254, mcs1_mcs_mat1_2_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_8255, mcs1_mcs_mat1_2_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_7776, mcs1_mcs_mat1_2_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_8734, mcs1_mcs_mat1_2_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_8256, mcs1_mcs_mat1_2_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_6755, mcs1_mcs_mat1_2_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_8735, mcs1_mcs_mat1_2_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_7774, mcs1_mcs_mat1_2_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7412, mcs1_mcs_mat1_2_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8256, mcs1_mcs_mat1_2_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_7775, mcs1_mcs_mat1_2_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_7412, mcs1_mcs_mat1_2_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8257, mcs1_mcs_mat1_2_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[667]), .c ({new_AGEMA_signal_7776, mcs1_mcs_mat1_2_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[668]), .c ({new_AGEMA_signal_7028, mcs1_mcs_mat1_2_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7231, shiftr_out[87]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[669]), .c ({new_AGEMA_signal_7412, mcs1_mcs_mat1_2_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_10138, mcs1_mcs_mat1_2_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_8258, mcs1_mcs_mat1_2_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_10379, mcs1_mcs_mat1_2_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_9449, mcs1_mcs_mat1_2_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_9448, mcs1_mcs_mat1_2_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_9691, mcs1_mcs_mat1_2_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({new_AGEMA_signal_10138, mcs1_mcs_mat1_2_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_10380, mcs1_mcs_mat1_2_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_9692, mcs1_mcs_mat1_2_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_9921, mcs1_mcs_mat1_2_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_10138, mcs1_mcs_mat1_2_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_9693, mcs1_mcs_mat1_2_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9450, mcs1_mcs_mat1_2_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_9921, mcs1_mcs_mat1_2_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_9693, mcs1_mcs_mat1_2_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9449, mcs1_mcs_mat1_2_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_9922, mcs1_mcs_mat1_2_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_9162, mcs1_mcs_mat1_2_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_9449, mcs1_mcs_mat1_2_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({new_AGEMA_signal_8736, mcs1_mcs_mat1_2_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_9162, mcs1_mcs_mat1_2_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9361, shiftr_out[53]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[670]), .c ({new_AGEMA_signal_9693, mcs1_mcs_mat1_2_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[671]), .c ({new_AGEMA_signal_8736, mcs1_mcs_mat1_2_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[672]), .c ({new_AGEMA_signal_9450, mcs1_mcs_mat1_2_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_7777, mcs1_mcs_mat1_2_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7413, mcs1_mcs_mat1_2_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_8259, mcs1_mcs_mat1_2_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_7029, mcs1_mcs_mat1_2_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_7255, mcs1_mcs_mat1_2_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_9163, mcs1_mcs_mat1_2_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_7778, mcs1_mcs_mat1_2_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_9451, mcs1_mcs_mat1_2_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7310, shiftr_out[21]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[673]), .c ({new_AGEMA_signal_7778, mcs1_mcs_mat1_2_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[674]), .c ({new_AGEMA_signal_7029, mcs1_mcs_mat1_2_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[675]), .c ({new_AGEMA_signal_7413, mcs1_mcs_mat1_2_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_8738, mcs1_mcs_mat1_2_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_8261, mcs1_mcs_mat1_2_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_9164, mcs1_mcs_mat1_2_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_7031, mcs1_mcs_mat1_2_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_8262, mcs1_mcs_mat1_2_mcs_out[29]}), .c ({new_AGEMA_signal_8738, mcs1_mcs_mat1_2_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_7030, mcs1_mcs_mat1_2_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_8261, mcs1_mcs_mat1_2_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_8739, mcs1_mcs_mat1_2_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_7781, mcs1_mcs_mat1_2_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_6612, shiftr_out[116]}), .c ({new_AGEMA_signal_8261, mcs1_mcs_mat1_2_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_8740, mcs1_mcs_mat1_2_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_7779, mcs1_mcs_mat1_2_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_9165, mcs1_mcs_mat1_2_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_8263, mcs1_mcs_mat1_2_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_7780, mcs1_mcs_mat1_2_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_8740, mcs1_mcs_mat1_2_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_7414, mcs1_mcs_mat1_2_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_7780, mcs1_mcs_mat1_2_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_7781, mcs1_mcs_mat1_2_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7031, mcs1_mcs_mat1_2_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_8263, mcs1_mcs_mat1_2_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[676]), .c ({new_AGEMA_signal_7781, mcs1_mcs_mat1_2_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[677]), .c ({new_AGEMA_signal_7031, mcs1_mcs_mat1_2_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[678]), .c ({new_AGEMA_signal_7414, mcs1_mcs_mat1_2_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_7782, mcs1_mcs_mat1_2_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_8264, mcs1_mcs_mat1_2_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_7415, mcs1_mcs_mat1_2_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7032, mcs1_mcs_mat1_2_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_7782, mcs1_mcs_mat1_2_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_8265, mcs1_mcs_mat1_2_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_8741, mcs1_mcs_mat1_2_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_7784, mcs1_mcs_mat1_2_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_7032, mcs1_mcs_mat1_2_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_8265, mcs1_mcs_mat1_2_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_8742, mcs1_mcs_mat1_2_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_6617, shiftr_out[84]}), .c ({new_AGEMA_signal_9166, mcs1_mcs_mat1_2_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_7784, mcs1_mcs_mat1_2_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8266, mcs1_mcs_mat1_2_mcs_out[24]}), .c ({new_AGEMA_signal_8742, mcs1_mcs_mat1_2_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_7783, mcs1_mcs_mat1_2_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_7231, shiftr_out[87]}), .c ({new_AGEMA_signal_8266, mcs1_mcs_mat1_2_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_7415, mcs1_mcs_mat1_2_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_6758, mcs1_mcs_mat1_2_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_7783, mcs1_mcs_mat1_2_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[679]), .c ({new_AGEMA_signal_7784, mcs1_mcs_mat1_2_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[680]), .c ({new_AGEMA_signal_7032, mcs1_mcs_mat1_2_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7231, shiftr_out[87]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[681]), .c ({new_AGEMA_signal_7415, mcs1_mcs_mat1_2_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_9694, mcs1_mcs_mat1_2_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_8099, shiftr_out[54]}), .c ({new_AGEMA_signal_9923, mcs1_mcs_mat1_2_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_9452, mcs1_mcs_mat1_2_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8743, mcs1_mcs_mat1_2_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_9694, mcs1_mcs_mat1_2_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_9924, mcs1_mcs_mat1_2_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_9361, shiftr_out[53]}), .c ({new_AGEMA_signal_10139, mcs1_mcs_mat1_2_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_9696, mcs1_mcs_mat1_2_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8743, mcs1_mcs_mat1_2_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_9924, mcs1_mcs_mat1_2_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_10140, mcs1_mcs_mat1_2_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_7619, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_10381, mcs1_mcs_mat1_2_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_9696, mcs1_mcs_mat1_2_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_9925, mcs1_mcs_mat1_2_mcs_out[20]}), .c ({new_AGEMA_signal_10140, mcs1_mcs_mat1_2_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_9695, mcs1_mcs_mat1_2_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_9925, mcs1_mcs_mat1_2_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_9452, mcs1_mcs_mat1_2_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8267, mcs1_mcs_mat1_2_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_9695, mcs1_mcs_mat1_2_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9361, shiftr_out[53]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[682]), .c ({new_AGEMA_signal_9696, mcs1_mcs_mat1_2_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[683]), .c ({new_AGEMA_signal_8743, mcs1_mcs_mat1_2_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[684]), .c ({new_AGEMA_signal_9452, mcs1_mcs_mat1_2_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_7785, mcs1_mcs_mat1_2_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_7788, mcs1_mcs_mat1_2_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_8268, mcs1_mcs_mat1_2_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_8269, mcs1_mcs_mat1_2_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_6759, mcs1_mcs_mat1_2_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_8744, mcs1_mcs_mat1_2_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_8745, mcs1_mcs_mat1_2_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_7033, mcs1_mcs_mat1_2_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_9167, mcs1_mcs_mat1_2_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_6630, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_8269, mcs1_mcs_mat1_2_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_8745, mcs1_mcs_mat1_2_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_7786, mcs1_mcs_mat1_2_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_7310, shiftr_out[21]}), .c ({new_AGEMA_signal_8269, mcs1_mcs_mat1_2_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_7416, mcs1_mcs_mat1_2_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_7417, mcs1_mcs_mat1_2_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_7786, mcs1_mcs_mat1_2_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_7787, mcs1_mcs_mat1_2_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_7033, mcs1_mcs_mat1_2_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_8270, mcs1_mcs_mat1_2_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7310, shiftr_out[21]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[685]), .c ({new_AGEMA_signal_7788, mcs1_mcs_mat1_2_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[686]), .c ({new_AGEMA_signal_7033, mcs1_mcs_mat1_2_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[687]), .c ({new_AGEMA_signal_7417, mcs1_mcs_mat1_2_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_8748, mcs1_mcs_mat1_2_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_7256, mcs1_mcs_mat1_2_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_9168, mcs1_mcs_mat1_2_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_8273, mcs1_mcs_mat1_2_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_8271, mcs1_mcs_mat1_2_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_8746, mcs1_mcs_mat1_2_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_7790, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_7034, mcs1_mcs_mat1_2_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8271, mcs1_mcs_mat1_2_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_7256, mcs1_mcs_mat1_2_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_8272, mcs1_mcs_mat1_2_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_8747, mcs1_mcs_mat1_2_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_7789, mcs1_mcs_mat1_2_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_7790, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_8272, mcs1_mcs_mat1_2_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_6760, mcs1_mcs_mat1_2_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_7034, mcs1_mcs_mat1_2_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_7256, mcs1_mcs_mat1_2_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_9169, mcs1_mcs_mat1_2_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_9453, mcs1_mcs_mat1_2_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_8748, mcs1_mcs_mat1_2_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_7790, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_9169, mcs1_mcs_mat1_2_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_8273, mcs1_mcs_mat1_2_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_8748, mcs1_mcs_mat1_2_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_7789, mcs1_mcs_mat1_2_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_8273, mcs1_mcs_mat1_2_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_6612, shiftr_out[116]}), .b ({new_AGEMA_signal_7418, mcs1_mcs_mat1_2_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_7789, mcs1_mcs_mat1_2_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7292, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[688]), .c ({new_AGEMA_signal_7790, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6680, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[689]), .c ({new_AGEMA_signal_7034, mcs1_mcs_mat1_2_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7226, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[690]), .c ({new_AGEMA_signal_7418, mcs1_mcs_mat1_2_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_7257, mcs1_mcs_mat1_2_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_7231, shiftr_out[87]}), .c ({new_AGEMA_signal_7419, mcs1_mcs_mat1_2_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_8275, mcs1_mcs_mat1_2_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_8749, mcs1_mcs_mat1_2_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_7791, mcs1_mcs_mat1_2_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_8274, mcs1_mcs_mat1_2_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_7420, mcs1_mcs_mat1_2_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_7257, mcs1_mcs_mat1_2_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_7791, mcs1_mcs_mat1_2_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_6761, mcs1_mcs_mat1_2_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_7035, mcs1_mcs_mat1_2_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_7257, mcs1_mcs_mat1_2_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_8750, mcs1_mcs_mat1_2_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_6617, shiftr_out[84]}), .c ({new_AGEMA_signal_9170, mcs1_mcs_mat1_2_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_6761, mcs1_mcs_mat1_2_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8275, mcs1_mcs_mat1_2_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_8750, mcs1_mcs_mat1_2_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_7792, mcs1_mcs_mat1_2_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_7420, mcs1_mcs_mat1_2_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_8275, mcs1_mcs_mat1_2_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7297, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[691]), .c ({new_AGEMA_signal_7792, mcs1_mcs_mat1_2_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6685, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[692]), .c ({new_AGEMA_signal_7035, mcs1_mcs_mat1_2_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7231, shiftr_out[87]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[693]), .c ({new_AGEMA_signal_7420, mcs1_mcs_mat1_2_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_10659, mcs1_mcs_mat1_2_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_9455, mcs1_mcs_mat1_2_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_10893, mcs1_mcs_mat1_2_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_10382, mcs1_mcs_mat1_2_mcs_out[7]}), .b ({new_AGEMA_signal_8099, shiftr_out[54]}), .c ({new_AGEMA_signal_10659, mcs1_mcs_mat1_2_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_10141, mcs1_mcs_mat1_2_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_9361, shiftr_out[53]}), .c ({new_AGEMA_signal_10382, mcs1_mcs_mat1_2_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_9926, mcs1_mcs_mat1_2_mcs_out[6]}), .b ({new_AGEMA_signal_8752, mcs1_mcs_mat1_2_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_10141, mcs1_mcs_mat1_2_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_8751, mcs1_mcs_mat1_2_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_9697, mcs1_mcs_mat1_2_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_9926, mcs1_mcs_mat1_2_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9361, shiftr_out[53]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[694]), .c ({new_AGEMA_signal_9697, mcs1_mcs_mat1_2_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8099, shiftr_out[54]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[695]), .c ({new_AGEMA_signal_8752, mcs1_mcs_mat1_2_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9057, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[696]), .c ({new_AGEMA_signal_9455, mcs1_mcs_mat1_2_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_7421, mcs1_mcs_mat1_2_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_7793, mcs1_mcs_mat1_2_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_8278, mcs1_mcs_mat1_2_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_7310, shiftr_out[21]}), .b ({new_AGEMA_signal_7422, mcs1_mcs_mat1_2_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_7793, mcs1_mcs_mat1_2_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_8279, mcs1_mcs_mat1_2_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_7036, mcs1_mcs_mat1_2_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_8753, mcs1_mcs_mat1_2_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_8280, mcs1_mcs_mat1_2_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_7795, mcs1_mcs_mat1_2_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_8754, mcs1_mcs_mat1_2_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_7796, mcs1_mcs_mat1_2_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_6762, mcs1_mcs_mat1_2_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8280, mcs1_mcs_mat1_2_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7310, shiftr_out[21]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[697]), .c ({new_AGEMA_signal_7796, mcs1_mcs_mat1_2_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6698, shiftr_out[22]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[698]), .c ({new_AGEMA_signal_7036, mcs1_mcs_mat1_2_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7244, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[699]), .c ({new_AGEMA_signal_7422, mcs1_mcs_mat1_2_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U96 ( .a ({new_AGEMA_signal_9456, mcs1_mcs_mat1_3_n128}), .b ({new_AGEMA_signal_10383, mcs1_mcs_mat1_3_n127}), .c ({temp_next_s1[81], temp_next_s0[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U95 ( .a ({new_AGEMA_signal_10164, mcs1_mcs_mat1_3_mcs_out[41]}), .b ({new_AGEMA_signal_7832, mcs1_mcs_mat1_3_mcs_out[45]}), .c ({new_AGEMA_signal_10383, mcs1_mcs_mat1_3_n127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U94 ( .a ({new_AGEMA_signal_7259, mcs1_mcs_mat1_3_mcs_out[33]}), .b ({new_AGEMA_signal_9197, mcs1_mcs_mat1_3_mcs_out[37]}), .c ({new_AGEMA_signal_9456, mcs1_mcs_mat1_3_n128}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U93 ( .a ({new_AGEMA_signal_9698, mcs1_mcs_mat1_3_n126}), .b ({new_AGEMA_signal_10142, mcs1_mcs_mat1_3_n125}), .c ({temp_next_s1[80], temp_next_s0[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U92 ( .a ({new_AGEMA_signal_9947, mcs1_mcs_mat1_3_mcs_out[40]}), .b ({new_AGEMA_signal_9482, mcs1_mcs_mat1_3_mcs_out[44]}), .c ({new_AGEMA_signal_10142, mcs1_mcs_mat1_3_n125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U91 ( .a ({new_AGEMA_signal_9485, mcs1_mcs_mat1_3_mcs_out[32]}), .b ({new_AGEMA_signal_8315, mcs1_mcs_mat1_3_mcs_out[36]}), .c ({new_AGEMA_signal_9698, mcs1_mcs_mat1_3_n126}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U90 ( .a ({new_AGEMA_signal_8755, mcs1_mcs_mat1_3_n124}), .b ({new_AGEMA_signal_10143, mcs1_mcs_mat1_3_n123}), .c ({temp_next_s1[51], temp_next_s0[51]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U89 ( .a ({new_AGEMA_signal_9948, mcs1_mcs_mat1_3_mcs_out[27]}), .b ({new_AGEMA_signal_9199, mcs1_mcs_mat1_3_mcs_out[31]}), .c ({new_AGEMA_signal_10143, mcs1_mcs_mat1_3_n123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U88 ( .a ({new_AGEMA_signal_8325, mcs1_mcs_mat1_3_mcs_out[19]}), .b ({new_AGEMA_signal_8322, mcs1_mcs_mat1_3_mcs_out[23]}), .c ({new_AGEMA_signal_8755, mcs1_mcs_mat1_3_n124}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U87 ( .a ({new_AGEMA_signal_9171, mcs1_mcs_mat1_3_n122}), .b ({new_AGEMA_signal_10386, mcs1_mcs_mat1_3_n121}), .c ({temp_next_s1[50], temp_next_s0[50]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U86 ( .a ({new_AGEMA_signal_10165, mcs1_mcs_mat1_3_mcs_out[26]}), .b ({new_AGEMA_signal_8800, mcs1_mcs_mat1_3_mcs_out[30]}), .c ({new_AGEMA_signal_10386, mcs1_mcs_mat1_3_n121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U85 ( .a ({new_AGEMA_signal_8805, mcs1_mcs_mat1_3_mcs_out[18]}), .b ({new_AGEMA_signal_8803, mcs1_mcs_mat1_3_mcs_out[22]}), .c ({new_AGEMA_signal_9171, mcs1_mcs_mat1_3_n122}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U84 ( .a ({new_AGEMA_signal_9457, mcs1_mcs_mat1_3_n120}), .b ({new_AGEMA_signal_10662, mcs1_mcs_mat1_3_n119}), .c ({temp_next_s1[49], temp_next_s0[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U83 ( .a ({new_AGEMA_signal_10405, mcs1_mcs_mat1_3_mcs_out[25]}), .b ({new_AGEMA_signal_8319, mcs1_mcs_mat1_3_mcs_out[29]}), .c ({new_AGEMA_signal_10662, mcs1_mcs_mat1_3_n119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U82 ( .a ({new_AGEMA_signal_9202, mcs1_mcs_mat1_3_mcs_out[17]}), .b ({new_AGEMA_signal_9201, mcs1_mcs_mat1_3_mcs_out[21]}), .c ({new_AGEMA_signal_9457, mcs1_mcs_mat1_3_n120}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U81 ( .a ({new_AGEMA_signal_8756, mcs1_mcs_mat1_3_n118}), .b ({new_AGEMA_signal_10144, mcs1_mcs_mat1_3_n117}), .c ({temp_next_s1[48], temp_next_s0[48]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U80 ( .a ({new_AGEMA_signal_9950, mcs1_mcs_mat1_3_mcs_out[24]}), .b ({new_AGEMA_signal_9200, mcs1_mcs_mat1_3_mcs_out[28]}), .c ({new_AGEMA_signal_10144, mcs1_mcs_mat1_3_n117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U79 ( .a ({new_AGEMA_signal_8327, mcs1_mcs_mat1_3_mcs_out[16]}), .b ({new_AGEMA_signal_8324, mcs1_mcs_mat1_3_mcs_out[20]}), .c ({new_AGEMA_signal_8756, mcs1_mcs_mat1_3_n118}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U78 ( .a ({new_AGEMA_signal_9699, mcs1_mcs_mat1_3_n116}), .b ({new_AGEMA_signal_9458, mcs1_mcs_mat1_3_n115}), .c ({temp_next_s1[19], temp_next_s0[19]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U77 ( .a ({new_AGEMA_signal_8333, mcs1_mcs_mat1_3_mcs_out[3]}), .b ({new_AGEMA_signal_9206, mcs1_mcs_mat1_3_mcs_out[7]}), .c ({new_AGEMA_signal_9458, mcs1_mcs_mat1_3_n115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U76 ( .a ({new_AGEMA_signal_9488, mcs1_mcs_mat1_3_mcs_out[11]}), .b ({new_AGEMA_signal_9203, mcs1_mcs_mat1_3_mcs_out[15]}), .c ({new_AGEMA_signal_9699, mcs1_mcs_mat1_3_n116}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U75 ( .a ({new_AGEMA_signal_9459, mcs1_mcs_mat1_3_n114}), .b ({new_AGEMA_signal_10663, mcs1_mcs_mat1_3_n113}), .c ({new_AGEMA_signal_10895, mcs_out[243]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U74 ( .a ({new_AGEMA_signal_10400, mcs1_mcs_mat1_3_mcs_out[123]}), .b ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_10663, mcs1_mcs_mat1_3_n113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U73 ( .a ({new_AGEMA_signal_8767, mcs1_mcs_mat1_3_mcs_out[115]}), .b ({new_AGEMA_signal_9177, mcs1_mcs_mat1_3_mcs_out[119]}), .c ({new_AGEMA_signal_9459, mcs1_mcs_mat1_3_n114}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U72 ( .a ({new_AGEMA_signal_9460, mcs1_mcs_mat1_3_n112}), .b ({new_AGEMA_signal_9928, mcs1_mcs_mat1_3_n111}), .c ({new_AGEMA_signal_10145, mcs_out[242]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U71 ( .a ({new_AGEMA_signal_9706, mcs1_mcs_mat1_3_mcs_out[122]}), .b ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_9928, mcs1_mcs_mat1_3_n111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U70 ( .a ({new_AGEMA_signal_8284, mcs1_mcs_mat1_3_mcs_out[114]}), .b ({new_AGEMA_signal_9178, mcs1_mcs_mat1_3_mcs_out[118]}), .c ({new_AGEMA_signal_9460, mcs1_mcs_mat1_3_n112}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U69 ( .a ({new_AGEMA_signal_10388, mcs1_mcs_mat1_3_n110}), .b ({new_AGEMA_signal_8757, mcs1_mcs_mat1_3_n109}), .c ({temp_next_s1[18], temp_next_s0[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U68 ( .a ({new_AGEMA_signal_8334, mcs1_mcs_mat1_3_mcs_out[2]}), .b ({new_AGEMA_signal_8332, mcs1_mcs_mat1_3_mcs_out[6]}), .c ({new_AGEMA_signal_8757, mcs1_mcs_mat1_3_n109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U67 ( .a ({new_AGEMA_signal_10167, mcs1_mcs_mat1_3_mcs_out[10]}), .b ({new_AGEMA_signal_8807, mcs1_mcs_mat1_3_mcs_out[14]}), .c ({new_AGEMA_signal_10388, mcs1_mcs_mat1_3_n110}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U66 ( .a ({new_AGEMA_signal_9172, mcs1_mcs_mat1_3_n108}), .b ({new_AGEMA_signal_10665, mcs1_mcs_mat1_3_n107}), .c ({new_AGEMA_signal_10896, mcs_out[241]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U65 ( .a ({new_AGEMA_signal_10401, mcs1_mcs_mat1_3_mcs_out[121]}), .b ({new_AGEMA_signal_7423, mcs1_mcs_mat1_3_mcs_out[125]}), .c ({new_AGEMA_signal_10665, mcs1_mcs_mat1_3_n107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U64 ( .a ({new_AGEMA_signal_7800, mcs1_mcs_mat1_3_mcs_out[113]}), .b ({new_AGEMA_signal_8766, mcs1_mcs_mat1_3_mcs_out[117]}), .c ({new_AGEMA_signal_9172, mcs1_mcs_mat1_3_n108}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U63 ( .a ({new_AGEMA_signal_9461, mcs1_mcs_mat1_3_n106}), .b ({new_AGEMA_signal_10389, mcs1_mcs_mat1_3_n105}), .c ({new_AGEMA_signal_10666, mcs_out[240]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U62 ( .a ({new_AGEMA_signal_10154, mcs1_mcs_mat1_3_mcs_out[120]}), .b ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_10389, mcs1_mcs_mat1_3_n105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U61 ( .a ({new_AGEMA_signal_9179, mcs1_mcs_mat1_3_mcs_out[112]}), .b ({new_AGEMA_signal_8283, mcs1_mcs_mat1_3_mcs_out[116]}), .c ({new_AGEMA_signal_9461, mcs1_mcs_mat1_3_n106}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U60 ( .a ({new_AGEMA_signal_10390, mcs1_mcs_mat1_3_n104}), .b ({new_AGEMA_signal_9462, mcs1_mcs_mat1_3_n103}), .c ({new_AGEMA_signal_10667, mcs_out[211]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U59 ( .a ({new_AGEMA_signal_9180, mcs1_mcs_mat1_3_mcs_out[111]}), .b ({new_AGEMA_signal_9184, mcs1_mcs_mat1_3_mcs_out[99]}), .c ({new_AGEMA_signal_9462, mcs1_mcs_mat1_3_n103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U58 ( .a ({new_AGEMA_signal_8772, mcs1_mcs_mat1_3_mcs_out[103]}), .b ({new_AGEMA_signal_10155, mcs1_mcs_mat1_3_mcs_out[107]}), .c ({new_AGEMA_signal_10390, mcs1_mcs_mat1_3_n104}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U57 ( .a ({new_AGEMA_signal_10391, mcs1_mcs_mat1_3_n102}), .b ({new_AGEMA_signal_9463, mcs1_mcs_mat1_3_n101}), .c ({new_AGEMA_signal_10668, mcs_out[210]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U56 ( .a ({new_AGEMA_signal_9181, mcs1_mcs_mat1_3_mcs_out[110]}), .b ({new_AGEMA_signal_8293, mcs1_mcs_mat1_3_mcs_out[98]}), .c ({new_AGEMA_signal_9463, mcs1_mcs_mat1_3_n101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U55 ( .a ({new_AGEMA_signal_7805, mcs1_mcs_mat1_3_mcs_out[102]}), .b ({new_AGEMA_signal_10156, mcs1_mcs_mat1_3_mcs_out[106]}), .c ({new_AGEMA_signal_10391, mcs1_mcs_mat1_3_n102}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U54 ( .a ({new_AGEMA_signal_10392, mcs1_mcs_mat1_3_n100}), .b ({new_AGEMA_signal_9464, mcs1_mcs_mat1_3_n99}), .c ({new_AGEMA_signal_10669, mcs_out[209]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U53 ( .a ({new_AGEMA_signal_9182, mcs1_mcs_mat1_3_mcs_out[109]}), .b ({new_AGEMA_signal_7432, mcs1_mcs_mat1_3_mcs_out[97]}), .c ({new_AGEMA_signal_9464, mcs1_mcs_mat1_3_n99}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U52 ( .a ({new_AGEMA_signal_8291, mcs1_mcs_mat1_3_mcs_out[101]}), .b ({new_AGEMA_signal_10157, mcs1_mcs_mat1_3_mcs_out[105]}), .c ({new_AGEMA_signal_10392, mcs1_mcs_mat1_3_n100}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U51 ( .a ({new_AGEMA_signal_10670, mcs1_mcs_mat1_3_n98}), .b ({new_AGEMA_signal_9929, mcs1_mcs_mat1_3_n97}), .c ({new_AGEMA_signal_10897, mcs_out[208]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U50 ( .a ({new_AGEMA_signal_9183, mcs1_mcs_mat1_3_mcs_out[108]}), .b ({new_AGEMA_signal_9710, mcs1_mcs_mat1_3_mcs_out[96]}), .c ({new_AGEMA_signal_9929, mcs1_mcs_mat1_3_n97}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U49 ( .a ({new_AGEMA_signal_8773, mcs1_mcs_mat1_3_mcs_out[100]}), .b ({new_AGEMA_signal_10402, mcs1_mcs_mat1_3_mcs_out[104]}), .c ({new_AGEMA_signal_10670, mcs1_mcs_mat1_3_n98}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U48 ( .a ({new_AGEMA_signal_8758, mcs1_mcs_mat1_3_n96}), .b ({new_AGEMA_signal_9700, mcs1_mcs_mat1_3_n95}), .c ({new_AGEMA_signal_9930, mcs_out[179]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U47 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_8775, mcs1_mcs_mat1_3_mcs_out[95]}), .c ({new_AGEMA_signal_9700, mcs1_mcs_mat1_3_n95}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U46 ( .a ({new_AGEMA_signal_8296, mcs1_mcs_mat1_3_mcs_out[83]}), .b ({new_AGEMA_signal_7813, mcs1_mcs_mat1_3_mcs_out[87]}), .c ({new_AGEMA_signal_8758, mcs1_mcs_mat1_3_n96}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U45 ( .a ({new_AGEMA_signal_8759, mcs1_mcs_mat1_3_n94}), .b ({new_AGEMA_signal_9701, mcs1_mcs_mat1_3_n93}), .c ({new_AGEMA_signal_9931, mcs_out[178]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U43 ( .a ({new_AGEMA_signal_8297, mcs1_mcs_mat1_3_mcs_out[82]}), .b ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_8759, mcs1_mcs_mat1_3_n94}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U42 ( .a ({new_AGEMA_signal_8760, mcs1_mcs_mat1_3_n92}), .b ({new_AGEMA_signal_9702, mcs1_mcs_mat1_3_n91}), .c ({new_AGEMA_signal_9932, mcs_out[177]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U41 ( .a ({new_AGEMA_signal_9478, mcs1_mcs_mat1_3_mcs_out[89]}), .b ({new_AGEMA_signal_7811, mcs1_mcs_mat1_3_mcs_out[93]}), .c ({new_AGEMA_signal_9702, mcs1_mcs_mat1_3_n91}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U40 ( .a ({new_AGEMA_signal_8298, mcs1_mcs_mat1_3_mcs_out[81]}), .b ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_8760, mcs1_mcs_mat1_3_n92}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U39 ( .a ({new_AGEMA_signal_9173, mcs1_mcs_mat1_3_n90}), .b ({new_AGEMA_signal_9465, mcs1_mcs_mat1_3_n89}), .c ({new_AGEMA_signal_9703, mcs_out[176]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U38 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_9185, mcs1_mcs_mat1_3_mcs_out[92]}), .c ({new_AGEMA_signal_9465, mcs1_mcs_mat1_3_n89}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U37 ( .a ({new_AGEMA_signal_8777, mcs1_mcs_mat1_3_mcs_out[80]}), .b ({new_AGEMA_signal_8295, mcs1_mcs_mat1_3_mcs_out[84]}), .c ({new_AGEMA_signal_9173, mcs1_mcs_mat1_3_n90}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U36 ( .a ({new_AGEMA_signal_9174, mcs1_mcs_mat1_3_n88}), .b ({new_AGEMA_signal_10146, mcs1_mcs_mat1_3_n87}), .c ({temp_next_s1[17], temp_next_s0[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U35 ( .a ({new_AGEMA_signal_7455, mcs1_mcs_mat1_3_mcs_out[5]}), .b ({new_AGEMA_signal_9951, mcs1_mcs_mat1_3_mcs_out[9]}), .c ({new_AGEMA_signal_10146, mcs1_mcs_mat1_3_n87}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U34 ( .a ({new_AGEMA_signal_8808, mcs1_mcs_mat1_3_mcs_out[13]}), .b ({new_AGEMA_signal_8812, mcs1_mcs_mat1_3_mcs_out[1]}), .c ({new_AGEMA_signal_9174, mcs1_mcs_mat1_3_n88}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U33 ( .a ({new_AGEMA_signal_9466, mcs1_mcs_mat1_3_n86}), .b ({new_AGEMA_signal_9933, mcs1_mcs_mat1_3_n85}), .c ({new_AGEMA_signal_10147, mcs_out[147]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U32 ( .a ({new_AGEMA_signal_9711, mcs1_mcs_mat1_3_mcs_out[75]}), .b ({new_AGEMA_signal_8778, mcs1_mcs_mat1_3_mcs_out[79]}), .c ({new_AGEMA_signal_9933, mcs1_mcs_mat1_3_n85}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U31 ( .a ({new_AGEMA_signal_9190, mcs1_mcs_mat1_3_mcs_out[67]}), .b ({new_AGEMA_signal_8782, mcs1_mcs_mat1_3_mcs_out[71]}), .c ({new_AGEMA_signal_9466, mcs1_mcs_mat1_3_n86}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U30 ( .a ({new_AGEMA_signal_9467, mcs1_mcs_mat1_3_n84}), .b ({new_AGEMA_signal_10671, mcs1_mcs_mat1_3_n83}), .c ({new_AGEMA_signal_10898, mcs_out[146]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U29 ( .a ({new_AGEMA_signal_10403, mcs1_mcs_mat1_3_mcs_out[74]}), .b ({new_AGEMA_signal_7046, mcs1_mcs_mat1_3_mcs_out[78]}), .c ({new_AGEMA_signal_10671, mcs1_mcs_mat1_3_n83}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U28 ( .a ({new_AGEMA_signal_8785, mcs1_mcs_mat1_3_mcs_out[66]}), .b ({new_AGEMA_signal_9188, mcs1_mcs_mat1_3_mcs_out[70]}), .c ({new_AGEMA_signal_9467, mcs1_mcs_mat1_3_n84}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U27 ( .a ({new_AGEMA_signal_9468, mcs1_mcs_mat1_3_n82}), .b ({new_AGEMA_signal_10148, mcs1_mcs_mat1_3_n81}), .c ({new_AGEMA_signal_10394, mcs_out[145]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U26 ( .a ({new_AGEMA_signal_9939, mcs1_mcs_mat1_3_mcs_out[73]}), .b ({new_AGEMA_signal_7818, mcs1_mcs_mat1_3_mcs_out[77]}), .c ({new_AGEMA_signal_10148, mcs1_mcs_mat1_3_n81}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U25 ( .a ({new_AGEMA_signal_7823, mcs1_mcs_mat1_3_mcs_out[65]}), .b ({new_AGEMA_signal_9189, mcs1_mcs_mat1_3_mcs_out[69]}), .c ({new_AGEMA_signal_9468, mcs1_mcs_mat1_3_n82}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U24 ( .a ({new_AGEMA_signal_9704, mcs1_mcs_mat1_3_n80}), .b ({new_AGEMA_signal_10672, mcs1_mcs_mat1_3_n79}), .c ({new_AGEMA_signal_10899, mcs_out[144]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U23 ( .a ({new_AGEMA_signal_10404, mcs1_mcs_mat1_3_mcs_out[72]}), .b ({new_AGEMA_signal_9186, mcs1_mcs_mat1_3_mcs_out[76]}), .c ({new_AGEMA_signal_10672, mcs1_mcs_mat1_3_n79}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U22 ( .a ({new_AGEMA_signal_9480, mcs1_mcs_mat1_3_mcs_out[64]}), .b ({new_AGEMA_signal_8784, mcs1_mcs_mat1_3_mcs_out[68]}), .c ({new_AGEMA_signal_9704, mcs1_mcs_mat1_3_n80}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U21 ( .a ({new_AGEMA_signal_9175, mcs1_mcs_mat1_3_n78}), .b ({new_AGEMA_signal_10149, mcs1_mcs_mat1_3_n77}), .c ({temp_next_s1[115], temp_next_s0[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U20 ( .a ({new_AGEMA_signal_9941, mcs1_mcs_mat1_3_mcs_out[59]}), .b ({new_AGEMA_signal_8787, mcs1_mcs_mat1_3_mcs_out[63]}), .c ({new_AGEMA_signal_10149, mcs1_mcs_mat1_3_n77}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U19 ( .a ({new_AGEMA_signal_7831, mcs1_mcs_mat1_3_mcs_out[51]}), .b ({new_AGEMA_signal_8792, mcs1_mcs_mat1_3_mcs_out[55]}), .c ({new_AGEMA_signal_9175, mcs1_mcs_mat1_3_n78}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U18 ( .a ({new_AGEMA_signal_9469, mcs1_mcs_mat1_3_n76}), .b ({new_AGEMA_signal_9934, mcs1_mcs_mat1_3_n75}), .c ({temp_next_s1[114], temp_next_s0[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U17 ( .a ({new_AGEMA_signal_9714, mcs1_mcs_mat1_3_mcs_out[58]}), .b ({new_AGEMA_signal_8305, mcs1_mcs_mat1_3_mcs_out[62]}), .c ({new_AGEMA_signal_9934, mcs1_mcs_mat1_3_n75}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U16 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_9193, mcs1_mcs_mat1_3_mcs_out[54]}), .c ({new_AGEMA_signal_9469, mcs1_mcs_mat1_3_n76}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U15 ( .a ({new_AGEMA_signal_9470, mcs1_mcs_mat1_3_n74}), .b ({new_AGEMA_signal_10151, mcs1_mcs_mat1_3_n73}), .c ({temp_next_s1[113], temp_next_s0[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U14 ( .a ({new_AGEMA_signal_9942, mcs1_mcs_mat1_3_mcs_out[57]}), .b ({new_AGEMA_signal_8306, mcs1_mcs_mat1_3_mcs_out[61]}), .c ({new_AGEMA_signal_10151, mcs1_mcs_mat1_3_n73}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U13 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_9194, mcs1_mcs_mat1_3_mcs_out[53]}), .c ({new_AGEMA_signal_9470, mcs1_mcs_mat1_3_n74}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U12 ( .a ({new_AGEMA_signal_9176, mcs1_mcs_mat1_3_n72}), .b ({new_AGEMA_signal_10397, mcs1_mcs_mat1_3_n71}), .c ({temp_next_s1[112], temp_next_s0[112]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U11 ( .a ({new_AGEMA_signal_10161, mcs1_mcs_mat1_3_mcs_out[56]}), .b ({new_AGEMA_signal_9192, mcs1_mcs_mat1_3_mcs_out[60]}), .c ({new_AGEMA_signal_10397, mcs1_mcs_mat1_3_n71}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U10 ( .a ({new_AGEMA_signal_8311, mcs1_mcs_mat1_3_mcs_out[48]}), .b ({new_AGEMA_signal_8794, mcs1_mcs_mat1_3_mcs_out[52]}), .c ({new_AGEMA_signal_9176, mcs1_mcs_mat1_3_n72}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U9 ( .a ({new_AGEMA_signal_9471, mcs1_mcs_mat1_3_n70}), .b ({new_AGEMA_signal_10398, mcs1_mcs_mat1_3_n69}), .c ({temp_next_s1[83], temp_next_s0[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U8 ( .a ({new_AGEMA_signal_10162, mcs1_mcs_mat1_3_mcs_out[43]}), .b ({new_AGEMA_signal_8795, mcs1_mcs_mat1_3_mcs_out[47]}), .c ({new_AGEMA_signal_10398, mcs1_mcs_mat1_3_n69}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U7 ( .a ({new_AGEMA_signal_8798, mcs1_mcs_mat1_3_mcs_out[35]}), .b ({new_AGEMA_signal_9196, mcs1_mcs_mat1_3_mcs_out[39]}), .c ({new_AGEMA_signal_9471, mcs1_mcs_mat1_3_n70}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U6 ( .a ({new_AGEMA_signal_8761, mcs1_mcs_mat1_3_n68}), .b ({new_AGEMA_signal_10399, mcs1_mcs_mat1_3_n67}), .c ({temp_next_s1[82], temp_next_s0[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U5 ( .a ({new_AGEMA_signal_10163, mcs1_mcs_mat1_3_mcs_out[42]}), .b ({new_AGEMA_signal_7444, mcs1_mcs_mat1_3_mcs_out[46]}), .c ({new_AGEMA_signal_10399, mcs1_mcs_mat1_3_n67}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U4 ( .a ({new_AGEMA_signal_8316, mcs1_mcs_mat1_3_mcs_out[34]}), .b ({new_AGEMA_signal_7834, mcs1_mcs_mat1_3_mcs_out[38]}), .c ({new_AGEMA_signal_8761, mcs1_mcs_mat1_3_n68}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U3 ( .a ({new_AGEMA_signal_9705, mcs1_mcs_mat1_3_n66}), .b ({new_AGEMA_signal_10676, mcs1_mcs_mat1_3_n65}), .c ({temp_next_s1[16], temp_next_s0[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U2 ( .a ({new_AGEMA_signal_9726, mcs1_mcs_mat1_3_mcs_out[4]}), .b ({new_AGEMA_signal_10406, mcs1_mcs_mat1_3_mcs_out[8]}), .c ({new_AGEMA_signal_10676, mcs1_mcs_mat1_3_n65}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_U1 ( .a ({new_AGEMA_signal_8813, mcs1_mcs_mat1_3_mcs_out[0]}), .b ({new_AGEMA_signal_9487, mcs1_mcs_mat1_3_mcs_out[12]}), .c ({new_AGEMA_signal_9705, mcs1_mcs_mat1_3_n66}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_10152, mcs1_mcs_mat1_3_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_10400, mcs1_mcs_mat1_3_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_9935, mcs1_mcs_mat1_3_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_8281, mcs1_mcs_mat1_3_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_10152, mcs1_mcs_mat1_3_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_8762, mcs1_mcs_mat1_3_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_9472, mcs1_mcs_mat1_3_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_9706, mcs1_mcs_mat1_3_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_8763, mcs1_mcs_mat1_3_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_9055, shiftr_out[83]}), .c ({new_AGEMA_signal_9472, mcs1_mcs_mat1_3_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_10153, mcs1_mcs_mat1_3_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_9055, shiftr_out[83]}), .c ({new_AGEMA_signal_10401, mcs1_mcs_mat1_3_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_9935, mcs1_mcs_mat1_3_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_10153, mcs1_mcs_mat1_3_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_9707, mcs1_mcs_mat1_3_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9473, mcs1_mcs_mat1_3_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_9935, mcs1_mcs_mat1_3_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_9936, mcs1_mcs_mat1_3_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_10154, mcs1_mcs_mat1_3_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_9707, mcs1_mcs_mat1_3_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_8763, mcs1_mcs_mat1_3_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_9936, mcs1_mcs_mat1_3_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[700]), .c ({new_AGEMA_signal_9707, mcs1_mcs_mat1_3_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[701]), .c ({new_AGEMA_signal_8763, mcs1_mcs_mat1_3_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9055, shiftr_out[83]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[702]), .c ({new_AGEMA_signal_9473, mcs1_mcs_mat1_3_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_8764, mcs1_mcs_mat1_3_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_6691, shiftr_out[50]}), .c ({new_AGEMA_signal_9177, mcs1_mcs_mat1_3_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_8282, mcs1_mcs_mat1_3_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7426, mcs1_mcs_mat1_3_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_8764, mcs1_mcs_mat1_3_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_8765, mcs1_mcs_mat1_3_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_7798, mcs1_mcs_mat1_3_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_9178, mcs1_mcs_mat1_3_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_8282, mcs1_mcs_mat1_3_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7303, shiftr_out[49]}), .c ({new_AGEMA_signal_8765, mcs1_mcs_mat1_3_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_8282, mcs1_mcs_mat1_3_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7797, mcs1_mcs_mat1_3_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_8766, mcs1_mcs_mat1_3_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_7799, mcs1_mcs_mat1_3_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_7037, mcs1_mcs_mat1_3_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_8282, mcs1_mcs_mat1_3_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_7425, mcs1_mcs_mat1_3_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_7798, mcs1_mcs_mat1_3_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_8283, mcs1_mcs_mat1_3_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_6763, mcs1_mcs_mat1_3_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7426, mcs1_mcs_mat1_3_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_7798, mcs1_mcs_mat1_3_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_7037, mcs1_mcs_mat1_3_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_7425, mcs1_mcs_mat1_3_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7303, shiftr_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[703]), .c ({new_AGEMA_signal_7799, mcs1_mcs_mat1_3_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[704]), .c ({new_AGEMA_signal_7037, mcs1_mcs_mat1_3_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[705]), .c ({new_AGEMA_signal_7426, mcs1_mcs_mat1_3_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_8285, mcs1_mcs_mat1_3_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_7038, mcs1_mcs_mat1_3_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_8767, mcs1_mcs_mat1_3_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_7427, mcs1_mcs_mat1_3_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_7428, mcs1_mcs_mat1_3_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_7800, mcs1_mcs_mat1_3_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_8286, mcs1_mcs_mat1_3_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_8768, mcs1_mcs_mat1_3_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_9179, mcs1_mcs_mat1_3_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_8285, mcs1_mcs_mat1_3_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_8768, mcs1_mcs_mat1_3_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_6764, mcs1_mcs_mat1_3_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_7802, mcs1_mcs_mat1_3_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_8285, mcs1_mcs_mat1_3_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_7039, mcs1_mcs_mat1_3_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_7801, mcs1_mcs_mat1_3_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8286, mcs1_mcs_mat1_3_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7309, shiftr_out[17]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[706]), .c ({new_AGEMA_signal_7802, mcs1_mcs_mat1_3_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[707]), .c ({new_AGEMA_signal_7039, mcs1_mcs_mat1_3_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[708]), .c ({new_AGEMA_signal_7428, mcs1_mcs_mat1_3_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({new_AGEMA_signal_8769, mcs1_mcs_mat1_3_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9180, mcs1_mcs_mat1_3_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({new_AGEMA_signal_8770, mcs1_mcs_mat1_3_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9181, mcs1_mcs_mat1_3_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_7429, mcs1_mcs_mat1_3_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_8769, mcs1_mcs_mat1_3_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9182, mcs1_mcs_mat1_3_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_7040, mcs1_mcs_mat1_3_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_8287, mcs1_mcs_mat1_3_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_8769, mcs1_mcs_mat1_3_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_7803, mcs1_mcs_mat1_3_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8770, mcs1_mcs_mat1_3_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9183, mcs1_mcs_mat1_3_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_8288, mcs1_mcs_mat1_3_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_8770, mcs1_mcs_mat1_3_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_7429, mcs1_mcs_mat1_3_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_7804, mcs1_mcs_mat1_3_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_8288, mcs1_mcs_mat1_3_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[709]), .c ({new_AGEMA_signal_7804, mcs1_mcs_mat1_3_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[710]), .c ({new_AGEMA_signal_7040, mcs1_mcs_mat1_3_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[711]), .c ({new_AGEMA_signal_7429, mcs1_mcs_mat1_3_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_9938, mcs1_mcs_mat1_3_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_9937, mcs1_mcs_mat1_3_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_10155, mcs1_mcs_mat1_3_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_9937, mcs1_mcs_mat1_3_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_9474, mcs1_mcs_mat1_3_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_10156, mcs1_mcs_mat1_3_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_8771, mcs1_mcs_mat1_3_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_9055, shiftr_out[83]}), .c ({new_AGEMA_signal_9474, mcs1_mcs_mat1_3_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_9937, mcs1_mcs_mat1_3_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_10157, mcs1_mcs_mat1_3_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_9709, mcs1_mcs_mat1_3_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_8289, mcs1_mcs_mat1_3_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_9937, mcs1_mcs_mat1_3_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_10158, mcs1_mcs_mat1_3_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_10402, mcs1_mcs_mat1_3_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_9938, mcs1_mcs_mat1_3_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_9709, mcs1_mcs_mat1_3_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_10158, mcs1_mcs_mat1_3_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_9708, mcs1_mcs_mat1_3_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_7617, shiftr_out[80]}), .c ({new_AGEMA_signal_9938, mcs1_mcs_mat1_3_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_8771, mcs1_mcs_mat1_3_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_9475, mcs1_mcs_mat1_3_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_9708, mcs1_mcs_mat1_3_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[712]), .c ({new_AGEMA_signal_9709, mcs1_mcs_mat1_3_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[713]), .c ({new_AGEMA_signal_8771, mcs1_mcs_mat1_3_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9055, shiftr_out[83]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[714]), .c ({new_AGEMA_signal_9475, mcs1_mcs_mat1_3_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_7430, mcs1_mcs_mat1_3_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_8290, mcs1_mcs_mat1_3_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_8772, mcs1_mcs_mat1_3_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_7808, mcs1_mcs_mat1_3_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_8290, mcs1_mcs_mat1_3_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_7806, mcs1_mcs_mat1_3_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_7431, mcs1_mcs_mat1_3_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_8291, mcs1_mcs_mat1_3_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_7807, mcs1_mcs_mat1_3_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_8292, mcs1_mcs_mat1_3_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_8773, mcs1_mcs_mat1_3_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_6766, mcs1_mcs_mat1_3_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7808, mcs1_mcs_mat1_3_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_8292, mcs1_mcs_mat1_3_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_7041, mcs1_mcs_mat1_3_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_7303, shiftr_out[49]}), .c ({new_AGEMA_signal_7807, mcs1_mcs_mat1_3_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7303, shiftr_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[715]), .c ({new_AGEMA_signal_7808, mcs1_mcs_mat1_3_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[716]), .c ({new_AGEMA_signal_7041, mcs1_mcs_mat1_3_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[717]), .c ({new_AGEMA_signal_7431, mcs1_mcs_mat1_3_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_9476, mcs1_mcs_mat1_3_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_7433, mcs1_mcs_mat1_3_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_9710, mcs1_mcs_mat1_3_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_9184, mcs1_mcs_mat1_3_mcs_out[99]}), .b ({new_AGEMA_signal_6697, shiftr_out[18]}), .c ({new_AGEMA_signal_9476, mcs1_mcs_mat1_3_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_8774, mcs1_mcs_mat1_3_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_7309, shiftr_out[17]}), .c ({new_AGEMA_signal_9184, mcs1_mcs_mat1_3_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_8293, mcs1_mcs_mat1_3_mcs_out[98]}), .b ({new_AGEMA_signal_7043, mcs1_mcs_mat1_3_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_8774, mcs1_mcs_mat1_3_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_7042, mcs1_mcs_mat1_3_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_7809, mcs1_mcs_mat1_3_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_8293, mcs1_mcs_mat1_3_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7309, shiftr_out[17]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[718]), .c ({new_AGEMA_signal_7809, mcs1_mcs_mat1_3_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[719]), .c ({new_AGEMA_signal_7043, mcs1_mcs_mat1_3_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[720]), .c ({new_AGEMA_signal_7433, mcs1_mcs_mat1_3_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_8294, mcs1_mcs_mat1_3_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_8775, mcs1_mcs_mat1_3_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_7435, mcs1_mcs_mat1_3_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_7436, mcs1_mcs_mat1_3_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_7811, mcs1_mcs_mat1_3_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_8776, mcs1_mcs_mat1_3_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_7044, mcs1_mcs_mat1_3_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_9185, mcs1_mcs_mat1_3_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_8294, mcs1_mcs_mat1_3_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_8776, mcs1_mcs_mat1_3_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_6768, mcs1_mcs_mat1_3_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7812, mcs1_mcs_mat1_3_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_8294, mcs1_mcs_mat1_3_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[721]), .c ({new_AGEMA_signal_7812, mcs1_mcs_mat1_3_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[722]), .c ({new_AGEMA_signal_7044, mcs1_mcs_mat1_3_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[723]), .c ({new_AGEMA_signal_7436, mcs1_mcs_mat1_3_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_7816, mcs1_mcs_mat1_3_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_7817, mcs1_mcs_mat1_3_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_8296, mcs1_mcs_mat1_3_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_7814, mcs1_mcs_mat1_3_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_6769, mcs1_mcs_mat1_3_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_8297, mcs1_mcs_mat1_3_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_7437, mcs1_mcs_mat1_3_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_7814, mcs1_mcs_mat1_3_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_7815, mcs1_mcs_mat1_3_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_8298, mcs1_mcs_mat1_3_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_7045, mcs1_mcs_mat1_3_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_7437, mcs1_mcs_mat1_3_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_7815, mcs1_mcs_mat1_3_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_8299, mcs1_mcs_mat1_3_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_6697, shiftr_out[18]}), .c ({new_AGEMA_signal_8777, mcs1_mcs_mat1_3_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_7816, mcs1_mcs_mat1_3_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_7045, mcs1_mcs_mat1_3_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_8299, mcs1_mcs_mat1_3_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7309, shiftr_out[17]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[724]), .c ({new_AGEMA_signal_7817, mcs1_mcs_mat1_3_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[725]), .c ({new_AGEMA_signal_7045, mcs1_mcs_mat1_3_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[726]), .c ({new_AGEMA_signal_7437, mcs1_mcs_mat1_3_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_8300, mcs1_mcs_mat1_3_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_8778, mcs1_mcs_mat1_3_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_7438, mcs1_mcs_mat1_3_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_7818, mcs1_mcs_mat1_3_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_8779, mcs1_mcs_mat1_3_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_7047, mcs1_mcs_mat1_3_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_9186, mcs1_mcs_mat1_3_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_8300, mcs1_mcs_mat1_3_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_6611, shiftr_out[112]}), .c ({new_AGEMA_signal_8779, mcs1_mcs_mat1_3_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_6770, mcs1_mcs_mat1_3_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7819, mcs1_mcs_mat1_3_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_8300, mcs1_mcs_mat1_3_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[727]), .c ({new_AGEMA_signal_7819, mcs1_mcs_mat1_3_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[728]), .c ({new_AGEMA_signal_7047, mcs1_mcs_mat1_3_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[729]), .c ({new_AGEMA_signal_7438, mcs1_mcs_mat1_3_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_10159, mcs1_mcs_mat1_3_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_10403, mcs1_mcs_mat1_3_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_9940, mcs1_mcs_mat1_3_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9712, mcs1_mcs_mat1_3_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_10159, mcs1_mcs_mat1_3_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_9187, mcs1_mcs_mat1_3_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_9711, mcs1_mcs_mat1_3_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_9712, mcs1_mcs_mat1_3_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_9187, mcs1_mcs_mat1_3_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_9939, mcs1_mcs_mat1_3_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_8780, mcs1_mcs_mat1_3_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_8781, mcs1_mcs_mat1_3_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_9187, mcs1_mcs_mat1_3_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_9479, mcs1_mcs_mat1_3_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_7617, shiftr_out[80]}), .c ({new_AGEMA_signal_9712, mcs1_mcs_mat1_3_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_10160, mcs1_mcs_mat1_3_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_8780, mcs1_mcs_mat1_3_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_10404, mcs1_mcs_mat1_3_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_9940, mcs1_mcs_mat1_3_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9479, mcs1_mcs_mat1_3_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_10160, mcs1_mcs_mat1_3_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_9055, shiftr_out[83]}), .b ({new_AGEMA_signal_9713, mcs1_mcs_mat1_3_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_9940, mcs1_mcs_mat1_3_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[730]), .c ({new_AGEMA_signal_9713, mcs1_mcs_mat1_3_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[731]), .c ({new_AGEMA_signal_8781, mcs1_mcs_mat1_3_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9055, shiftr_out[83]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[732]), .c ({new_AGEMA_signal_9479, mcs1_mcs_mat1_3_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_8302, mcs1_mcs_mat1_3_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_7439, mcs1_mcs_mat1_3_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_8782, mcs1_mcs_mat1_3_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_7821, mcs1_mcs_mat1_3_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_8783, mcs1_mcs_mat1_3_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9188, mcs1_mcs_mat1_3_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_8302, mcs1_mcs_mat1_3_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_8783, mcs1_mcs_mat1_3_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9189, mcs1_mcs_mat1_3_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_7439, mcs1_mcs_mat1_3_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_8303, mcs1_mcs_mat1_3_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_8783, mcs1_mcs_mat1_3_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({new_AGEMA_signal_7048, mcs1_mcs_mat1_3_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_7439, mcs1_mcs_mat1_3_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_7820, mcs1_mcs_mat1_3_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_7303, shiftr_out[49]}), .c ({new_AGEMA_signal_8302, mcs1_mcs_mat1_3_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_7440, mcs1_mcs_mat1_3_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6771, mcs1_mcs_mat1_3_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_7820, mcs1_mcs_mat1_3_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_8303, mcs1_mcs_mat1_3_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_7821, mcs1_mcs_mat1_3_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_8784, mcs1_mcs_mat1_3_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_7440, mcs1_mcs_mat1_3_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_7821, mcs1_mcs_mat1_3_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({new_AGEMA_signal_7822, mcs1_mcs_mat1_3_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_8303, mcs1_mcs_mat1_3_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7303, shiftr_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[733]), .c ({new_AGEMA_signal_7822, mcs1_mcs_mat1_3_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[734]), .c ({new_AGEMA_signal_7048, mcs1_mcs_mat1_3_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[735]), .c ({new_AGEMA_signal_7440, mcs1_mcs_mat1_3_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_8786, mcs1_mcs_mat1_3_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_9190, mcs1_mcs_mat1_3_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({new_AGEMA_signal_8304, mcs1_mcs_mat1_3_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_8785, mcs1_mcs_mat1_3_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_9191, mcs1_mcs_mat1_3_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_7441, mcs1_mcs_mat1_3_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_9480, mcs1_mcs_mat1_3_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_8786, mcs1_mcs_mat1_3_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .c ({new_AGEMA_signal_9191, mcs1_mcs_mat1_3_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_7049, mcs1_mcs_mat1_3_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_8304, mcs1_mcs_mat1_3_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_8786, mcs1_mcs_mat1_3_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_6772, mcs1_mcs_mat1_3_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7824, mcs1_mcs_mat1_3_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_8304, mcs1_mcs_mat1_3_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7309, shiftr_out[17]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[736]), .c ({new_AGEMA_signal_7824, mcs1_mcs_mat1_3_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[737]), .c ({new_AGEMA_signal_7049, mcs1_mcs_mat1_3_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[738]), .c ({new_AGEMA_signal_7441, mcs1_mcs_mat1_3_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_8307, mcs1_mcs_mat1_3_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7442, mcs1_mcs_mat1_3_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_8787, mcs1_mcs_mat1_3_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_7050, mcs1_mcs_mat1_3_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_7825, mcs1_mcs_mat1_3_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8305, mcs1_mcs_mat1_3_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({new_AGEMA_signal_7826, mcs1_mcs_mat1_3_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_8306, mcs1_mcs_mat1_3_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[739]), .c ({new_AGEMA_signal_7826, mcs1_mcs_mat1_3_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[740]), .c ({new_AGEMA_signal_7050, mcs1_mcs_mat1_3_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[741]), .c ({new_AGEMA_signal_7442, mcs1_mcs_mat1_3_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_8790, mcs1_mcs_mat1_3_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_9481, mcs1_mcs_mat1_3_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_9714, mcs1_mcs_mat1_3_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_8791, mcs1_mcs_mat1_3_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_9715, mcs1_mcs_mat1_3_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_9942, mcs1_mcs_mat1_3_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_9943, mcs1_mcs_mat1_3_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_9716, mcs1_mcs_mat1_3_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_10161, mcs1_mcs_mat1_3_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_9717, mcs1_mcs_mat1_3_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_9943, mcs1_mcs_mat1_3_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[742]), .c ({new_AGEMA_signal_9717, mcs1_mcs_mat1_3_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[743]), .c ({new_AGEMA_signal_8791, mcs1_mcs_mat1_3_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9055, shiftr_out[83]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[744]), .c ({new_AGEMA_signal_9481, mcs1_mcs_mat1_3_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_7828, mcs1_mcs_mat1_3_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8309, mcs1_mcs_mat1_3_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_8792, mcs1_mcs_mat1_3_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_8793, mcs1_mcs_mat1_3_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_7827, mcs1_mcs_mat1_3_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_9193, mcs1_mcs_mat1_3_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_7443, mcs1_mcs_mat1_3_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_7827, mcs1_mcs_mat1_3_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({new_AGEMA_signal_8793, mcs1_mcs_mat1_3_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_9194, mcs1_mcs_mat1_3_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_6774, mcs1_mcs_mat1_3_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_8309, mcs1_mcs_mat1_3_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_8793, mcs1_mcs_mat1_3_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_7051, mcs1_mcs_mat1_3_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_7830, mcs1_mcs_mat1_3_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_8309, mcs1_mcs_mat1_3_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_7829, mcs1_mcs_mat1_3_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_8310, mcs1_mcs_mat1_3_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_8794, mcs1_mcs_mat1_3_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_7828, mcs1_mcs_mat1_3_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_7051, mcs1_mcs_mat1_3_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_8310, mcs1_mcs_mat1_3_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_7443, mcs1_mcs_mat1_3_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_7828, mcs1_mcs_mat1_3_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7303, shiftr_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[745]), .c ({new_AGEMA_signal_7830, mcs1_mcs_mat1_3_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[746]), .c ({new_AGEMA_signal_7051, mcs1_mcs_mat1_3_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[747]), .c ({new_AGEMA_signal_7443, mcs1_mcs_mat1_3_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_7445, mcs1_mcs_mat1_3_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_7832, mcs1_mcs_mat1_3_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_9195, mcs1_mcs_mat1_3_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_7052, mcs1_mcs_mat1_3_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_9482, mcs1_mcs_mat1_3_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_8795, mcs1_mcs_mat1_3_mcs_out[47]}), .b ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_9195, mcs1_mcs_mat1_3_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_8312, mcs1_mcs_mat1_3_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_6611, shiftr_out[112]}), .c ({new_AGEMA_signal_8795, mcs1_mcs_mat1_3_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_6775, mcs1_mcs_mat1_3_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_7833, mcs1_mcs_mat1_3_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_8312, mcs1_mcs_mat1_3_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[748]), .c ({new_AGEMA_signal_7833, mcs1_mcs_mat1_3_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[749]), .c ({new_AGEMA_signal_7052, mcs1_mcs_mat1_3_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[750]), .c ({new_AGEMA_signal_7445, mcs1_mcs_mat1_3_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_9944, mcs1_mcs_mat1_3_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_9483, mcs1_mcs_mat1_3_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_10162, mcs1_mcs_mat1_3_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_9718, mcs1_mcs_mat1_3_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8796, mcs1_mcs_mat1_3_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_9944, mcs1_mcs_mat1_3_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_9945, mcs1_mcs_mat1_3_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_9720, mcs1_mcs_mat1_3_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_10163, mcs1_mcs_mat1_3_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_9946, mcs1_mcs_mat1_3_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_8313, mcs1_mcs_mat1_3_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_10164, mcs1_mcs_mat1_3_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_9718, mcs1_mcs_mat1_3_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9484, mcs1_mcs_mat1_3_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_9946, mcs1_mcs_mat1_3_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_9719, mcs1_mcs_mat1_3_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_9484, mcs1_mcs_mat1_3_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_9947, mcs1_mcs_mat1_3_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[751]), .c ({new_AGEMA_signal_9720, mcs1_mcs_mat1_3_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[752]), .c ({new_AGEMA_signal_8796, mcs1_mcs_mat1_3_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9055, shiftr_out[83]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[753]), .c ({new_AGEMA_signal_9484, mcs1_mcs_mat1_3_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_8797, mcs1_mcs_mat1_3_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_6776, mcs1_mcs_mat1_3_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9196, mcs1_mcs_mat1_3_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_7447, mcs1_mcs_mat1_3_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_7446, mcs1_mcs_mat1_3_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_7834, mcs1_mcs_mat1_3_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({new_AGEMA_signal_8797, mcs1_mcs_mat1_3_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_9197, mcs1_mcs_mat1_3_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_7835, mcs1_mcs_mat1_3_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_8314, mcs1_mcs_mat1_3_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_8797, mcs1_mcs_mat1_3_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_7836, mcs1_mcs_mat1_3_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7448, mcs1_mcs_mat1_3_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_8314, mcs1_mcs_mat1_3_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_7836, mcs1_mcs_mat1_3_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7447, mcs1_mcs_mat1_3_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_8315, mcs1_mcs_mat1_3_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_7258, mcs1_mcs_mat1_3_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_7447, mcs1_mcs_mat1_3_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({new_AGEMA_signal_7053, mcs1_mcs_mat1_3_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_7258, mcs1_mcs_mat1_3_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7303, shiftr_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[754]), .c ({new_AGEMA_signal_7836, mcs1_mcs_mat1_3_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[755]), .c ({new_AGEMA_signal_7053, mcs1_mcs_mat1_3_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[756]), .c ({new_AGEMA_signal_7448, mcs1_mcs_mat1_3_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_7837, mcs1_mcs_mat1_3_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7449, mcs1_mcs_mat1_3_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_8316, mcs1_mcs_mat1_3_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_7054, mcs1_mcs_mat1_3_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_7259, mcs1_mcs_mat1_3_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_9198, mcs1_mcs_mat1_3_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_7838, mcs1_mcs_mat1_3_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_9485, mcs1_mcs_mat1_3_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7309, shiftr_out[17]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[757]), .c ({new_AGEMA_signal_7838, mcs1_mcs_mat1_3_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[758]), .c ({new_AGEMA_signal_7054, mcs1_mcs_mat1_3_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[759]), .c ({new_AGEMA_signal_7449, mcs1_mcs_mat1_3_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_8799, mcs1_mcs_mat1_3_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_8318, mcs1_mcs_mat1_3_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_9199, mcs1_mcs_mat1_3_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_7056, mcs1_mcs_mat1_3_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_8319, mcs1_mcs_mat1_3_mcs_out[29]}), .c ({new_AGEMA_signal_8799, mcs1_mcs_mat1_3_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_7055, mcs1_mcs_mat1_3_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_8318, mcs1_mcs_mat1_3_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_8800, mcs1_mcs_mat1_3_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_7841, mcs1_mcs_mat1_3_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_6611, shiftr_out[112]}), .c ({new_AGEMA_signal_8318, mcs1_mcs_mat1_3_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_8801, mcs1_mcs_mat1_3_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_7839, mcs1_mcs_mat1_3_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_9200, mcs1_mcs_mat1_3_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_8320, mcs1_mcs_mat1_3_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_7840, mcs1_mcs_mat1_3_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_8801, mcs1_mcs_mat1_3_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_7450, mcs1_mcs_mat1_3_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_7840, mcs1_mcs_mat1_3_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_7841, mcs1_mcs_mat1_3_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7056, mcs1_mcs_mat1_3_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_8320, mcs1_mcs_mat1_3_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[760]), .c ({new_AGEMA_signal_7841, mcs1_mcs_mat1_3_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[761]), .c ({new_AGEMA_signal_7056, mcs1_mcs_mat1_3_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[762]), .c ({new_AGEMA_signal_7450, mcs1_mcs_mat1_3_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_9721, mcs1_mcs_mat1_3_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_9948, mcs1_mcs_mat1_3_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_9486, mcs1_mcs_mat1_3_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8802, mcs1_mcs_mat1_3_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_9721, mcs1_mcs_mat1_3_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_9949, mcs1_mcs_mat1_3_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_10165, mcs1_mcs_mat1_3_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_9723, mcs1_mcs_mat1_3_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8802, mcs1_mcs_mat1_3_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_9949, mcs1_mcs_mat1_3_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_10166, mcs1_mcs_mat1_3_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_7617, shiftr_out[80]}), .c ({new_AGEMA_signal_10405, mcs1_mcs_mat1_3_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_9723, mcs1_mcs_mat1_3_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_9950, mcs1_mcs_mat1_3_mcs_out[24]}), .c ({new_AGEMA_signal_10166, mcs1_mcs_mat1_3_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_9722, mcs1_mcs_mat1_3_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_9055, shiftr_out[83]}), .c ({new_AGEMA_signal_9950, mcs1_mcs_mat1_3_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_9486, mcs1_mcs_mat1_3_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8321, mcs1_mcs_mat1_3_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_9722, mcs1_mcs_mat1_3_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[763]), .c ({new_AGEMA_signal_9723, mcs1_mcs_mat1_3_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[764]), .c ({new_AGEMA_signal_8802, mcs1_mcs_mat1_3_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9055, shiftr_out[83]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[765]), .c ({new_AGEMA_signal_9486, mcs1_mcs_mat1_3_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_7842, mcs1_mcs_mat1_3_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_6691, shiftr_out[50]}), .c ({new_AGEMA_signal_8322, mcs1_mcs_mat1_3_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_7451, mcs1_mcs_mat1_3_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7057, mcs1_mcs_mat1_3_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_7842, mcs1_mcs_mat1_3_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_8323, mcs1_mcs_mat1_3_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_7303, shiftr_out[49]}), .c ({new_AGEMA_signal_8803, mcs1_mcs_mat1_3_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_7844, mcs1_mcs_mat1_3_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_7057, mcs1_mcs_mat1_3_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_8323, mcs1_mcs_mat1_3_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_8804, mcs1_mcs_mat1_3_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_6623, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_9201, mcs1_mcs_mat1_3_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_7844, mcs1_mcs_mat1_3_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8324, mcs1_mcs_mat1_3_mcs_out[20]}), .c ({new_AGEMA_signal_8804, mcs1_mcs_mat1_3_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_7843, mcs1_mcs_mat1_3_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_8324, mcs1_mcs_mat1_3_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_7451, mcs1_mcs_mat1_3_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_6779, mcs1_mcs_mat1_3_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_7843, mcs1_mcs_mat1_3_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7303, shiftr_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[766]), .c ({new_AGEMA_signal_7844, mcs1_mcs_mat1_3_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[767]), .c ({new_AGEMA_signal_7057, mcs1_mcs_mat1_3_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[768]), .c ({new_AGEMA_signal_7451, mcs1_mcs_mat1_3_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_7845, mcs1_mcs_mat1_3_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_7848, mcs1_mcs_mat1_3_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_8325, mcs1_mcs_mat1_3_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_8326, mcs1_mcs_mat1_3_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_6780, mcs1_mcs_mat1_3_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_8805, mcs1_mcs_mat1_3_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_8806, mcs1_mcs_mat1_3_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_7058, mcs1_mcs_mat1_3_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_9202, mcs1_mcs_mat1_3_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_6629, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_8326, mcs1_mcs_mat1_3_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_8806, mcs1_mcs_mat1_3_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_7846, mcs1_mcs_mat1_3_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_7309, shiftr_out[17]}), .c ({new_AGEMA_signal_8326, mcs1_mcs_mat1_3_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_7452, mcs1_mcs_mat1_3_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_7453, mcs1_mcs_mat1_3_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_7846, mcs1_mcs_mat1_3_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_7847, mcs1_mcs_mat1_3_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_7058, mcs1_mcs_mat1_3_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_8327, mcs1_mcs_mat1_3_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7309, shiftr_out[17]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[769]), .c ({new_AGEMA_signal_7848, mcs1_mcs_mat1_3_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[770]), .c ({new_AGEMA_signal_7058, mcs1_mcs_mat1_3_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[771]), .c ({new_AGEMA_signal_7453, mcs1_mcs_mat1_3_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_8809, mcs1_mcs_mat1_3_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_7260, mcs1_mcs_mat1_3_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_9203, mcs1_mcs_mat1_3_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_8330, mcs1_mcs_mat1_3_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_8328, mcs1_mcs_mat1_3_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_8807, mcs1_mcs_mat1_3_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_7850, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_7059, mcs1_mcs_mat1_3_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8328, mcs1_mcs_mat1_3_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_7260, mcs1_mcs_mat1_3_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_8329, mcs1_mcs_mat1_3_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_8808, mcs1_mcs_mat1_3_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_7849, mcs1_mcs_mat1_3_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_7850, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_8329, mcs1_mcs_mat1_3_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_6781, mcs1_mcs_mat1_3_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_7059, mcs1_mcs_mat1_3_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_7260, mcs1_mcs_mat1_3_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_9204, mcs1_mcs_mat1_3_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_9487, mcs1_mcs_mat1_3_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_8809, mcs1_mcs_mat1_3_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_7850, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_9204, mcs1_mcs_mat1_3_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_8330, mcs1_mcs_mat1_3_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_8809, mcs1_mcs_mat1_3_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_7849, mcs1_mcs_mat1_3_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_8330, mcs1_mcs_mat1_3_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_6611, shiftr_out[112]}), .b ({new_AGEMA_signal_7454, mcs1_mcs_mat1_3_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_7849, mcs1_mcs_mat1_3_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7291, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[772]), .c ({new_AGEMA_signal_7850, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6679, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[773]), .c ({new_AGEMA_signal_7059, mcs1_mcs_mat1_3_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7225, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[774]), .c ({new_AGEMA_signal_7454, mcs1_mcs_mat1_3_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_9205, mcs1_mcs_mat1_3_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_9055, shiftr_out[83]}), .c ({new_AGEMA_signal_9488, mcs1_mcs_mat1_3_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_9952, mcs1_mcs_mat1_3_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_10167, mcs1_mcs_mat1_3_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_9724, mcs1_mcs_mat1_3_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_9951, mcs1_mcs_mat1_3_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_9489, mcs1_mcs_mat1_3_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_9205, mcs1_mcs_mat1_3_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_9724, mcs1_mcs_mat1_3_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_8331, mcs1_mcs_mat1_3_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8810, mcs1_mcs_mat1_3_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_9205, mcs1_mcs_mat1_3_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_10168, mcs1_mcs_mat1_3_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_7617, shiftr_out[80]}), .c ({new_AGEMA_signal_10406, mcs1_mcs_mat1_3_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_8331, mcs1_mcs_mat1_3_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_9952, mcs1_mcs_mat1_3_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_10168, mcs1_mcs_mat1_3_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_9725, mcs1_mcs_mat1_3_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_9489, mcs1_mcs_mat1_3_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_9952, mcs1_mcs_mat1_3_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9359, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[775]), .c ({new_AGEMA_signal_9725, mcs1_mcs_mat1_3_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8097, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[776]), .c ({new_AGEMA_signal_8810, mcs1_mcs_mat1_3_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9055, shiftr_out[83]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[777]), .c ({new_AGEMA_signal_9489, mcs1_mcs_mat1_3_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_9490, mcs1_mcs_mat1_3_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_7456, mcs1_mcs_mat1_3_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_9726, mcs1_mcs_mat1_3_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_9206, mcs1_mcs_mat1_3_mcs_out[7]}), .b ({new_AGEMA_signal_6691, shiftr_out[50]}), .c ({new_AGEMA_signal_9490, mcs1_mcs_mat1_3_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_8811, mcs1_mcs_mat1_3_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_7303, shiftr_out[49]}), .c ({new_AGEMA_signal_9206, mcs1_mcs_mat1_3_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_8332, mcs1_mcs_mat1_3_mcs_out[6]}), .b ({new_AGEMA_signal_7061, mcs1_mcs_mat1_3_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_8811, mcs1_mcs_mat1_3_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_7060, mcs1_mcs_mat1_3_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_7851, mcs1_mcs_mat1_3_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_8332, mcs1_mcs_mat1_3_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7303, shiftr_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[778]), .c ({new_AGEMA_signal_7851, mcs1_mcs_mat1_3_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6691, shiftr_out[50]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[779]), .c ({new_AGEMA_signal_7061, mcs1_mcs_mat1_3_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7237, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[780]), .c ({new_AGEMA_signal_7456, mcs1_mcs_mat1_3_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_7457, mcs1_mcs_mat1_3_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_7852, mcs1_mcs_mat1_3_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_8334, mcs1_mcs_mat1_3_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_7309, shiftr_out[17]}), .b ({new_AGEMA_signal_7458, mcs1_mcs_mat1_3_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_7852, mcs1_mcs_mat1_3_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_8335, mcs1_mcs_mat1_3_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_7062, mcs1_mcs_mat1_3_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_8812, mcs1_mcs_mat1_3_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_8336, mcs1_mcs_mat1_3_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_7854, mcs1_mcs_mat1_3_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_8813, mcs1_mcs_mat1_3_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_7855, mcs1_mcs_mat1_3_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_6783, mcs1_mcs_mat1_3_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8336, mcs1_mcs_mat1_3_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7309, shiftr_out[17]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[781]), .c ({new_AGEMA_signal_7855, mcs1_mcs_mat1_3_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6697, shiftr_out[18]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[782]), .c ({new_AGEMA_signal_7062, mcs1_mcs_mat1_3_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7243, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[783]), .c ({new_AGEMA_signal_7458, mcs1_mcs_mat1_3_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U96 ( .a ({new_AGEMA_signal_9491, mcs1_mcs_mat1_4_n128}), .b ({new_AGEMA_signal_9953, mcs1_mcs_mat1_4_n127}), .c ({temp_next_s1[77], temp_next_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U95 ( .a ({new_AGEMA_signal_8857, mcs1_mcs_mat1_4_mcs_out[41]}), .b ({new_AGEMA_signal_9745, mcs1_mcs_mat1_4_mcs_out[45]}), .c ({new_AGEMA_signal_9953, mcs1_mcs_mat1_4_n127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U94 ( .a ({new_AGEMA_signal_7263, mcs1_mcs_mat1_4_mcs_out[33]}), .b ({new_AGEMA_signal_9231, mcs1_mcs_mat1_4_mcs_out[37]}), .c ({new_AGEMA_signal_9491, mcs1_mcs_mat1_4_n128}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U93 ( .a ({new_AGEMA_signal_9727, mcs1_mcs_mat1_4_n126}), .b ({new_AGEMA_signal_10901, mcs1_mcs_mat1_4_n125}), .c ({temp_next_s1[76], temp_next_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U92 ( .a ({new_AGEMA_signal_8374, mcs1_mcs_mat1_4_mcs_out[40]}), .b ({new_AGEMA_signal_10694, mcs1_mcs_mat1_4_mcs_out[44]}), .c ({new_AGEMA_signal_10901, mcs1_mcs_mat1_4_n125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U91 ( .a ({new_AGEMA_signal_9518, mcs1_mcs_mat1_4_mcs_out[32]}), .b ({new_AGEMA_signal_8376, mcs1_mcs_mat1_4_mcs_out[36]}), .c ({new_AGEMA_signal_9727, mcs1_mcs_mat1_4_n126}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U90 ( .a ({new_AGEMA_signal_8814, mcs1_mcs_mat1_4_n124}), .b ({new_AGEMA_signal_10677, mcs1_mcs_mat1_4_n123}), .c ({temp_next_s1[47], temp_next_s0[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U89 ( .a ({new_AGEMA_signal_8380, mcs1_mcs_mat1_4_mcs_out[27]}), .b ({new_AGEMA_signal_10425, mcs1_mcs_mat1_4_mcs_out[31]}), .c ({new_AGEMA_signal_10677, mcs1_mcs_mat1_4_n123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U88 ( .a ({new_AGEMA_signal_8386, mcs1_mcs_mat1_4_mcs_out[19]}), .b ({new_AGEMA_signal_8383, mcs1_mcs_mat1_4_mcs_out[23]}), .c ({new_AGEMA_signal_8814, mcs1_mcs_mat1_4_n124}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U87 ( .a ({new_AGEMA_signal_9207, mcs1_mcs_mat1_4_n122}), .b ({new_AGEMA_signal_10407, mcs1_mcs_mat1_4_n121}), .c ({temp_next_s1[46], temp_next_s0[46]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U86 ( .a ({new_AGEMA_signal_8862, mcs1_mcs_mat1_4_mcs_out[26]}), .b ({new_AGEMA_signal_10186, mcs1_mcs_mat1_4_mcs_out[30]}), .c ({new_AGEMA_signal_10407, mcs1_mcs_mat1_4_n121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U85 ( .a ({new_AGEMA_signal_8866, mcs1_mcs_mat1_4_mcs_out[18]}), .b ({new_AGEMA_signal_8864, mcs1_mcs_mat1_4_mcs_out[22]}), .c ({new_AGEMA_signal_9207, mcs1_mcs_mat1_4_n122}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U84 ( .a ({new_AGEMA_signal_9492, mcs1_mcs_mat1_4_n120}), .b ({new_AGEMA_signal_10170, mcs1_mcs_mat1_4_n119}), .c ({temp_next_s1[45], temp_next_s0[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U83 ( .a ({new_AGEMA_signal_9233, mcs1_mcs_mat1_4_mcs_out[25]}), .b ({new_AGEMA_signal_9970, mcs1_mcs_mat1_4_mcs_out[29]}), .c ({new_AGEMA_signal_10170, mcs1_mcs_mat1_4_n119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U82 ( .a ({new_AGEMA_signal_9235, mcs1_mcs_mat1_4_mcs_out[17]}), .b ({new_AGEMA_signal_9234, mcs1_mcs_mat1_4_mcs_out[21]}), .c ({new_AGEMA_signal_9492, mcs1_mcs_mat1_4_n120}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U81 ( .a ({new_AGEMA_signal_8815, mcs1_mcs_mat1_4_n118}), .b ({new_AGEMA_signal_10679, mcs1_mcs_mat1_4_n117}), .c ({temp_next_s1[44], temp_next_s0[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U80 ( .a ({new_AGEMA_signal_8382, mcs1_mcs_mat1_4_mcs_out[24]}), .b ({new_AGEMA_signal_10426, mcs1_mcs_mat1_4_mcs_out[28]}), .c ({new_AGEMA_signal_10679, mcs1_mcs_mat1_4_n117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U79 ( .a ({new_AGEMA_signal_8388, mcs1_mcs_mat1_4_mcs_out[16]}), .b ({new_AGEMA_signal_8385, mcs1_mcs_mat1_4_mcs_out[20]}), .c ({new_AGEMA_signal_8815, mcs1_mcs_mat1_4_n118}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U78 ( .a ({new_AGEMA_signal_10680, mcs1_mcs_mat1_4_n116}), .b ({new_AGEMA_signal_9493, mcs1_mcs_mat1_4_n115}), .c ({temp_next_s1[15], temp_next_s0[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U77 ( .a ({new_AGEMA_signal_8393, mcs1_mcs_mat1_4_mcs_out[3]}), .b ({new_AGEMA_signal_9238, mcs1_mcs_mat1_4_mcs_out[7]}), .c ({new_AGEMA_signal_9493, mcs1_mcs_mat1_4_n115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U76 ( .a ({new_AGEMA_signal_7491, mcs1_mcs_mat1_4_mcs_out[11]}), .b ({new_AGEMA_signal_10427, mcs1_mcs_mat1_4_mcs_out[15]}), .c ({new_AGEMA_signal_10680, mcs1_mcs_mat1_4_n116}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U75 ( .a ({new_AGEMA_signal_9495, mcs1_mcs_mat1_4_n114}), .b ({new_AGEMA_signal_9494, mcs1_mcs_mat1_4_n113}), .c ({new_AGEMA_signal_9728, mcs_out[239]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U74 ( .a ({new_AGEMA_signal_9215, mcs1_mcs_mat1_4_mcs_out[123]}), .b ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_9494, mcs1_mcs_mat1_4_n113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U73 ( .a ({new_AGEMA_signal_8828, mcs1_mcs_mat1_4_mcs_out[115]}), .b ({new_AGEMA_signal_9217, mcs1_mcs_mat1_4_mcs_out[119]}), .c ({new_AGEMA_signal_9495, mcs1_mcs_mat1_4_n114}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U72 ( .a ({new_AGEMA_signal_9496, mcs1_mcs_mat1_4_n112}), .b ({new_AGEMA_signal_9729, mcs1_mcs_mat1_4_n111}), .c ({new_AGEMA_signal_9954, mcs_out[238]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U71 ( .a ({new_AGEMA_signal_7856, mcs1_mcs_mat1_4_mcs_out[122]}), .b ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_9729, mcs1_mcs_mat1_4_n111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U70 ( .a ({new_AGEMA_signal_8341, mcs1_mcs_mat1_4_mcs_out[114]}), .b ({new_AGEMA_signal_9218, mcs1_mcs_mat1_4_mcs_out[118]}), .c ({new_AGEMA_signal_9496, mcs1_mcs_mat1_4_n112}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U69 ( .a ({new_AGEMA_signal_10409, mcs1_mcs_mat1_4_n110}), .b ({new_AGEMA_signal_8816, mcs1_mcs_mat1_4_n109}), .c ({temp_next_s1[14], temp_next_s0[14]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U68 ( .a ({new_AGEMA_signal_8394, mcs1_mcs_mat1_4_mcs_out[2]}), .b ({new_AGEMA_signal_8392, mcs1_mcs_mat1_4_mcs_out[6]}), .c ({new_AGEMA_signal_8816, mcs1_mcs_mat1_4_n109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U67 ( .a ({new_AGEMA_signal_8869, mcs1_mcs_mat1_4_mcs_out[10]}), .b ({new_AGEMA_signal_10188, mcs1_mcs_mat1_4_mcs_out[14]}), .c ({new_AGEMA_signal_10409, mcs1_mcs_mat1_4_n110}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U66 ( .a ({new_AGEMA_signal_9208, mcs1_mcs_mat1_4_n108}), .b ({new_AGEMA_signal_9730, mcs1_mcs_mat1_4_n107}), .c ({new_AGEMA_signal_9955, mcs_out[237]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U65 ( .a ({new_AGEMA_signal_9216, mcs1_mcs_mat1_4_mcs_out[121]}), .b ({new_AGEMA_signal_9507, mcs1_mcs_mat1_4_mcs_out[125]}), .c ({new_AGEMA_signal_9730, mcs1_mcs_mat1_4_n107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U64 ( .a ({new_AGEMA_signal_7861, mcs1_mcs_mat1_4_mcs_out[113]}), .b ({new_AGEMA_signal_8827, mcs1_mcs_mat1_4_mcs_out[117]}), .c ({new_AGEMA_signal_9208, mcs1_mcs_mat1_4_n108}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U63 ( .a ({new_AGEMA_signal_9498, mcs1_mcs_mat1_4_n106}), .b ({new_AGEMA_signal_9497, mcs1_mcs_mat1_4_n105}), .c ({new_AGEMA_signal_9731, mcs_out[236]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U62 ( .a ({new_AGEMA_signal_8824, mcs1_mcs_mat1_4_mcs_out[120]}), .b ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_9497, mcs1_mcs_mat1_4_n105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U61 ( .a ({new_AGEMA_signal_9219, mcs1_mcs_mat1_4_mcs_out[112]}), .b ({new_AGEMA_signal_8340, mcs1_mcs_mat1_4_mcs_out[116]}), .c ({new_AGEMA_signal_9498, mcs1_mcs_mat1_4_n106}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U60 ( .a ({new_AGEMA_signal_9209, mcs1_mcs_mat1_4_n104}), .b ({new_AGEMA_signal_10682, mcs1_mcs_mat1_4_n103}), .c ({new_AGEMA_signal_10905, mcs_out[207]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U59 ( .a ({new_AGEMA_signal_10417, mcs1_mcs_mat1_4_mcs_out[111]}), .b ({new_AGEMA_signal_9221, mcs1_mcs_mat1_4_mcs_out[99]}), .c ({new_AGEMA_signal_10682, mcs1_mcs_mat1_4_n103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U58 ( .a ({new_AGEMA_signal_8835, mcs1_mcs_mat1_4_mcs_out[103]}), .b ({new_AGEMA_signal_8831, mcs1_mcs_mat1_4_mcs_out[107]}), .c ({new_AGEMA_signal_9209, mcs1_mcs_mat1_4_n104}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U57 ( .a ({new_AGEMA_signal_9210, mcs1_mcs_mat1_4_n102}), .b ({new_AGEMA_signal_10683, mcs1_mcs_mat1_4_n101}), .c ({new_AGEMA_signal_10906, mcs_out[206]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U56 ( .a ({new_AGEMA_signal_10418, mcs1_mcs_mat1_4_mcs_out[110]}), .b ({new_AGEMA_signal_8350, mcs1_mcs_mat1_4_mcs_out[98]}), .c ({new_AGEMA_signal_10683, mcs1_mcs_mat1_4_n101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U55 ( .a ({new_AGEMA_signal_7866, mcs1_mcs_mat1_4_mcs_out[102]}), .b ({new_AGEMA_signal_8832, mcs1_mcs_mat1_4_mcs_out[106]}), .c ({new_AGEMA_signal_9210, mcs1_mcs_mat1_4_n102}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U54 ( .a ({new_AGEMA_signal_9211, mcs1_mcs_mat1_4_n100}), .b ({new_AGEMA_signal_10684, mcs1_mcs_mat1_4_n99}), .c ({new_AGEMA_signal_10907, mcs_out[205]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U53 ( .a ({new_AGEMA_signal_10419, mcs1_mcs_mat1_4_mcs_out[109]}), .b ({new_AGEMA_signal_7470, mcs1_mcs_mat1_4_mcs_out[97]}), .c ({new_AGEMA_signal_10684, mcs1_mcs_mat1_4_n99}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U52 ( .a ({new_AGEMA_signal_8348, mcs1_mcs_mat1_4_mcs_out[101]}), .b ({new_AGEMA_signal_8833, mcs1_mcs_mat1_4_mcs_out[105]}), .c ({new_AGEMA_signal_9211, mcs1_mcs_mat1_4_n100}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U51 ( .a ({new_AGEMA_signal_9499, mcs1_mcs_mat1_4_n98}), .b ({new_AGEMA_signal_10685, mcs1_mcs_mat1_4_n97}), .c ({new_AGEMA_signal_10908, mcs_out[204]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U50 ( .a ({new_AGEMA_signal_10420, mcs1_mcs_mat1_4_mcs_out[108]}), .b ({new_AGEMA_signal_9737, mcs1_mcs_mat1_4_mcs_out[96]}), .c ({new_AGEMA_signal_10685, mcs1_mcs_mat1_4_n97}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U49 ( .a ({new_AGEMA_signal_8836, mcs1_mcs_mat1_4_mcs_out[100]}), .b ({new_AGEMA_signal_9220, mcs1_mcs_mat1_4_mcs_out[104]}), .c ({new_AGEMA_signal_9499, mcs1_mcs_mat1_4_n98}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U48 ( .a ({new_AGEMA_signal_8817, mcs1_mcs_mat1_4_n96}), .b ({new_AGEMA_signal_10410, mcs1_mcs_mat1_4_n95}), .c ({new_AGEMA_signal_10686, mcs_out[175]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U47 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_10178, mcs1_mcs_mat1_4_mcs_out[95]}), .c ({new_AGEMA_signal_10410, mcs1_mcs_mat1_4_n95}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U46 ( .a ({new_AGEMA_signal_8353, mcs1_mcs_mat1_4_mcs_out[83]}), .b ({new_AGEMA_signal_7871, mcs1_mcs_mat1_4_mcs_out[87]}), .c ({new_AGEMA_signal_8817, mcs1_mcs_mat1_4_n96}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U45 ( .a ({new_AGEMA_signal_8818, mcs1_mcs_mat1_4_n94}), .b ({new_AGEMA_signal_9956, mcs1_mcs_mat1_4_n93}), .c ({new_AGEMA_signal_10171, mcs_out[174]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U43 ( .a ({new_AGEMA_signal_8354, mcs1_mcs_mat1_4_mcs_out[82]}), .b ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_8818, mcs1_mcs_mat1_4_n94}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U42 ( .a ({new_AGEMA_signal_8819, mcs1_mcs_mat1_4_n92}), .b ({new_AGEMA_signal_9957, mcs1_mcs_mat1_4_n91}), .c ({new_AGEMA_signal_10172, mcs_out[173]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U41 ( .a ({new_AGEMA_signal_7473, mcs1_mcs_mat1_4_mcs_out[89]}), .b ({new_AGEMA_signal_9739, mcs1_mcs_mat1_4_mcs_out[93]}), .c ({new_AGEMA_signal_9957, mcs1_mcs_mat1_4_n91}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U40 ( .a ({new_AGEMA_signal_8355, mcs1_mcs_mat1_4_mcs_out[81]}), .b ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_8819, mcs1_mcs_mat1_4_n92}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U39 ( .a ({new_AGEMA_signal_9212, mcs1_mcs_mat1_4_n90}), .b ({new_AGEMA_signal_10687, mcs1_mcs_mat1_4_n89}), .c ({new_AGEMA_signal_10909, mcs_out[172]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U38 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_10421, mcs1_mcs_mat1_4_mcs_out[92]}), .c ({new_AGEMA_signal_10687, mcs1_mcs_mat1_4_n89}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U37 ( .a ({new_AGEMA_signal_8839, mcs1_mcs_mat1_4_mcs_out[80]}), .b ({new_AGEMA_signal_8352, mcs1_mcs_mat1_4_mcs_out[84]}), .c ({new_AGEMA_signal_9212, mcs1_mcs_mat1_4_n90}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U36 ( .a ({new_AGEMA_signal_10411, mcs1_mcs_mat1_4_n88}), .b ({new_AGEMA_signal_8820, mcs1_mcs_mat1_4_n87}), .c ({temp_next_s1[13], temp_next_s0[13]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U35 ( .a ({new_AGEMA_signal_7493, mcs1_mcs_mat1_4_mcs_out[5]}), .b ({new_AGEMA_signal_8390, mcs1_mcs_mat1_4_mcs_out[9]}), .c ({new_AGEMA_signal_8820, mcs1_mcs_mat1_4_n87}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U34 ( .a ({new_AGEMA_signal_10189, mcs1_mcs_mat1_4_mcs_out[13]}), .b ({new_AGEMA_signal_8872, mcs1_mcs_mat1_4_mcs_out[1]}), .c ({new_AGEMA_signal_10411, mcs1_mcs_mat1_4_n88}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U33 ( .a ({new_AGEMA_signal_9500, mcs1_mcs_mat1_4_n86}), .b ({new_AGEMA_signal_10412, mcs1_mcs_mat1_4_n85}), .c ({new_AGEMA_signal_10689, mcs_out[143]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U32 ( .a ({new_AGEMA_signal_7876, mcs1_mcs_mat1_4_mcs_out[75]}), .b ({new_AGEMA_signal_10180, mcs1_mcs_mat1_4_mcs_out[79]}), .c ({new_AGEMA_signal_10412, mcs1_mcs_mat1_4_n85}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U31 ( .a ({new_AGEMA_signal_9226, mcs1_mcs_mat1_4_mcs_out[67]}), .b ({new_AGEMA_signal_8844, mcs1_mcs_mat1_4_mcs_out[71]}), .c ({new_AGEMA_signal_9500, mcs1_mcs_mat1_4_n86}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U30 ( .a ({new_AGEMA_signal_9502, mcs1_mcs_mat1_4_n84}), .b ({new_AGEMA_signal_9501, mcs1_mcs_mat1_4_n83}), .c ({new_AGEMA_signal_9732, mcs_out[142]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U29 ( .a ({new_AGEMA_signal_9222, mcs1_mcs_mat1_4_mcs_out[74]}), .b ({new_AGEMA_signal_8840, mcs1_mcs_mat1_4_mcs_out[78]}), .c ({new_AGEMA_signal_9501, mcs1_mcs_mat1_4_n83}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U28 ( .a ({new_AGEMA_signal_8847, mcs1_mcs_mat1_4_mcs_out[66]}), .b ({new_AGEMA_signal_9224, mcs1_mcs_mat1_4_mcs_out[70]}), .c ({new_AGEMA_signal_9502, mcs1_mcs_mat1_4_n84}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U27 ( .a ({new_AGEMA_signal_9503, mcs1_mcs_mat1_4_n82}), .b ({new_AGEMA_signal_9958, mcs1_mcs_mat1_4_n81}), .c ({new_AGEMA_signal_10173, mcs_out[141]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U26 ( .a ({new_AGEMA_signal_8358, mcs1_mcs_mat1_4_mcs_out[73]}), .b ({new_AGEMA_signal_9741, mcs1_mcs_mat1_4_mcs_out[77]}), .c ({new_AGEMA_signal_9958, mcs1_mcs_mat1_4_n81}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U25 ( .a ({new_AGEMA_signal_7882, mcs1_mcs_mat1_4_mcs_out[65]}), .b ({new_AGEMA_signal_9225, mcs1_mcs_mat1_4_mcs_out[69]}), .c ({new_AGEMA_signal_9503, mcs1_mcs_mat1_4_n82}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U24 ( .a ({new_AGEMA_signal_9733, mcs1_mcs_mat1_4_n80}), .b ({new_AGEMA_signal_10690, mcs1_mcs_mat1_4_n79}), .c ({new_AGEMA_signal_10910, mcs_out[140]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U23 ( .a ({new_AGEMA_signal_9223, mcs1_mcs_mat1_4_mcs_out[72]}), .b ({new_AGEMA_signal_10422, mcs1_mcs_mat1_4_mcs_out[76]}), .c ({new_AGEMA_signal_10690, mcs1_mcs_mat1_4_n79}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U22 ( .a ({new_AGEMA_signal_9514, mcs1_mcs_mat1_4_mcs_out[64]}), .b ({new_AGEMA_signal_8846, mcs1_mcs_mat1_4_mcs_out[68]}), .c ({new_AGEMA_signal_9733, mcs1_mcs_mat1_4_n80}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U21 ( .a ({new_AGEMA_signal_9213, mcs1_mcs_mat1_4_n78}), .b ({new_AGEMA_signal_10413, mcs1_mcs_mat1_4_n77}), .c ({temp_next_s1[111], temp_next_s0[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U20 ( .a ({new_AGEMA_signal_8364, mcs1_mcs_mat1_4_mcs_out[59]}), .b ({new_AGEMA_signal_10182, mcs1_mcs_mat1_4_mcs_out[63]}), .c ({new_AGEMA_signal_10413, mcs1_mcs_mat1_4_n77}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U19 ( .a ({new_AGEMA_signal_7892, mcs1_mcs_mat1_4_mcs_out[51]}), .b ({new_AGEMA_signal_8851, mcs1_mcs_mat1_4_mcs_out[55]}), .c ({new_AGEMA_signal_9213, mcs1_mcs_mat1_4_n78}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U18 ( .a ({new_AGEMA_signal_9504, mcs1_mcs_mat1_4_n76}), .b ({new_AGEMA_signal_10174, mcs1_mcs_mat1_4_n75}), .c ({temp_next_s1[110], temp_next_s0[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U17 ( .a ({new_AGEMA_signal_7884, mcs1_mcs_mat1_4_mcs_out[58]}), .b ({new_AGEMA_signal_9965, mcs1_mcs_mat1_4_mcs_out[62]}), .c ({new_AGEMA_signal_10174, mcs1_mcs_mat1_4_n75}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U16 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_9228, mcs1_mcs_mat1_4_mcs_out[54]}), .c ({new_AGEMA_signal_9504, mcs1_mcs_mat1_4_n76}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U15 ( .a ({new_AGEMA_signal_9505, mcs1_mcs_mat1_4_n74}), .b ({new_AGEMA_signal_10175, mcs1_mcs_mat1_4_n73}), .c ({temp_next_s1[109], temp_next_s0[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U14 ( .a ({new_AGEMA_signal_8365, mcs1_mcs_mat1_4_mcs_out[57]}), .b ({new_AGEMA_signal_9966, mcs1_mcs_mat1_4_mcs_out[61]}), .c ({new_AGEMA_signal_10175, mcs1_mcs_mat1_4_n73}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U13 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_9229, mcs1_mcs_mat1_4_mcs_out[53]}), .c ({new_AGEMA_signal_9505, mcs1_mcs_mat1_4_n74}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U12 ( .a ({new_AGEMA_signal_9214, mcs1_mcs_mat1_4_n72}), .b ({new_AGEMA_signal_10692, mcs1_mcs_mat1_4_n71}), .c ({temp_next_s1[108], temp_next_s0[108]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U11 ( .a ({new_AGEMA_signal_8850, mcs1_mcs_mat1_4_mcs_out[56]}), .b ({new_AGEMA_signal_10423, mcs1_mcs_mat1_4_mcs_out[60]}), .c ({new_AGEMA_signal_10692, mcs1_mcs_mat1_4_n71}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U10 ( .a ({new_AGEMA_signal_8369, mcs1_mcs_mat1_4_mcs_out[48]}), .b ({new_AGEMA_signal_8853, mcs1_mcs_mat1_4_mcs_out[52]}), .c ({new_AGEMA_signal_9214, mcs1_mcs_mat1_4_n72}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U9 ( .a ({new_AGEMA_signal_9506, mcs1_mcs_mat1_4_n70}), .b ({new_AGEMA_signal_10416, mcs1_mcs_mat1_4_n69}), .c ({temp_next_s1[79], temp_next_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U8 ( .a ({new_AGEMA_signal_8855, mcs1_mcs_mat1_4_mcs_out[43]}), .b ({new_AGEMA_signal_10184, mcs1_mcs_mat1_4_mcs_out[47]}), .c ({new_AGEMA_signal_10416, mcs1_mcs_mat1_4_n69}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U7 ( .a ({new_AGEMA_signal_8859, mcs1_mcs_mat1_4_mcs_out[35]}), .b ({new_AGEMA_signal_9230, mcs1_mcs_mat1_4_mcs_out[39]}), .c ({new_AGEMA_signal_9506, mcs1_mcs_mat1_4_n70}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U6 ( .a ({new_AGEMA_signal_8821, mcs1_mcs_mat1_4_n68}), .b ({new_AGEMA_signal_9734, mcs1_mcs_mat1_4_n67}), .c ({temp_next_s1[78], temp_next_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U5 ( .a ({new_AGEMA_signal_8856, mcs1_mcs_mat1_4_mcs_out[42]}), .b ({new_AGEMA_signal_9516, mcs1_mcs_mat1_4_mcs_out[46]}), .c ({new_AGEMA_signal_9734, mcs1_mcs_mat1_4_n67}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U4 ( .a ({new_AGEMA_signal_8377, mcs1_mcs_mat1_4_mcs_out[34]}), .b ({new_AGEMA_signal_7896, mcs1_mcs_mat1_4_mcs_out[38]}), .c ({new_AGEMA_signal_8821, mcs1_mcs_mat1_4_n68}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U3 ( .a ({new_AGEMA_signal_10912, mcs1_mcs_mat1_4_n66}), .b ({new_AGEMA_signal_9960, mcs1_mcs_mat1_4_n65}), .c ({temp_next_s1[12], temp_next_s0[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U2 ( .a ({new_AGEMA_signal_9752, mcs1_mcs_mat1_4_mcs_out[4]}), .b ({new_AGEMA_signal_9237, mcs1_mcs_mat1_4_mcs_out[8]}), .c ({new_AGEMA_signal_9960, mcs1_mcs_mat1_4_n65}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_U1 ( .a ({new_AGEMA_signal_8873, mcs1_mcs_mat1_4_mcs_out[0]}), .b ({new_AGEMA_signal_10695, mcs1_mcs_mat1_4_mcs_out[12]}), .c ({new_AGEMA_signal_10912, mcs1_mcs_mat1_4_n66}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_8822, mcs1_mcs_mat1_4_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_9215, mcs1_mcs_mat1_4_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_8337, mcs1_mcs_mat1_4_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_6784, mcs1_mcs_mat1_4_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8822, mcs1_mcs_mat1_4_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_7063, mcs1_mcs_mat1_4_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_7459, mcs1_mcs_mat1_4_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_7856, mcs1_mcs_mat1_4_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_7064, mcs1_mcs_mat1_4_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_7230, shiftr_out[79]}), .c ({new_AGEMA_signal_7459, mcs1_mcs_mat1_4_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_8823, mcs1_mcs_mat1_4_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_7230, shiftr_out[79]}), .c ({new_AGEMA_signal_9216, mcs1_mcs_mat1_4_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_8337, mcs1_mcs_mat1_4_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_8823, mcs1_mcs_mat1_4_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_7857, mcs1_mcs_mat1_4_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_7460, mcs1_mcs_mat1_4_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_8337, mcs1_mcs_mat1_4_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_8338, mcs1_mcs_mat1_4_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_8824, mcs1_mcs_mat1_4_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_7857, mcs1_mcs_mat1_4_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_7064, mcs1_mcs_mat1_4_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_8338, mcs1_mcs_mat1_4_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[784]), .c ({new_AGEMA_signal_7857, mcs1_mcs_mat1_4_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[785]), .c ({new_AGEMA_signal_7064, mcs1_mcs_mat1_4_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7230, shiftr_out[79]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[786]), .c ({new_AGEMA_signal_7460, mcs1_mcs_mat1_4_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_8825, mcs1_mcs_mat1_4_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_6690, shiftr_out[46]}), .c ({new_AGEMA_signal_9217, mcs1_mcs_mat1_4_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_8339, mcs1_mcs_mat1_4_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7463, mcs1_mcs_mat1_4_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_8825, mcs1_mcs_mat1_4_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_8826, mcs1_mcs_mat1_4_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_7859, mcs1_mcs_mat1_4_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_9218, mcs1_mcs_mat1_4_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_8339, mcs1_mcs_mat1_4_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7302, shiftr_out[45]}), .c ({new_AGEMA_signal_8826, mcs1_mcs_mat1_4_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_8339, mcs1_mcs_mat1_4_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7858, mcs1_mcs_mat1_4_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_8827, mcs1_mcs_mat1_4_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_7860, mcs1_mcs_mat1_4_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_7065, mcs1_mcs_mat1_4_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_8339, mcs1_mcs_mat1_4_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_7462, mcs1_mcs_mat1_4_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_7859, mcs1_mcs_mat1_4_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_8340, mcs1_mcs_mat1_4_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_6785, mcs1_mcs_mat1_4_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7463, mcs1_mcs_mat1_4_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_7859, mcs1_mcs_mat1_4_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_7065, mcs1_mcs_mat1_4_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_7462, mcs1_mcs_mat1_4_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7302, shiftr_out[45]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[787]), .c ({new_AGEMA_signal_7860, mcs1_mcs_mat1_4_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[788]), .c ({new_AGEMA_signal_7065, mcs1_mcs_mat1_4_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[789]), .c ({new_AGEMA_signal_7463, mcs1_mcs_mat1_4_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_8342, mcs1_mcs_mat1_4_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_7066, mcs1_mcs_mat1_4_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_8828, mcs1_mcs_mat1_4_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_7464, mcs1_mcs_mat1_4_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_7465, mcs1_mcs_mat1_4_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_7861, mcs1_mcs_mat1_4_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_8343, mcs1_mcs_mat1_4_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_8829, mcs1_mcs_mat1_4_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_9219, mcs1_mcs_mat1_4_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_8342, mcs1_mcs_mat1_4_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_8829, mcs1_mcs_mat1_4_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_6786, mcs1_mcs_mat1_4_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_7863, mcs1_mcs_mat1_4_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_8342, mcs1_mcs_mat1_4_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_7067, mcs1_mcs_mat1_4_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_7862, mcs1_mcs_mat1_4_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8343, mcs1_mcs_mat1_4_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7308, shiftr_out[13]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[790]), .c ({new_AGEMA_signal_7863, mcs1_mcs_mat1_4_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[791]), .c ({new_AGEMA_signal_7067, mcs1_mcs_mat1_4_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[792]), .c ({new_AGEMA_signal_7465, mcs1_mcs_mat1_4_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({new_AGEMA_signal_10176, mcs1_mcs_mat1_4_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_10417, mcs1_mcs_mat1_4_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({new_AGEMA_signal_10177, mcs1_mcs_mat1_4_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_10418, mcs1_mcs_mat1_4_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_9508, mcs1_mcs_mat1_4_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_10176, mcs1_mcs_mat1_4_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_10419, mcs1_mcs_mat1_4_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_8830, mcs1_mcs_mat1_4_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_9961, mcs1_mcs_mat1_4_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_10176, mcs1_mcs_mat1_4_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_9735, mcs1_mcs_mat1_4_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_10177, mcs1_mcs_mat1_4_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_10420, mcs1_mcs_mat1_4_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_9962, mcs1_mcs_mat1_4_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_10177, mcs1_mcs_mat1_4_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_9508, mcs1_mcs_mat1_4_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_9736, mcs1_mcs_mat1_4_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_9962, mcs1_mcs_mat1_4_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[793]), .c ({new_AGEMA_signal_9736, mcs1_mcs_mat1_4_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[794]), .c ({new_AGEMA_signal_8830, mcs1_mcs_mat1_4_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[795]), .c ({new_AGEMA_signal_9508, mcs1_mcs_mat1_4_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_8346, mcs1_mcs_mat1_4_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_8345, mcs1_mcs_mat1_4_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8831, mcs1_mcs_mat1_4_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_8345, mcs1_mcs_mat1_4_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_7466, mcs1_mcs_mat1_4_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_8832, mcs1_mcs_mat1_4_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_7068, mcs1_mcs_mat1_4_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7230, shiftr_out[79]}), .c ({new_AGEMA_signal_7466, mcs1_mcs_mat1_4_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_8345, mcs1_mcs_mat1_4_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8833, mcs1_mcs_mat1_4_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_7865, mcs1_mcs_mat1_4_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_6787, mcs1_mcs_mat1_4_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_8345, mcs1_mcs_mat1_4_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_8834, mcs1_mcs_mat1_4_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_9220, mcs1_mcs_mat1_4_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_8346, mcs1_mcs_mat1_4_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_7865, mcs1_mcs_mat1_4_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_8834, mcs1_mcs_mat1_4_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_7864, mcs1_mcs_mat1_4_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_6616, shiftr_out[76]}), .c ({new_AGEMA_signal_8346, mcs1_mcs_mat1_4_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_7068, mcs1_mcs_mat1_4_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7467, mcs1_mcs_mat1_4_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_7864, mcs1_mcs_mat1_4_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[796]), .c ({new_AGEMA_signal_7865, mcs1_mcs_mat1_4_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[797]), .c ({new_AGEMA_signal_7068, mcs1_mcs_mat1_4_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7230, shiftr_out[79]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[798]), .c ({new_AGEMA_signal_7467, mcs1_mcs_mat1_4_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_7468, mcs1_mcs_mat1_4_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_8347, mcs1_mcs_mat1_4_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_8835, mcs1_mcs_mat1_4_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_7869, mcs1_mcs_mat1_4_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_8347, mcs1_mcs_mat1_4_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_7867, mcs1_mcs_mat1_4_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_7469, mcs1_mcs_mat1_4_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_8348, mcs1_mcs_mat1_4_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_7868, mcs1_mcs_mat1_4_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_8349, mcs1_mcs_mat1_4_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_8836, mcs1_mcs_mat1_4_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_6788, mcs1_mcs_mat1_4_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7869, mcs1_mcs_mat1_4_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_8349, mcs1_mcs_mat1_4_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_7069, mcs1_mcs_mat1_4_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_7302, shiftr_out[45]}), .c ({new_AGEMA_signal_7868, mcs1_mcs_mat1_4_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7302, shiftr_out[45]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[799]), .c ({new_AGEMA_signal_7869, mcs1_mcs_mat1_4_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[800]), .c ({new_AGEMA_signal_7069, mcs1_mcs_mat1_4_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[801]), .c ({new_AGEMA_signal_7469, mcs1_mcs_mat1_4_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_9509, mcs1_mcs_mat1_4_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_7471, mcs1_mcs_mat1_4_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_9737, mcs1_mcs_mat1_4_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_9221, mcs1_mcs_mat1_4_mcs_out[99]}), .b ({new_AGEMA_signal_6696, shiftr_out[14]}), .c ({new_AGEMA_signal_9509, mcs1_mcs_mat1_4_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_8837, mcs1_mcs_mat1_4_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_7308, shiftr_out[13]}), .c ({new_AGEMA_signal_9221, mcs1_mcs_mat1_4_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_8350, mcs1_mcs_mat1_4_mcs_out[98]}), .b ({new_AGEMA_signal_7071, mcs1_mcs_mat1_4_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_8837, mcs1_mcs_mat1_4_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_7070, mcs1_mcs_mat1_4_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_7870, mcs1_mcs_mat1_4_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_8350, mcs1_mcs_mat1_4_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7308, shiftr_out[13]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[802]), .c ({new_AGEMA_signal_7870, mcs1_mcs_mat1_4_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[803]), .c ({new_AGEMA_signal_7071, mcs1_mcs_mat1_4_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[804]), .c ({new_AGEMA_signal_7471, mcs1_mcs_mat1_4_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_9963, mcs1_mcs_mat1_4_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_10178, mcs1_mcs_mat1_4_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_9511, mcs1_mcs_mat1_4_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_9512, mcs1_mcs_mat1_4_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_9739, mcs1_mcs_mat1_4_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_10179, mcs1_mcs_mat1_4_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_8838, mcs1_mcs_mat1_4_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_10421, mcs1_mcs_mat1_4_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_9963, mcs1_mcs_mat1_4_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_10179, mcs1_mcs_mat1_4_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_8351, mcs1_mcs_mat1_4_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_9740, mcs1_mcs_mat1_4_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_9963, mcs1_mcs_mat1_4_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[805]), .c ({new_AGEMA_signal_9740, mcs1_mcs_mat1_4_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[806]), .c ({new_AGEMA_signal_8838, mcs1_mcs_mat1_4_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[807]), .c ({new_AGEMA_signal_9512, mcs1_mcs_mat1_4_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_7874, mcs1_mcs_mat1_4_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_7875, mcs1_mcs_mat1_4_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_8353, mcs1_mcs_mat1_4_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_7872, mcs1_mcs_mat1_4_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_6790, mcs1_mcs_mat1_4_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_8354, mcs1_mcs_mat1_4_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_7474, mcs1_mcs_mat1_4_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_7872, mcs1_mcs_mat1_4_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_7873, mcs1_mcs_mat1_4_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_8355, mcs1_mcs_mat1_4_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_7072, mcs1_mcs_mat1_4_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_7474, mcs1_mcs_mat1_4_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_7873, mcs1_mcs_mat1_4_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_8356, mcs1_mcs_mat1_4_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_6696, shiftr_out[14]}), .c ({new_AGEMA_signal_8839, mcs1_mcs_mat1_4_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_7874, mcs1_mcs_mat1_4_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_7072, mcs1_mcs_mat1_4_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_8356, mcs1_mcs_mat1_4_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7308, shiftr_out[13]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[808]), .c ({new_AGEMA_signal_7875, mcs1_mcs_mat1_4_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[809]), .c ({new_AGEMA_signal_7072, mcs1_mcs_mat1_4_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[810]), .c ({new_AGEMA_signal_7474, mcs1_mcs_mat1_4_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_9964, mcs1_mcs_mat1_4_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_10180, mcs1_mcs_mat1_4_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_9513, mcs1_mcs_mat1_4_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_9741, mcs1_mcs_mat1_4_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_10181, mcs1_mcs_mat1_4_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_8841, mcs1_mcs_mat1_4_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_10422, mcs1_mcs_mat1_4_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_9964, mcs1_mcs_mat1_4_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7614, shiftr_out[108]}), .c ({new_AGEMA_signal_10181, mcs1_mcs_mat1_4_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_8357, mcs1_mcs_mat1_4_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_9742, mcs1_mcs_mat1_4_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_9964, mcs1_mcs_mat1_4_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[811]), .c ({new_AGEMA_signal_9742, mcs1_mcs_mat1_4_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[812]), .c ({new_AGEMA_signal_8841, mcs1_mcs_mat1_4_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[813]), .c ({new_AGEMA_signal_9513, mcs1_mcs_mat1_4_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_8842, mcs1_mcs_mat1_4_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_9222, mcs1_mcs_mat1_4_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_8359, mcs1_mcs_mat1_4_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7877, mcs1_mcs_mat1_4_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_8842, mcs1_mcs_mat1_4_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_7261, mcs1_mcs_mat1_4_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_7876, mcs1_mcs_mat1_4_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_7877, mcs1_mcs_mat1_4_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_7261, mcs1_mcs_mat1_4_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_8358, mcs1_mcs_mat1_4_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_7073, mcs1_mcs_mat1_4_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_7074, mcs1_mcs_mat1_4_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_7261, mcs1_mcs_mat1_4_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_7475, mcs1_mcs_mat1_4_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_6616, shiftr_out[76]}), .c ({new_AGEMA_signal_7877, mcs1_mcs_mat1_4_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_8843, mcs1_mcs_mat1_4_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_7073, mcs1_mcs_mat1_4_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_9223, mcs1_mcs_mat1_4_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_8359, mcs1_mcs_mat1_4_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7475, mcs1_mcs_mat1_4_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_8843, mcs1_mcs_mat1_4_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_7230, shiftr_out[79]}), .b ({new_AGEMA_signal_7878, mcs1_mcs_mat1_4_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_8359, mcs1_mcs_mat1_4_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[814]), .c ({new_AGEMA_signal_7878, mcs1_mcs_mat1_4_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[815]), .c ({new_AGEMA_signal_7074, mcs1_mcs_mat1_4_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7230, shiftr_out[79]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[816]), .c ({new_AGEMA_signal_7475, mcs1_mcs_mat1_4_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_8360, mcs1_mcs_mat1_4_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_7476, mcs1_mcs_mat1_4_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_8844, mcs1_mcs_mat1_4_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_7880, mcs1_mcs_mat1_4_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_8845, mcs1_mcs_mat1_4_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9224, mcs1_mcs_mat1_4_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_8360, mcs1_mcs_mat1_4_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_8845, mcs1_mcs_mat1_4_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9225, mcs1_mcs_mat1_4_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_7476, mcs1_mcs_mat1_4_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_8361, mcs1_mcs_mat1_4_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_8845, mcs1_mcs_mat1_4_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({new_AGEMA_signal_7075, mcs1_mcs_mat1_4_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_7476, mcs1_mcs_mat1_4_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_7879, mcs1_mcs_mat1_4_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_7302, shiftr_out[45]}), .c ({new_AGEMA_signal_8360, mcs1_mcs_mat1_4_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_7477, mcs1_mcs_mat1_4_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6792, mcs1_mcs_mat1_4_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_7879, mcs1_mcs_mat1_4_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_8361, mcs1_mcs_mat1_4_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_7880, mcs1_mcs_mat1_4_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_8846, mcs1_mcs_mat1_4_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_7477, mcs1_mcs_mat1_4_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_7880, mcs1_mcs_mat1_4_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({new_AGEMA_signal_7881, mcs1_mcs_mat1_4_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_8361, mcs1_mcs_mat1_4_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7302, shiftr_out[45]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[817]), .c ({new_AGEMA_signal_7881, mcs1_mcs_mat1_4_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[818]), .c ({new_AGEMA_signal_7075, mcs1_mcs_mat1_4_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[819]), .c ({new_AGEMA_signal_7477, mcs1_mcs_mat1_4_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_8848, mcs1_mcs_mat1_4_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_9226, mcs1_mcs_mat1_4_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({new_AGEMA_signal_8362, mcs1_mcs_mat1_4_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_8847, mcs1_mcs_mat1_4_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_9227, mcs1_mcs_mat1_4_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_7478, mcs1_mcs_mat1_4_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_9514, mcs1_mcs_mat1_4_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_8848, mcs1_mcs_mat1_4_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .c ({new_AGEMA_signal_9227, mcs1_mcs_mat1_4_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_7076, mcs1_mcs_mat1_4_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_8362, mcs1_mcs_mat1_4_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_8848, mcs1_mcs_mat1_4_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_6793, mcs1_mcs_mat1_4_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7883, mcs1_mcs_mat1_4_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_8362, mcs1_mcs_mat1_4_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7308, shiftr_out[13]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[820]), .c ({new_AGEMA_signal_7883, mcs1_mcs_mat1_4_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[821]), .c ({new_AGEMA_signal_7076, mcs1_mcs_mat1_4_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[822]), .c ({new_AGEMA_signal_7478, mcs1_mcs_mat1_4_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_9967, mcs1_mcs_mat1_4_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_9515, mcs1_mcs_mat1_4_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_10182, mcs1_mcs_mat1_4_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_8849, mcs1_mcs_mat1_4_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_9743, mcs1_mcs_mat1_4_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_9965, mcs1_mcs_mat1_4_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({new_AGEMA_signal_9744, mcs1_mcs_mat1_4_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_9966, mcs1_mcs_mat1_4_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[823]), .c ({new_AGEMA_signal_9744, mcs1_mcs_mat1_4_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[824]), .c ({new_AGEMA_signal_8849, mcs1_mcs_mat1_4_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[825]), .c ({new_AGEMA_signal_9515, mcs1_mcs_mat1_4_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_7078, mcs1_mcs_mat1_4_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_7479, mcs1_mcs_mat1_4_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_7884, mcs1_mcs_mat1_4_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_7079, mcs1_mcs_mat1_4_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_7885, mcs1_mcs_mat1_4_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_8365, mcs1_mcs_mat1_4_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_8366, mcs1_mcs_mat1_4_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_7886, mcs1_mcs_mat1_4_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_8850, mcs1_mcs_mat1_4_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_7887, mcs1_mcs_mat1_4_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_8366, mcs1_mcs_mat1_4_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[826]), .c ({new_AGEMA_signal_7887, mcs1_mcs_mat1_4_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[827]), .c ({new_AGEMA_signal_7079, mcs1_mcs_mat1_4_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7230, shiftr_out[79]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[828]), .c ({new_AGEMA_signal_7479, mcs1_mcs_mat1_4_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_7889, mcs1_mcs_mat1_4_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8367, mcs1_mcs_mat1_4_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_8851, mcs1_mcs_mat1_4_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_8852, mcs1_mcs_mat1_4_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_7888, mcs1_mcs_mat1_4_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_9228, mcs1_mcs_mat1_4_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_7480, mcs1_mcs_mat1_4_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_7888, mcs1_mcs_mat1_4_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({new_AGEMA_signal_8852, mcs1_mcs_mat1_4_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_9229, mcs1_mcs_mat1_4_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_6795, mcs1_mcs_mat1_4_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_8367, mcs1_mcs_mat1_4_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_8852, mcs1_mcs_mat1_4_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_7080, mcs1_mcs_mat1_4_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_7891, mcs1_mcs_mat1_4_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_8367, mcs1_mcs_mat1_4_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_7890, mcs1_mcs_mat1_4_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_8368, mcs1_mcs_mat1_4_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_8853, mcs1_mcs_mat1_4_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_7889, mcs1_mcs_mat1_4_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_7080, mcs1_mcs_mat1_4_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_8368, mcs1_mcs_mat1_4_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_7480, mcs1_mcs_mat1_4_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_7889, mcs1_mcs_mat1_4_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7302, shiftr_out[45]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[829]), .c ({new_AGEMA_signal_7891, mcs1_mcs_mat1_4_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[830]), .c ({new_AGEMA_signal_7080, mcs1_mcs_mat1_4_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[831]), .c ({new_AGEMA_signal_7480, mcs1_mcs_mat1_4_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_9517, mcs1_mcs_mat1_4_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_9745, mcs1_mcs_mat1_4_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_8854, mcs1_mcs_mat1_4_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_10694, mcs1_mcs_mat1_4_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_10184, mcs1_mcs_mat1_4_mcs_out[47]}), .b ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_9968, mcs1_mcs_mat1_4_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_7614, shiftr_out[108]}), .c ({new_AGEMA_signal_10184, mcs1_mcs_mat1_4_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_8370, mcs1_mcs_mat1_4_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_9746, mcs1_mcs_mat1_4_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_9968, mcs1_mcs_mat1_4_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[832]), .c ({new_AGEMA_signal_9746, mcs1_mcs_mat1_4_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[833]), .c ({new_AGEMA_signal_8854, mcs1_mcs_mat1_4_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[834]), .c ({new_AGEMA_signal_9517, mcs1_mcs_mat1_4_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_8371, mcs1_mcs_mat1_4_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_7481, mcs1_mcs_mat1_4_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_8855, mcs1_mcs_mat1_4_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_7893, mcs1_mcs_mat1_4_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7081, mcs1_mcs_mat1_4_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_8371, mcs1_mcs_mat1_4_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_8372, mcs1_mcs_mat1_4_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_7895, mcs1_mcs_mat1_4_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_8856, mcs1_mcs_mat1_4_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_8373, mcs1_mcs_mat1_4_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_6796, mcs1_mcs_mat1_4_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_8857, mcs1_mcs_mat1_4_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_7893, mcs1_mcs_mat1_4_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7482, mcs1_mcs_mat1_4_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8373, mcs1_mcs_mat1_4_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_7894, mcs1_mcs_mat1_4_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_7482, mcs1_mcs_mat1_4_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8374, mcs1_mcs_mat1_4_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[835]), .c ({new_AGEMA_signal_7895, mcs1_mcs_mat1_4_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[836]), .c ({new_AGEMA_signal_7081, mcs1_mcs_mat1_4_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7230, shiftr_out[79]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[837]), .c ({new_AGEMA_signal_7482, mcs1_mcs_mat1_4_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_8858, mcs1_mcs_mat1_4_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_6797, mcs1_mcs_mat1_4_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9230, mcs1_mcs_mat1_4_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_7484, mcs1_mcs_mat1_4_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_7483, mcs1_mcs_mat1_4_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_7896, mcs1_mcs_mat1_4_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({new_AGEMA_signal_8858, mcs1_mcs_mat1_4_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_9231, mcs1_mcs_mat1_4_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_7897, mcs1_mcs_mat1_4_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_8375, mcs1_mcs_mat1_4_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_8858, mcs1_mcs_mat1_4_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_7898, mcs1_mcs_mat1_4_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7485, mcs1_mcs_mat1_4_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_8375, mcs1_mcs_mat1_4_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_7898, mcs1_mcs_mat1_4_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7484, mcs1_mcs_mat1_4_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_8376, mcs1_mcs_mat1_4_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_7262, mcs1_mcs_mat1_4_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_7484, mcs1_mcs_mat1_4_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({new_AGEMA_signal_7082, mcs1_mcs_mat1_4_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_7262, mcs1_mcs_mat1_4_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7302, shiftr_out[45]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[838]), .c ({new_AGEMA_signal_7898, mcs1_mcs_mat1_4_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[839]), .c ({new_AGEMA_signal_7082, mcs1_mcs_mat1_4_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[840]), .c ({new_AGEMA_signal_7485, mcs1_mcs_mat1_4_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_7899, mcs1_mcs_mat1_4_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7486, mcs1_mcs_mat1_4_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_8377, mcs1_mcs_mat1_4_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_7083, mcs1_mcs_mat1_4_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_7263, mcs1_mcs_mat1_4_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_9232, mcs1_mcs_mat1_4_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_7900, mcs1_mcs_mat1_4_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_9518, mcs1_mcs_mat1_4_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7308, shiftr_out[13]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[841]), .c ({new_AGEMA_signal_7900, mcs1_mcs_mat1_4_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[842]), .c ({new_AGEMA_signal_7083, mcs1_mcs_mat1_4_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[843]), .c ({new_AGEMA_signal_7486, mcs1_mcs_mat1_4_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_10185, mcs1_mcs_mat1_4_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_9969, mcs1_mcs_mat1_4_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_10425, mcs1_mcs_mat1_4_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_8861, mcs1_mcs_mat1_4_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_9970, mcs1_mcs_mat1_4_mcs_out[29]}), .c ({new_AGEMA_signal_10185, mcs1_mcs_mat1_4_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_9969, mcs1_mcs_mat1_4_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_10186, mcs1_mcs_mat1_4_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_9749, mcs1_mcs_mat1_4_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7614, shiftr_out[108]}), .c ({new_AGEMA_signal_9969, mcs1_mcs_mat1_4_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_10187, mcs1_mcs_mat1_4_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_9747, mcs1_mcs_mat1_4_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_10426, mcs1_mcs_mat1_4_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_9971, mcs1_mcs_mat1_4_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_9748, mcs1_mcs_mat1_4_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_10187, mcs1_mcs_mat1_4_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_9519, mcs1_mcs_mat1_4_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_9748, mcs1_mcs_mat1_4_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_9749, mcs1_mcs_mat1_4_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8861, mcs1_mcs_mat1_4_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_9971, mcs1_mcs_mat1_4_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[844]), .c ({new_AGEMA_signal_9749, mcs1_mcs_mat1_4_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[845]), .c ({new_AGEMA_signal_8861, mcs1_mcs_mat1_4_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[846]), .c ({new_AGEMA_signal_9519, mcs1_mcs_mat1_4_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_7901, mcs1_mcs_mat1_4_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_8380, mcs1_mcs_mat1_4_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_7487, mcs1_mcs_mat1_4_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7084, mcs1_mcs_mat1_4_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_7901, mcs1_mcs_mat1_4_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_8381, mcs1_mcs_mat1_4_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_8862, mcs1_mcs_mat1_4_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_7903, mcs1_mcs_mat1_4_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_7084, mcs1_mcs_mat1_4_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_8381, mcs1_mcs_mat1_4_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_8863, mcs1_mcs_mat1_4_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_6616, shiftr_out[76]}), .c ({new_AGEMA_signal_9233, mcs1_mcs_mat1_4_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_7903, mcs1_mcs_mat1_4_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8382, mcs1_mcs_mat1_4_mcs_out[24]}), .c ({new_AGEMA_signal_8863, mcs1_mcs_mat1_4_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_7902, mcs1_mcs_mat1_4_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_7230, shiftr_out[79]}), .c ({new_AGEMA_signal_8382, mcs1_mcs_mat1_4_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_7487, mcs1_mcs_mat1_4_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_6799, mcs1_mcs_mat1_4_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_7902, mcs1_mcs_mat1_4_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[847]), .c ({new_AGEMA_signal_7903, mcs1_mcs_mat1_4_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[848]), .c ({new_AGEMA_signal_7084, mcs1_mcs_mat1_4_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7230, shiftr_out[79]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[849]), .c ({new_AGEMA_signal_7487, mcs1_mcs_mat1_4_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_7904, mcs1_mcs_mat1_4_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_6690, shiftr_out[46]}), .c ({new_AGEMA_signal_8383, mcs1_mcs_mat1_4_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_7488, mcs1_mcs_mat1_4_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7085, mcs1_mcs_mat1_4_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_7904, mcs1_mcs_mat1_4_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_8384, mcs1_mcs_mat1_4_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_7302, shiftr_out[45]}), .c ({new_AGEMA_signal_8864, mcs1_mcs_mat1_4_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_7906, mcs1_mcs_mat1_4_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_7085, mcs1_mcs_mat1_4_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_8384, mcs1_mcs_mat1_4_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_8865, mcs1_mcs_mat1_4_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_6622, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_9234, mcs1_mcs_mat1_4_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_7906, mcs1_mcs_mat1_4_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8385, mcs1_mcs_mat1_4_mcs_out[20]}), .c ({new_AGEMA_signal_8865, mcs1_mcs_mat1_4_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_7905, mcs1_mcs_mat1_4_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_8385, mcs1_mcs_mat1_4_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_7488, mcs1_mcs_mat1_4_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_6800, mcs1_mcs_mat1_4_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_7905, mcs1_mcs_mat1_4_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7302, shiftr_out[45]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[850]), .c ({new_AGEMA_signal_7906, mcs1_mcs_mat1_4_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[851]), .c ({new_AGEMA_signal_7085, mcs1_mcs_mat1_4_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[852]), .c ({new_AGEMA_signal_7488, mcs1_mcs_mat1_4_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_7907, mcs1_mcs_mat1_4_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_7910, mcs1_mcs_mat1_4_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_8386, mcs1_mcs_mat1_4_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_8387, mcs1_mcs_mat1_4_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_6801, mcs1_mcs_mat1_4_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_8866, mcs1_mcs_mat1_4_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_8867, mcs1_mcs_mat1_4_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_7086, mcs1_mcs_mat1_4_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_9235, mcs1_mcs_mat1_4_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_6628, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_8387, mcs1_mcs_mat1_4_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_8867, mcs1_mcs_mat1_4_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_7908, mcs1_mcs_mat1_4_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_7308, shiftr_out[13]}), .c ({new_AGEMA_signal_8387, mcs1_mcs_mat1_4_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_7489, mcs1_mcs_mat1_4_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_7490, mcs1_mcs_mat1_4_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_7908, mcs1_mcs_mat1_4_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_7909, mcs1_mcs_mat1_4_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_7086, mcs1_mcs_mat1_4_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_8388, mcs1_mcs_mat1_4_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7308, shiftr_out[13]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[853]), .c ({new_AGEMA_signal_7910, mcs1_mcs_mat1_4_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[854]), .c ({new_AGEMA_signal_7086, mcs1_mcs_mat1_4_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[855]), .c ({new_AGEMA_signal_7490, mcs1_mcs_mat1_4_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_10190, mcs1_mcs_mat1_4_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_9236, mcs1_mcs_mat1_4_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_10427, mcs1_mcs_mat1_4_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_9974, mcs1_mcs_mat1_4_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_9972, mcs1_mcs_mat1_4_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_10188, mcs1_mcs_mat1_4_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_9751, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_8868, mcs1_mcs_mat1_4_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_9972, mcs1_mcs_mat1_4_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_9236, mcs1_mcs_mat1_4_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_9973, mcs1_mcs_mat1_4_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_10189, mcs1_mcs_mat1_4_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_9750, mcs1_mcs_mat1_4_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_9751, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_9973, mcs1_mcs_mat1_4_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_8389, mcs1_mcs_mat1_4_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_8868, mcs1_mcs_mat1_4_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_9236, mcs1_mcs_mat1_4_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_10428, mcs1_mcs_mat1_4_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_10695, mcs1_mcs_mat1_4_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_10190, mcs1_mcs_mat1_4_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_9751, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_10428, mcs1_mcs_mat1_4_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_9974, mcs1_mcs_mat1_4_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_10190, mcs1_mcs_mat1_4_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_9750, mcs1_mcs_mat1_4_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_9974, mcs1_mcs_mat1_4_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_7614, shiftr_out[108]}), .b ({new_AGEMA_signal_9520, mcs1_mcs_mat1_4_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_9750, mcs1_mcs_mat1_4_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9356, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[856]), .c ({new_AGEMA_signal_9751, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8094, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[857]), .c ({new_AGEMA_signal_8868, mcs1_mcs_mat1_4_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9052, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[858]), .c ({new_AGEMA_signal_9520, mcs1_mcs_mat1_4_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_7264, mcs1_mcs_mat1_4_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_7230, shiftr_out[79]}), .c ({new_AGEMA_signal_7491, mcs1_mcs_mat1_4_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_8391, mcs1_mcs_mat1_4_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_8869, mcs1_mcs_mat1_4_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_7911, mcs1_mcs_mat1_4_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_8390, mcs1_mcs_mat1_4_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_7492, mcs1_mcs_mat1_4_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_7264, mcs1_mcs_mat1_4_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_7911, mcs1_mcs_mat1_4_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_6802, mcs1_mcs_mat1_4_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_7087, mcs1_mcs_mat1_4_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_7264, mcs1_mcs_mat1_4_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_8870, mcs1_mcs_mat1_4_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_6616, shiftr_out[76]}), .c ({new_AGEMA_signal_9237, mcs1_mcs_mat1_4_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_6802, mcs1_mcs_mat1_4_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8391, mcs1_mcs_mat1_4_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_8870, mcs1_mcs_mat1_4_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_7912, mcs1_mcs_mat1_4_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_7492, mcs1_mcs_mat1_4_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_8391, mcs1_mcs_mat1_4_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7296, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[859]), .c ({new_AGEMA_signal_7912, mcs1_mcs_mat1_4_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6684, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[860]), .c ({new_AGEMA_signal_7087, mcs1_mcs_mat1_4_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7230, shiftr_out[79]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[861]), .c ({new_AGEMA_signal_7492, mcs1_mcs_mat1_4_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_9521, mcs1_mcs_mat1_4_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_7494, mcs1_mcs_mat1_4_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_9752, mcs1_mcs_mat1_4_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_9238, mcs1_mcs_mat1_4_mcs_out[7]}), .b ({new_AGEMA_signal_6690, shiftr_out[46]}), .c ({new_AGEMA_signal_9521, mcs1_mcs_mat1_4_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_8871, mcs1_mcs_mat1_4_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_7302, shiftr_out[45]}), .c ({new_AGEMA_signal_9238, mcs1_mcs_mat1_4_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_8392, mcs1_mcs_mat1_4_mcs_out[6]}), .b ({new_AGEMA_signal_7089, mcs1_mcs_mat1_4_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_8871, mcs1_mcs_mat1_4_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_7088, mcs1_mcs_mat1_4_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_7913, mcs1_mcs_mat1_4_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_8392, mcs1_mcs_mat1_4_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7302, shiftr_out[45]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[862]), .c ({new_AGEMA_signal_7913, mcs1_mcs_mat1_4_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6690, shiftr_out[46]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[863]), .c ({new_AGEMA_signal_7089, mcs1_mcs_mat1_4_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7236, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[864]), .c ({new_AGEMA_signal_7494, mcs1_mcs_mat1_4_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_7495, mcs1_mcs_mat1_4_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_7914, mcs1_mcs_mat1_4_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_8394, mcs1_mcs_mat1_4_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_7308, shiftr_out[13]}), .b ({new_AGEMA_signal_7496, mcs1_mcs_mat1_4_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_7914, mcs1_mcs_mat1_4_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_8395, mcs1_mcs_mat1_4_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_7090, mcs1_mcs_mat1_4_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_8872, mcs1_mcs_mat1_4_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_8396, mcs1_mcs_mat1_4_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_7916, mcs1_mcs_mat1_4_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_8873, mcs1_mcs_mat1_4_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_7917, mcs1_mcs_mat1_4_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_6804, mcs1_mcs_mat1_4_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8396, mcs1_mcs_mat1_4_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7308, shiftr_out[13]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[865]), .c ({new_AGEMA_signal_7917, mcs1_mcs_mat1_4_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6696, shiftr_out[14]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[866]), .c ({new_AGEMA_signal_7090, mcs1_mcs_mat1_4_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7242, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[867]), .c ({new_AGEMA_signal_7496, mcs1_mcs_mat1_4_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U96 ( .a ({new_AGEMA_signal_9522, mcs1_mcs_mat1_5_n128}), .b ({new_AGEMA_signal_9239, mcs1_mcs_mat1_5_n127}), .c ({temp_next_s1[73], temp_next_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U95 ( .a ({new_AGEMA_signal_8916, mcs1_mcs_mat1_5_mcs_out[41]}), .b ({new_AGEMA_signal_7953, mcs1_mcs_mat1_5_mcs_out[45]}), .c ({new_AGEMA_signal_9239, mcs1_mcs_mat1_5_n127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U94 ( .a ({new_AGEMA_signal_9272, mcs1_mcs_mat1_5_mcs_out[33]}), .b ({new_AGEMA_signal_9271, mcs1_mcs_mat1_5_mcs_out[37]}), .c ({new_AGEMA_signal_9522, mcs1_mcs_mat1_5_n128}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U93 ( .a ({new_AGEMA_signal_10913, mcs1_mcs_mat1_5_n126}), .b ({new_AGEMA_signal_9754, mcs1_mcs_mat1_5_n125}), .c ({temp_next_s1[72], temp_next_s0[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U92 ( .a ({new_AGEMA_signal_8434, mcs1_mcs_mat1_5_mcs_out[40]}), .b ({new_AGEMA_signal_9542, mcs1_mcs_mat1_5_mcs_out[44]}), .c ({new_AGEMA_signal_9754, mcs1_mcs_mat1_5_n125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U91 ( .a ({new_AGEMA_signal_10709, mcs1_mcs_mat1_5_mcs_out[32]}), .b ({new_AGEMA_signal_8436, mcs1_mcs_mat1_5_mcs_out[36]}), .c ({new_AGEMA_signal_10913, mcs1_mcs_mat1_5_n126}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U90 ( .a ({new_AGEMA_signal_10191, mcs1_mcs_mat1_5_n124}), .b ({new_AGEMA_signal_9523, mcs1_mcs_mat1_5_n123}), .c ({temp_next_s1[43], temp_next_s0[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U89 ( .a ({new_AGEMA_signal_8441, mcs1_mcs_mat1_5_mcs_out[27]}), .b ({new_AGEMA_signal_9273, mcs1_mcs_mat1_5_mcs_out[31]}), .c ({new_AGEMA_signal_9523, mcs1_mcs_mat1_5_n123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U88 ( .a ({new_AGEMA_signal_9992, mcs1_mcs_mat1_5_mcs_out[19]}), .b ({new_AGEMA_signal_8444, mcs1_mcs_mat1_5_mcs_out[23]}), .c ({new_AGEMA_signal_10191, mcs1_mcs_mat1_5_n124}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U87 ( .a ({new_AGEMA_signal_10430, mcs1_mcs_mat1_5_n122}), .b ({new_AGEMA_signal_9240, mcs1_mcs_mat1_5_n121}), .c ({temp_next_s1[42], temp_next_s0[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U86 ( .a ({new_AGEMA_signal_8922, mcs1_mcs_mat1_5_mcs_out[26]}), .b ({new_AGEMA_signal_8920, mcs1_mcs_mat1_5_mcs_out[30]}), .c ({new_AGEMA_signal_9240, mcs1_mcs_mat1_5_n121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U85 ( .a ({new_AGEMA_signal_10212, mcs1_mcs_mat1_5_mcs_out[18]}), .b ({new_AGEMA_signal_8924, mcs1_mcs_mat1_5_mcs_out[22]}), .c ({new_AGEMA_signal_10430, mcs1_mcs_mat1_5_n122}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U84 ( .a ({new_AGEMA_signal_10697, mcs1_mcs_mat1_5_n120}), .b ({new_AGEMA_signal_9524, mcs1_mcs_mat1_5_n119}), .c ({temp_next_s1[41], temp_next_s0[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U83 ( .a ({new_AGEMA_signal_9275, mcs1_mcs_mat1_5_mcs_out[25]}), .b ({new_AGEMA_signal_8439, mcs1_mcs_mat1_5_mcs_out[29]}), .c ({new_AGEMA_signal_9524, mcs1_mcs_mat1_5_n119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U82 ( .a ({new_AGEMA_signal_10452, mcs1_mcs_mat1_5_mcs_out[17]}), .b ({new_AGEMA_signal_9276, mcs1_mcs_mat1_5_mcs_out[21]}), .c ({new_AGEMA_signal_10697, mcs1_mcs_mat1_5_n120}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U81 ( .a ({new_AGEMA_signal_10192, mcs1_mcs_mat1_5_n118}), .b ({new_AGEMA_signal_9525, mcs1_mcs_mat1_5_n117}), .c ({temp_next_s1[40], temp_next_s0[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U80 ( .a ({new_AGEMA_signal_8443, mcs1_mcs_mat1_5_mcs_out[24]}), .b ({new_AGEMA_signal_9274, mcs1_mcs_mat1_5_mcs_out[28]}), .c ({new_AGEMA_signal_9525, mcs1_mcs_mat1_5_n117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U79 ( .a ({new_AGEMA_signal_9994, mcs1_mcs_mat1_5_mcs_out[16]}), .b ({new_AGEMA_signal_8446, mcs1_mcs_mat1_5_mcs_out[20]}), .c ({new_AGEMA_signal_10192, mcs1_mcs_mat1_5_n118}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U78 ( .a ({new_AGEMA_signal_9526, mcs1_mcs_mat1_5_n116}), .b ({new_AGEMA_signal_10193, mcs1_mcs_mat1_5_n115}), .c ({temp_next_s1[11], temp_next_s0[11]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U77 ( .a ({new_AGEMA_signal_9995, mcs1_mcs_mat1_5_mcs_out[3]}), .b ({new_AGEMA_signal_9280, mcs1_mcs_mat1_5_mcs_out[7]}), .c ({new_AGEMA_signal_10193, mcs1_mcs_mat1_5_n115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U76 ( .a ({new_AGEMA_signal_7531, mcs1_mcs_mat1_5_mcs_out[11]}), .b ({new_AGEMA_signal_9277, mcs1_mcs_mat1_5_mcs_out[15]}), .c ({new_AGEMA_signal_9526, mcs1_mcs_mat1_5_n116}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U75 ( .a ({new_AGEMA_signal_10433, mcs1_mcs_mat1_5_n114}), .b ({new_AGEMA_signal_9527, mcs1_mcs_mat1_5_n113}), .c ({new_AGEMA_signal_10698, mcs_out[235]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U74 ( .a ({new_AGEMA_signal_9251, mcs1_mcs_mat1_5_mcs_out[123]}), .b ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_9527, mcs1_mcs_mat1_5_n113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U73 ( .a ({new_AGEMA_signal_10205, mcs1_mcs_mat1_5_mcs_out[115]}), .b ({new_AGEMA_signal_9253, mcs1_mcs_mat1_5_mcs_out[119]}), .c ({new_AGEMA_signal_10433, mcs1_mcs_mat1_5_n114}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U72 ( .a ({new_AGEMA_signal_10194, mcs1_mcs_mat1_5_n112}), .b ({new_AGEMA_signal_8397, mcs1_mcs_mat1_5_n111}), .c ({new_AGEMA_signal_10434, mcs_out[234]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U71 ( .a ({new_AGEMA_signal_7918, mcs1_mcs_mat1_5_mcs_out[122]}), .b ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_8397, mcs1_mcs_mat1_5_n111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U70 ( .a ({new_AGEMA_signal_9980, mcs1_mcs_mat1_5_mcs_out[114]}), .b ({new_AGEMA_signal_9254, mcs1_mcs_mat1_5_mcs_out[118]}), .c ({new_AGEMA_signal_10194, mcs1_mcs_mat1_5_n112}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U69 ( .a ({new_AGEMA_signal_9241, mcs1_mcs_mat1_5_n110}), .b ({new_AGEMA_signal_10195, mcs1_mcs_mat1_5_n109}), .c ({temp_next_s1[10], temp_next_s0[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U68 ( .a ({new_AGEMA_signal_9996, mcs1_mcs_mat1_5_mcs_out[2]}), .b ({new_AGEMA_signal_8453, mcs1_mcs_mat1_5_mcs_out[6]}), .c ({new_AGEMA_signal_10195, mcs1_mcs_mat1_5_n109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U67 ( .a ({new_AGEMA_signal_8930, mcs1_mcs_mat1_5_mcs_out[10]}), .b ({new_AGEMA_signal_8927, mcs1_mcs_mat1_5_mcs_out[14]}), .c ({new_AGEMA_signal_9241, mcs1_mcs_mat1_5_n110}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U66 ( .a ({new_AGEMA_signal_9975, mcs1_mcs_mat1_5_n108}), .b ({new_AGEMA_signal_9528, mcs1_mcs_mat1_5_n107}), .c ({new_AGEMA_signal_10196, mcs_out[233]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U65 ( .a ({new_AGEMA_signal_9252, mcs1_mcs_mat1_5_mcs_out[121]}), .b ({new_AGEMA_signal_7497, mcs1_mcs_mat1_5_mcs_out[125]}), .c ({new_AGEMA_signal_9528, mcs1_mcs_mat1_5_n107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U64 ( .a ({new_AGEMA_signal_9758, mcs1_mcs_mat1_5_mcs_out[113]}), .b ({new_AGEMA_signal_8883, mcs1_mcs_mat1_5_mcs_out[117]}), .c ({new_AGEMA_signal_9975, mcs1_mcs_mat1_5_n108}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U63 ( .a ({new_AGEMA_signal_10699, mcs1_mcs_mat1_5_n106}), .b ({new_AGEMA_signal_9242, mcs1_mcs_mat1_5_n105}), .c ({new_AGEMA_signal_10915, mcs_out[232]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U62 ( .a ({new_AGEMA_signal_8880, mcs1_mcs_mat1_5_mcs_out[120]}), .b ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_9242, mcs1_mcs_mat1_5_n105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U61 ( .a ({new_AGEMA_signal_10447, mcs1_mcs_mat1_5_mcs_out[112]}), .b ({new_AGEMA_signal_8403, mcs1_mcs_mat1_5_mcs_out[116]}), .c ({new_AGEMA_signal_10699, mcs1_mcs_mat1_5_n106}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U60 ( .a ({new_AGEMA_signal_9243, mcs1_mcs_mat1_5_n104}), .b ({new_AGEMA_signal_10700, mcs1_mcs_mat1_5_n103}), .c ({new_AGEMA_signal_10916, mcs_out[203]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U59 ( .a ({new_AGEMA_signal_9255, mcs1_mcs_mat1_5_mcs_out[111]}), .b ({new_AGEMA_signal_10448, mcs1_mcs_mat1_5_mcs_out[99]}), .c ({new_AGEMA_signal_10700, mcs1_mcs_mat1_5_n103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U58 ( .a ({new_AGEMA_signal_8892, mcs1_mcs_mat1_5_mcs_out[103]}), .b ({new_AGEMA_signal_8888, mcs1_mcs_mat1_5_mcs_out[107]}), .c ({new_AGEMA_signal_9243, mcs1_mcs_mat1_5_n104}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U57 ( .a ({new_AGEMA_signal_9244, mcs1_mcs_mat1_5_n102}), .b ({new_AGEMA_signal_10197, mcs1_mcs_mat1_5_n101}), .c ({new_AGEMA_signal_10436, mcs_out[202]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U56 ( .a ({new_AGEMA_signal_9256, mcs1_mcs_mat1_5_mcs_out[110]}), .b ({new_AGEMA_signal_9983, mcs1_mcs_mat1_5_mcs_out[98]}), .c ({new_AGEMA_signal_10197, mcs1_mcs_mat1_5_n101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U55 ( .a ({new_AGEMA_signal_7927, mcs1_mcs_mat1_5_mcs_out[102]}), .b ({new_AGEMA_signal_8889, mcs1_mcs_mat1_5_mcs_out[106]}), .c ({new_AGEMA_signal_9244, mcs1_mcs_mat1_5_n102}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U54 ( .a ({new_AGEMA_signal_9245, mcs1_mcs_mat1_5_n100}), .b ({new_AGEMA_signal_9755, mcs1_mcs_mat1_5_n99}), .c ({new_AGEMA_signal_9976, mcs_out[201]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U53 ( .a ({new_AGEMA_signal_9257, mcs1_mcs_mat1_5_mcs_out[109]}), .b ({new_AGEMA_signal_9538, mcs1_mcs_mat1_5_mcs_out[97]}), .c ({new_AGEMA_signal_9755, mcs1_mcs_mat1_5_n99}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U52 ( .a ({new_AGEMA_signal_8410, mcs1_mcs_mat1_5_mcs_out[101]}), .b ({new_AGEMA_signal_8890, mcs1_mcs_mat1_5_mcs_out[105]}), .c ({new_AGEMA_signal_9245, mcs1_mcs_mat1_5_n100}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U51 ( .a ({new_AGEMA_signal_9529, mcs1_mcs_mat1_5_n98}), .b ({new_AGEMA_signal_11053, mcs1_mcs_mat1_5_n97}), .c ({new_AGEMA_signal_11100, mcs_out[200]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U50 ( .a ({new_AGEMA_signal_9258, mcs1_mcs_mat1_5_mcs_out[108]}), .b ({new_AGEMA_signal_10919, mcs1_mcs_mat1_5_mcs_out[96]}), .c ({new_AGEMA_signal_11053, mcs1_mcs_mat1_5_n97}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U49 ( .a ({new_AGEMA_signal_8893, mcs1_mcs_mat1_5_mcs_out[100]}), .b ({new_AGEMA_signal_9259, mcs1_mcs_mat1_5_mcs_out[104]}), .c ({new_AGEMA_signal_9529, mcs1_mcs_mat1_5_n98}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U48 ( .a ({new_AGEMA_signal_10198, mcs1_mcs_mat1_5_n96}), .b ({new_AGEMA_signal_9246, mcs1_mcs_mat1_5_n95}), .c ({new_AGEMA_signal_10437, mcs_out[171]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U47 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_8896, mcs1_mcs_mat1_5_mcs_out[95]}), .c ({new_AGEMA_signal_9246, mcs1_mcs_mat1_5_n95}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U46 ( .a ({new_AGEMA_signal_9984, mcs1_mcs_mat1_5_mcs_out[83]}), .b ({new_AGEMA_signal_7934, mcs1_mcs_mat1_5_mcs_out[87]}), .c ({new_AGEMA_signal_10198, mcs1_mcs_mat1_5_n96}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U45 ( .a ({new_AGEMA_signal_10199, mcs1_mcs_mat1_5_n94}), .b ({new_AGEMA_signal_8398, mcs1_mcs_mat1_5_n93}), .c ({new_AGEMA_signal_10438, mcs_out[170]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U43 ( .a ({new_AGEMA_signal_9985, mcs1_mcs_mat1_5_mcs_out[82]}), .b ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_10199, mcs1_mcs_mat1_5_n94}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U42 ( .a ({new_AGEMA_signal_10200, mcs1_mcs_mat1_5_n92}), .b ({new_AGEMA_signal_8399, mcs1_mcs_mat1_5_n91}), .c ({new_AGEMA_signal_10439, mcs_out[169]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U41 ( .a ({new_AGEMA_signal_7512, mcs1_mcs_mat1_5_mcs_out[89]}), .b ({new_AGEMA_signal_7932, mcs1_mcs_mat1_5_mcs_out[93]}), .c ({new_AGEMA_signal_8399, mcs1_mcs_mat1_5_n91}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U40 ( .a ({new_AGEMA_signal_9986, mcs1_mcs_mat1_5_mcs_out[81]}), .b ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_10200, mcs1_mcs_mat1_5_n92}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U39 ( .a ({new_AGEMA_signal_10440, mcs1_mcs_mat1_5_n90}), .b ({new_AGEMA_signal_9530, mcs1_mcs_mat1_5_n89}), .c ({new_AGEMA_signal_10701, mcs_out[168]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U38 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_9260, mcs1_mcs_mat1_5_mcs_out[92]}), .c ({new_AGEMA_signal_9530, mcs1_mcs_mat1_5_n89}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U37 ( .a ({new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[80]}), .b ({new_AGEMA_signal_8414, mcs1_mcs_mat1_5_mcs_out[84]}), .c ({new_AGEMA_signal_10440, mcs1_mcs_mat1_5_n90}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U36 ( .a ({new_AGEMA_signal_10441, mcs1_mcs_mat1_5_n88}), .b ({new_AGEMA_signal_8874, mcs1_mcs_mat1_5_n87}), .c ({temp_next_s1[9], temp_next_s0[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U35 ( .a ({new_AGEMA_signal_7533, mcs1_mcs_mat1_5_mcs_out[5]}), .b ({new_AGEMA_signal_8451, mcs1_mcs_mat1_5_mcs_out[9]}), .c ({new_AGEMA_signal_8874, mcs1_mcs_mat1_5_n87}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U34 ( .a ({new_AGEMA_signal_8928, mcs1_mcs_mat1_5_mcs_out[13]}), .b ({new_AGEMA_signal_10214, mcs1_mcs_mat1_5_mcs_out[1]}), .c ({new_AGEMA_signal_10441, mcs1_mcs_mat1_5_n88}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U33 ( .a ({new_AGEMA_signal_10703, mcs1_mcs_mat1_5_n86}), .b ({new_AGEMA_signal_9247, mcs1_mcs_mat1_5_n85}), .c ({new_AGEMA_signal_10917, mcs_out[139]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U32 ( .a ({new_AGEMA_signal_7937, mcs1_mcs_mat1_5_mcs_out[75]}), .b ({new_AGEMA_signal_8899, mcs1_mcs_mat1_5_mcs_out[79]}), .c ({new_AGEMA_signal_9247, mcs1_mcs_mat1_5_n85}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U31 ( .a ({new_AGEMA_signal_10449, mcs1_mcs_mat1_5_mcs_out[67]}), .b ({new_AGEMA_signal_8903, mcs1_mcs_mat1_5_mcs_out[71]}), .c ({new_AGEMA_signal_10703, mcs1_mcs_mat1_5_n86}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U30 ( .a ({new_AGEMA_signal_10442, mcs1_mcs_mat1_5_n84}), .b ({new_AGEMA_signal_9531, mcs1_mcs_mat1_5_n83}), .c ({new_AGEMA_signal_10704, mcs_out[138]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U29 ( .a ({new_AGEMA_signal_9262, mcs1_mcs_mat1_5_mcs_out[74]}), .b ({new_AGEMA_signal_7098, mcs1_mcs_mat1_5_mcs_out[78]}), .c ({new_AGEMA_signal_9531, mcs1_mcs_mat1_5_n83}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U28 ( .a ({new_AGEMA_signal_10209, mcs1_mcs_mat1_5_mcs_out[66]}), .b ({new_AGEMA_signal_9264, mcs1_mcs_mat1_5_mcs_out[70]}), .c ({new_AGEMA_signal_10442, mcs1_mcs_mat1_5_n84}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U27 ( .a ({new_AGEMA_signal_9977, mcs1_mcs_mat1_5_n82}), .b ({new_AGEMA_signal_8875, mcs1_mcs_mat1_5_n81}), .c ({new_AGEMA_signal_10201, mcs_out[137]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U26 ( .a ({new_AGEMA_signal_8417, mcs1_mcs_mat1_5_mcs_out[73]}), .b ({new_AGEMA_signal_7935, mcs1_mcs_mat1_5_mcs_out[77]}), .c ({new_AGEMA_signal_8875, mcs1_mcs_mat1_5_n81}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U25 ( .a ({new_AGEMA_signal_9766, mcs1_mcs_mat1_5_mcs_out[65]}), .b ({new_AGEMA_signal_9265, mcs1_mcs_mat1_5_mcs_out[69]}), .c ({new_AGEMA_signal_9977, mcs1_mcs_mat1_5_n82}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U24 ( .a ({new_AGEMA_signal_10918, mcs1_mcs_mat1_5_n80}), .b ({new_AGEMA_signal_9532, mcs1_mcs_mat1_5_n79}), .c ({new_AGEMA_signal_11054, mcs_out[136]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U23 ( .a ({new_AGEMA_signal_9263, mcs1_mcs_mat1_5_mcs_out[72]}), .b ({new_AGEMA_signal_9261, mcs1_mcs_mat1_5_mcs_out[76]}), .c ({new_AGEMA_signal_9532, mcs1_mcs_mat1_5_n79}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U22 ( .a ({new_AGEMA_signal_10708, mcs1_mcs_mat1_5_mcs_out[64]}), .b ({new_AGEMA_signal_8905, mcs1_mcs_mat1_5_mcs_out[68]}), .c ({new_AGEMA_signal_10918, mcs1_mcs_mat1_5_n80}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U21 ( .a ({new_AGEMA_signal_9978, mcs1_mcs_mat1_5_n78}), .b ({new_AGEMA_signal_9248, mcs1_mcs_mat1_5_n77}), .c ({temp_next_s1[107], temp_next_s0[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U20 ( .a ({new_AGEMA_signal_8425, mcs1_mcs_mat1_5_mcs_out[59]}), .b ({new_AGEMA_signal_8907, mcs1_mcs_mat1_5_mcs_out[63]}), .c ({new_AGEMA_signal_9248, mcs1_mcs_mat1_5_n77}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U19 ( .a ({new_AGEMA_signal_9768, mcs1_mcs_mat1_5_mcs_out[51]}), .b ({new_AGEMA_signal_8910, mcs1_mcs_mat1_5_mcs_out[55]}), .c ({new_AGEMA_signal_9978, mcs1_mcs_mat1_5_n78}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U18 ( .a ({new_AGEMA_signal_9533, mcs1_mcs_mat1_5_n76}), .b ({new_AGEMA_signal_8876, mcs1_mcs_mat1_5_n75}), .c ({temp_next_s1[106], temp_next_s0[106]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U17 ( .a ({new_AGEMA_signal_7945, mcs1_mcs_mat1_5_mcs_out[58]}), .b ({new_AGEMA_signal_8422, mcs1_mcs_mat1_5_mcs_out[62]}), .c ({new_AGEMA_signal_8876, mcs1_mcs_mat1_5_n75}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U16 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_9267, mcs1_mcs_mat1_5_mcs_out[54]}), .c ({new_AGEMA_signal_9533, mcs1_mcs_mat1_5_n76}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U15 ( .a ({new_AGEMA_signal_9534, mcs1_mcs_mat1_5_n74}), .b ({new_AGEMA_signal_8877, mcs1_mcs_mat1_5_n73}), .c ({temp_next_s1[105], temp_next_s0[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U14 ( .a ({new_AGEMA_signal_8426, mcs1_mcs_mat1_5_mcs_out[57]}), .b ({new_AGEMA_signal_8423, mcs1_mcs_mat1_5_mcs_out[61]}), .c ({new_AGEMA_signal_8877, mcs1_mcs_mat1_5_n73}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U13 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_9268, mcs1_mcs_mat1_5_mcs_out[53]}), .c ({new_AGEMA_signal_9534, mcs1_mcs_mat1_5_n74}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U12 ( .a ({new_AGEMA_signal_10203, mcs1_mcs_mat1_5_n72}), .b ({new_AGEMA_signal_9535, mcs1_mcs_mat1_5_n71}), .c ({temp_next_s1[104], temp_next_s0[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U11 ( .a ({new_AGEMA_signal_8909, mcs1_mcs_mat1_5_mcs_out[56]}), .b ({new_AGEMA_signal_9266, mcs1_mcs_mat1_5_mcs_out[60]}), .c ({new_AGEMA_signal_9535, mcs1_mcs_mat1_5_n71}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U10 ( .a ({new_AGEMA_signal_9989, mcs1_mcs_mat1_5_mcs_out[48]}), .b ({new_AGEMA_signal_8912, mcs1_mcs_mat1_5_mcs_out[52]}), .c ({new_AGEMA_signal_10203, mcs1_mcs_mat1_5_n72}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U9 ( .a ({new_AGEMA_signal_10444, mcs1_mcs_mat1_5_n70}), .b ({new_AGEMA_signal_9249, mcs1_mcs_mat1_5_n69}), .c ({temp_next_s1[75], temp_next_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U8 ( .a ({new_AGEMA_signal_8914, mcs1_mcs_mat1_5_mcs_out[43]}), .b ({new_AGEMA_signal_8913, mcs1_mcs_mat1_5_mcs_out[47]}), .c ({new_AGEMA_signal_9249, mcs1_mcs_mat1_5_n69}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U7 ( .a ({new_AGEMA_signal_10211, mcs1_mcs_mat1_5_mcs_out[35]}), .b ({new_AGEMA_signal_9270, mcs1_mcs_mat1_5_mcs_out[39]}), .c ({new_AGEMA_signal_10444, mcs1_mcs_mat1_5_n70}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U6 ( .a ({new_AGEMA_signal_10204, mcs1_mcs_mat1_5_n68}), .b ({new_AGEMA_signal_9250, mcs1_mcs_mat1_5_n67}), .c ({temp_next_s1[74], temp_next_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U5 ( .a ({new_AGEMA_signal_8915, mcs1_mcs_mat1_5_mcs_out[42]}), .b ({new_AGEMA_signal_7520, mcs1_mcs_mat1_5_mcs_out[46]}), .c ({new_AGEMA_signal_9250, mcs1_mcs_mat1_5_n67}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U4 ( .a ({new_AGEMA_signal_9990, mcs1_mcs_mat1_5_mcs_out[34]}), .b ({new_AGEMA_signal_7958, mcs1_mcs_mat1_5_mcs_out[38]}), .c ({new_AGEMA_signal_10204, mcs1_mcs_mat1_5_n68}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U3 ( .a ({new_AGEMA_signal_10446, mcs1_mcs_mat1_5_n66}), .b ({new_AGEMA_signal_9979, mcs1_mcs_mat1_5_n65}), .c ({temp_next_s1[8], temp_next_s0[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U2 ( .a ({new_AGEMA_signal_9775, mcs1_mcs_mat1_5_mcs_out[4]}), .b ({new_AGEMA_signal_9279, mcs1_mcs_mat1_5_mcs_out[8]}), .c ({new_AGEMA_signal_9979, mcs1_mcs_mat1_5_n65}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_U1 ( .a ({new_AGEMA_signal_10215, mcs1_mcs_mat1_5_mcs_out[0]}), .b ({new_AGEMA_signal_9546, mcs1_mcs_mat1_5_mcs_out[12]}), .c ({new_AGEMA_signal_10446, mcs1_mcs_mat1_5_n66}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_8878, mcs1_mcs_mat1_5_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_9251, mcs1_mcs_mat1_5_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_8400, mcs1_mcs_mat1_5_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_6805, mcs1_mcs_mat1_5_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8878, mcs1_mcs_mat1_5_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_7091, mcs1_mcs_mat1_5_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_7498, mcs1_mcs_mat1_5_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_7918, mcs1_mcs_mat1_5_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_7092, mcs1_mcs_mat1_5_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_7229, shiftr_out[75]}), .c ({new_AGEMA_signal_7498, mcs1_mcs_mat1_5_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_8879, mcs1_mcs_mat1_5_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_7229, shiftr_out[75]}), .c ({new_AGEMA_signal_9252, mcs1_mcs_mat1_5_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_8400, mcs1_mcs_mat1_5_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_8879, mcs1_mcs_mat1_5_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_7919, mcs1_mcs_mat1_5_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_7499, mcs1_mcs_mat1_5_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_8400, mcs1_mcs_mat1_5_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_8401, mcs1_mcs_mat1_5_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_8880, mcs1_mcs_mat1_5_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_7919, mcs1_mcs_mat1_5_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_7092, mcs1_mcs_mat1_5_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_8401, mcs1_mcs_mat1_5_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[868]), .c ({new_AGEMA_signal_7919, mcs1_mcs_mat1_5_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[869]), .c ({new_AGEMA_signal_7092, mcs1_mcs_mat1_5_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7229, shiftr_out[75]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[870]), .c ({new_AGEMA_signal_7499, mcs1_mcs_mat1_5_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_8881, mcs1_mcs_mat1_5_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_6689, shiftr_out[42]}), .c ({new_AGEMA_signal_9253, mcs1_mcs_mat1_5_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_8402, mcs1_mcs_mat1_5_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7502, mcs1_mcs_mat1_5_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_8881, mcs1_mcs_mat1_5_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_8882, mcs1_mcs_mat1_5_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_7921, mcs1_mcs_mat1_5_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_9254, mcs1_mcs_mat1_5_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_8402, mcs1_mcs_mat1_5_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7301, shiftr_out[41]}), .c ({new_AGEMA_signal_8882, mcs1_mcs_mat1_5_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_8402, mcs1_mcs_mat1_5_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7920, mcs1_mcs_mat1_5_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_8883, mcs1_mcs_mat1_5_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_7922, mcs1_mcs_mat1_5_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_7093, mcs1_mcs_mat1_5_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_8402, mcs1_mcs_mat1_5_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_7501, mcs1_mcs_mat1_5_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_7921, mcs1_mcs_mat1_5_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_8403, mcs1_mcs_mat1_5_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_6806, mcs1_mcs_mat1_5_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7502, mcs1_mcs_mat1_5_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_7921, mcs1_mcs_mat1_5_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_7093, mcs1_mcs_mat1_5_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_7501, mcs1_mcs_mat1_5_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7301, shiftr_out[41]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[871]), .c ({new_AGEMA_signal_7922, mcs1_mcs_mat1_5_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[872]), .c ({new_AGEMA_signal_7093, mcs1_mcs_mat1_5_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[873]), .c ({new_AGEMA_signal_7502, mcs1_mcs_mat1_5_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_9981, mcs1_mcs_mat1_5_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_8884, mcs1_mcs_mat1_5_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_10205, mcs1_mcs_mat1_5_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_9536, mcs1_mcs_mat1_5_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_9537, mcs1_mcs_mat1_5_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_9758, mcs1_mcs_mat1_5_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_9982, mcs1_mcs_mat1_5_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_10206, mcs1_mcs_mat1_5_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_10447, mcs1_mcs_mat1_5_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_9981, mcs1_mcs_mat1_5_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_10206, mcs1_mcs_mat1_5_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_8404, mcs1_mcs_mat1_5_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9760, mcs1_mcs_mat1_5_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_9981, mcs1_mcs_mat1_5_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_8885, mcs1_mcs_mat1_5_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_9759, mcs1_mcs_mat1_5_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_9982, mcs1_mcs_mat1_5_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9362, shiftr_out[9]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[874]), .c ({new_AGEMA_signal_9760, mcs1_mcs_mat1_5_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[875]), .c ({new_AGEMA_signal_8885, mcs1_mcs_mat1_5_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[876]), .c ({new_AGEMA_signal_9537, mcs1_mcs_mat1_5_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({new_AGEMA_signal_8886, mcs1_mcs_mat1_5_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9255, mcs1_mcs_mat1_5_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({new_AGEMA_signal_8887, mcs1_mcs_mat1_5_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9256, mcs1_mcs_mat1_5_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_7503, mcs1_mcs_mat1_5_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_8886, mcs1_mcs_mat1_5_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9257, mcs1_mcs_mat1_5_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_7094, mcs1_mcs_mat1_5_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_8405, mcs1_mcs_mat1_5_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_8886, mcs1_mcs_mat1_5_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_7923, mcs1_mcs_mat1_5_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8887, mcs1_mcs_mat1_5_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9258, mcs1_mcs_mat1_5_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_8406, mcs1_mcs_mat1_5_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_8887, mcs1_mcs_mat1_5_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_7503, mcs1_mcs_mat1_5_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_7924, mcs1_mcs_mat1_5_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_8406, mcs1_mcs_mat1_5_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[877]), .c ({new_AGEMA_signal_7924, mcs1_mcs_mat1_5_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[878]), .c ({new_AGEMA_signal_7094, mcs1_mcs_mat1_5_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[879]), .c ({new_AGEMA_signal_7503, mcs1_mcs_mat1_5_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_8408, mcs1_mcs_mat1_5_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_8407, mcs1_mcs_mat1_5_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8888, mcs1_mcs_mat1_5_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_8407, mcs1_mcs_mat1_5_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_7504, mcs1_mcs_mat1_5_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_8889, mcs1_mcs_mat1_5_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_7095, mcs1_mcs_mat1_5_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7229, shiftr_out[75]}), .c ({new_AGEMA_signal_7504, mcs1_mcs_mat1_5_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_8407, mcs1_mcs_mat1_5_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8890, mcs1_mcs_mat1_5_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_7926, mcs1_mcs_mat1_5_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_6808, mcs1_mcs_mat1_5_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_8407, mcs1_mcs_mat1_5_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_8891, mcs1_mcs_mat1_5_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_9259, mcs1_mcs_mat1_5_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_8408, mcs1_mcs_mat1_5_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_7926, mcs1_mcs_mat1_5_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_8891, mcs1_mcs_mat1_5_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_7925, mcs1_mcs_mat1_5_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_6615, shiftr_out[72]}), .c ({new_AGEMA_signal_8408, mcs1_mcs_mat1_5_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_7095, mcs1_mcs_mat1_5_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7505, mcs1_mcs_mat1_5_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_7925, mcs1_mcs_mat1_5_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[880]), .c ({new_AGEMA_signal_7926, mcs1_mcs_mat1_5_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[881]), .c ({new_AGEMA_signal_7095, mcs1_mcs_mat1_5_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7229, shiftr_out[75]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[882]), .c ({new_AGEMA_signal_7505, mcs1_mcs_mat1_5_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_7506, mcs1_mcs_mat1_5_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_8409, mcs1_mcs_mat1_5_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_8892, mcs1_mcs_mat1_5_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_7930, mcs1_mcs_mat1_5_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_8409, mcs1_mcs_mat1_5_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_7928, mcs1_mcs_mat1_5_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_7507, mcs1_mcs_mat1_5_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_8410, mcs1_mcs_mat1_5_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_7929, mcs1_mcs_mat1_5_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_8411, mcs1_mcs_mat1_5_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_8893, mcs1_mcs_mat1_5_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_6809, mcs1_mcs_mat1_5_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_7930, mcs1_mcs_mat1_5_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_8411, mcs1_mcs_mat1_5_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_7096, mcs1_mcs_mat1_5_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_7301, shiftr_out[41]}), .c ({new_AGEMA_signal_7929, mcs1_mcs_mat1_5_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7301, shiftr_out[41]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[883]), .c ({new_AGEMA_signal_7930, mcs1_mcs_mat1_5_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[884]), .c ({new_AGEMA_signal_7096, mcs1_mcs_mat1_5_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[885]), .c ({new_AGEMA_signal_7507, mcs1_mcs_mat1_5_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_10707, mcs1_mcs_mat1_5_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_9539, mcs1_mcs_mat1_5_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_10919, mcs1_mcs_mat1_5_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_10448, mcs1_mcs_mat1_5_mcs_out[99]}), .b ({new_AGEMA_signal_8100, shiftr_out[10]}), .c ({new_AGEMA_signal_10707, mcs1_mcs_mat1_5_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_10207, mcs1_mcs_mat1_5_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_9362, shiftr_out[9]}), .c ({new_AGEMA_signal_10448, mcs1_mcs_mat1_5_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_9983, mcs1_mcs_mat1_5_mcs_out[98]}), .b ({new_AGEMA_signal_8895, mcs1_mcs_mat1_5_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_10207, mcs1_mcs_mat1_5_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_8894, mcs1_mcs_mat1_5_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_9761, mcs1_mcs_mat1_5_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_9983, mcs1_mcs_mat1_5_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9362, shiftr_out[9]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[886]), .c ({new_AGEMA_signal_9761, mcs1_mcs_mat1_5_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[887]), .c ({new_AGEMA_signal_8895, mcs1_mcs_mat1_5_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[888]), .c ({new_AGEMA_signal_9539, mcs1_mcs_mat1_5_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_8413, mcs1_mcs_mat1_5_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_8896, mcs1_mcs_mat1_5_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_7509, mcs1_mcs_mat1_5_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_7932, mcs1_mcs_mat1_5_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_8897, mcs1_mcs_mat1_5_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_7097, mcs1_mcs_mat1_5_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_9260, mcs1_mcs_mat1_5_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_8413, mcs1_mcs_mat1_5_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_8897, mcs1_mcs_mat1_5_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_6810, mcs1_mcs_mat1_5_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7933, mcs1_mcs_mat1_5_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_8413, mcs1_mcs_mat1_5_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[889]), .c ({new_AGEMA_signal_7933, mcs1_mcs_mat1_5_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[890]), .c ({new_AGEMA_signal_7097, mcs1_mcs_mat1_5_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[891]), .c ({new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_9764, mcs1_mcs_mat1_5_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_9765, mcs1_mcs_mat1_5_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_9984, mcs1_mcs_mat1_5_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_9762, mcs1_mcs_mat1_5_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_8415, mcs1_mcs_mat1_5_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_9985, mcs1_mcs_mat1_5_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_9540, mcs1_mcs_mat1_5_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_9762, mcs1_mcs_mat1_5_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_9763, mcs1_mcs_mat1_5_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_9986, mcs1_mcs_mat1_5_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_8898, mcs1_mcs_mat1_5_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_9540, mcs1_mcs_mat1_5_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_9763, mcs1_mcs_mat1_5_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_9987, mcs1_mcs_mat1_5_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_8100, shiftr_out[10]}), .c ({new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_9764, mcs1_mcs_mat1_5_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_8898, mcs1_mcs_mat1_5_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_9987, mcs1_mcs_mat1_5_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9362, shiftr_out[9]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[892]), .c ({new_AGEMA_signal_9765, mcs1_mcs_mat1_5_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[893]), .c ({new_AGEMA_signal_8898, mcs1_mcs_mat1_5_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[894]), .c ({new_AGEMA_signal_9540, mcs1_mcs_mat1_5_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_8416, mcs1_mcs_mat1_5_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_8899, mcs1_mcs_mat1_5_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_7513, mcs1_mcs_mat1_5_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_7935, mcs1_mcs_mat1_5_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_8900, mcs1_mcs_mat1_5_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_7099, mcs1_mcs_mat1_5_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_9261, mcs1_mcs_mat1_5_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_8416, mcs1_mcs_mat1_5_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_6610, shiftr_out[104]}), .c ({new_AGEMA_signal_8900, mcs1_mcs_mat1_5_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_6811, mcs1_mcs_mat1_5_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7936, mcs1_mcs_mat1_5_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_8416, mcs1_mcs_mat1_5_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[895]), .c ({new_AGEMA_signal_7936, mcs1_mcs_mat1_5_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[896]), .c ({new_AGEMA_signal_7099, mcs1_mcs_mat1_5_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[897]), .c ({new_AGEMA_signal_7513, mcs1_mcs_mat1_5_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_8901, mcs1_mcs_mat1_5_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_9262, mcs1_mcs_mat1_5_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_8418, mcs1_mcs_mat1_5_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7938, mcs1_mcs_mat1_5_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_8901, mcs1_mcs_mat1_5_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_7265, mcs1_mcs_mat1_5_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_7937, mcs1_mcs_mat1_5_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_7938, mcs1_mcs_mat1_5_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_7265, mcs1_mcs_mat1_5_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_8417, mcs1_mcs_mat1_5_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_7100, mcs1_mcs_mat1_5_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_7101, mcs1_mcs_mat1_5_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_7265, mcs1_mcs_mat1_5_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_7514, mcs1_mcs_mat1_5_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_6615, shiftr_out[72]}), .c ({new_AGEMA_signal_7938, mcs1_mcs_mat1_5_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_8902, mcs1_mcs_mat1_5_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_7100, mcs1_mcs_mat1_5_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_9263, mcs1_mcs_mat1_5_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_8418, mcs1_mcs_mat1_5_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7514, mcs1_mcs_mat1_5_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_8902, mcs1_mcs_mat1_5_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_7229, shiftr_out[75]}), .b ({new_AGEMA_signal_7939, mcs1_mcs_mat1_5_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_8418, mcs1_mcs_mat1_5_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[898]), .c ({new_AGEMA_signal_7939, mcs1_mcs_mat1_5_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[899]), .c ({new_AGEMA_signal_7101, mcs1_mcs_mat1_5_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7229, shiftr_out[75]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[900]), .c ({new_AGEMA_signal_7514, mcs1_mcs_mat1_5_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_8419, mcs1_mcs_mat1_5_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_7515, mcs1_mcs_mat1_5_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_8903, mcs1_mcs_mat1_5_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_7941, mcs1_mcs_mat1_5_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_8904, mcs1_mcs_mat1_5_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9264, mcs1_mcs_mat1_5_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_8419, mcs1_mcs_mat1_5_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_8904, mcs1_mcs_mat1_5_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9265, mcs1_mcs_mat1_5_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_7515, mcs1_mcs_mat1_5_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_8420, mcs1_mcs_mat1_5_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_8904, mcs1_mcs_mat1_5_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({new_AGEMA_signal_7102, mcs1_mcs_mat1_5_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_7515, mcs1_mcs_mat1_5_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_7940, mcs1_mcs_mat1_5_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_7301, shiftr_out[41]}), .c ({new_AGEMA_signal_8419, mcs1_mcs_mat1_5_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_7516, mcs1_mcs_mat1_5_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6813, mcs1_mcs_mat1_5_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_7940, mcs1_mcs_mat1_5_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_8420, mcs1_mcs_mat1_5_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_7941, mcs1_mcs_mat1_5_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_8905, mcs1_mcs_mat1_5_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_7516, mcs1_mcs_mat1_5_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_7941, mcs1_mcs_mat1_5_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({new_AGEMA_signal_7942, mcs1_mcs_mat1_5_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_8420, mcs1_mcs_mat1_5_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7301, shiftr_out[41]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[901]), .c ({new_AGEMA_signal_7942, mcs1_mcs_mat1_5_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[902]), .c ({new_AGEMA_signal_7102, mcs1_mcs_mat1_5_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[903]), .c ({new_AGEMA_signal_7516, mcs1_mcs_mat1_5_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_10210, mcs1_mcs_mat1_5_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_10449, mcs1_mcs_mat1_5_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({new_AGEMA_signal_9988, mcs1_mcs_mat1_5_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_10209, mcs1_mcs_mat1_5_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_10450, mcs1_mcs_mat1_5_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_9541, mcs1_mcs_mat1_5_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_10708, mcs1_mcs_mat1_5_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_10210, mcs1_mcs_mat1_5_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .c ({new_AGEMA_signal_10450, mcs1_mcs_mat1_5_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_8906, mcs1_mcs_mat1_5_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_9988, mcs1_mcs_mat1_5_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_10210, mcs1_mcs_mat1_5_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_8421, mcs1_mcs_mat1_5_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_9767, mcs1_mcs_mat1_5_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_9988, mcs1_mcs_mat1_5_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9362, shiftr_out[9]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[904]), .c ({new_AGEMA_signal_9767, mcs1_mcs_mat1_5_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[905]), .c ({new_AGEMA_signal_8906, mcs1_mcs_mat1_5_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[906]), .c ({new_AGEMA_signal_9541, mcs1_mcs_mat1_5_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_8424, mcs1_mcs_mat1_5_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7517, mcs1_mcs_mat1_5_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_8907, mcs1_mcs_mat1_5_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_7103, mcs1_mcs_mat1_5_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_7943, mcs1_mcs_mat1_5_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8422, mcs1_mcs_mat1_5_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({new_AGEMA_signal_7944, mcs1_mcs_mat1_5_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_8423, mcs1_mcs_mat1_5_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[907]), .c ({new_AGEMA_signal_7944, mcs1_mcs_mat1_5_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[908]), .c ({new_AGEMA_signal_7103, mcs1_mcs_mat1_5_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[909]), .c ({new_AGEMA_signal_7517, mcs1_mcs_mat1_5_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_7105, mcs1_mcs_mat1_5_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_7518, mcs1_mcs_mat1_5_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_7945, mcs1_mcs_mat1_5_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_7106, mcs1_mcs_mat1_5_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_7946, mcs1_mcs_mat1_5_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_8426, mcs1_mcs_mat1_5_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_8427, mcs1_mcs_mat1_5_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_7947, mcs1_mcs_mat1_5_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_8909, mcs1_mcs_mat1_5_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_7948, mcs1_mcs_mat1_5_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_8427, mcs1_mcs_mat1_5_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[910]), .c ({new_AGEMA_signal_7948, mcs1_mcs_mat1_5_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[911]), .c ({new_AGEMA_signal_7106, mcs1_mcs_mat1_5_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7229, shiftr_out[75]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[912]), .c ({new_AGEMA_signal_7518, mcs1_mcs_mat1_5_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_7950, mcs1_mcs_mat1_5_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8428, mcs1_mcs_mat1_5_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_8910, mcs1_mcs_mat1_5_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_8911, mcs1_mcs_mat1_5_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_7949, mcs1_mcs_mat1_5_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_9267, mcs1_mcs_mat1_5_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_7519, mcs1_mcs_mat1_5_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_7949, mcs1_mcs_mat1_5_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({new_AGEMA_signal_8911, mcs1_mcs_mat1_5_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_9268, mcs1_mcs_mat1_5_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_6816, mcs1_mcs_mat1_5_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_8428, mcs1_mcs_mat1_5_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_8911, mcs1_mcs_mat1_5_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_7107, mcs1_mcs_mat1_5_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_7952, mcs1_mcs_mat1_5_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_8428, mcs1_mcs_mat1_5_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_7951, mcs1_mcs_mat1_5_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_8429, mcs1_mcs_mat1_5_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_8912, mcs1_mcs_mat1_5_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_7950, mcs1_mcs_mat1_5_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_7107, mcs1_mcs_mat1_5_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_8429, mcs1_mcs_mat1_5_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_7519, mcs1_mcs_mat1_5_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_7950, mcs1_mcs_mat1_5_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7301, shiftr_out[41]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[913]), .c ({new_AGEMA_signal_7952, mcs1_mcs_mat1_5_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[914]), .c ({new_AGEMA_signal_7107, mcs1_mcs_mat1_5_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[915]), .c ({new_AGEMA_signal_7519, mcs1_mcs_mat1_5_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_7521, mcs1_mcs_mat1_5_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_7953, mcs1_mcs_mat1_5_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_9269, mcs1_mcs_mat1_5_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_7108, mcs1_mcs_mat1_5_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_9542, mcs1_mcs_mat1_5_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_8913, mcs1_mcs_mat1_5_mcs_out[47]}), .b ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_9269, mcs1_mcs_mat1_5_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_8430, mcs1_mcs_mat1_5_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_6610, shiftr_out[104]}), .c ({new_AGEMA_signal_8913, mcs1_mcs_mat1_5_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_6817, mcs1_mcs_mat1_5_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_7954, mcs1_mcs_mat1_5_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_8430, mcs1_mcs_mat1_5_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[916]), .c ({new_AGEMA_signal_7954, mcs1_mcs_mat1_5_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[917]), .c ({new_AGEMA_signal_7108, mcs1_mcs_mat1_5_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[918]), .c ({new_AGEMA_signal_7521, mcs1_mcs_mat1_5_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_8431, mcs1_mcs_mat1_5_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_7522, mcs1_mcs_mat1_5_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_8914, mcs1_mcs_mat1_5_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_7955, mcs1_mcs_mat1_5_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7109, mcs1_mcs_mat1_5_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_8431, mcs1_mcs_mat1_5_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_8432, mcs1_mcs_mat1_5_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_7957, mcs1_mcs_mat1_5_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_8915, mcs1_mcs_mat1_5_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_8433, mcs1_mcs_mat1_5_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_6818, mcs1_mcs_mat1_5_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_8916, mcs1_mcs_mat1_5_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_7955, mcs1_mcs_mat1_5_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7523, mcs1_mcs_mat1_5_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8433, mcs1_mcs_mat1_5_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_7956, mcs1_mcs_mat1_5_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_7523, mcs1_mcs_mat1_5_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8434, mcs1_mcs_mat1_5_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[919]), .c ({new_AGEMA_signal_7957, mcs1_mcs_mat1_5_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[920]), .c ({new_AGEMA_signal_7109, mcs1_mcs_mat1_5_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7229, shiftr_out[75]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[921]), .c ({new_AGEMA_signal_7523, mcs1_mcs_mat1_5_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_8917, mcs1_mcs_mat1_5_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_6819, mcs1_mcs_mat1_5_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9270, mcs1_mcs_mat1_5_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_7525, mcs1_mcs_mat1_5_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_7524, mcs1_mcs_mat1_5_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_7958, mcs1_mcs_mat1_5_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({new_AGEMA_signal_8917, mcs1_mcs_mat1_5_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_9271, mcs1_mcs_mat1_5_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_7959, mcs1_mcs_mat1_5_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_8435, mcs1_mcs_mat1_5_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_8917, mcs1_mcs_mat1_5_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_7960, mcs1_mcs_mat1_5_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7526, mcs1_mcs_mat1_5_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_8435, mcs1_mcs_mat1_5_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_7960, mcs1_mcs_mat1_5_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7525, mcs1_mcs_mat1_5_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_8436, mcs1_mcs_mat1_5_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_7266, mcs1_mcs_mat1_5_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_7525, mcs1_mcs_mat1_5_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({new_AGEMA_signal_7110, mcs1_mcs_mat1_5_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_7266, mcs1_mcs_mat1_5_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7301, shiftr_out[41]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[922]), .c ({new_AGEMA_signal_7960, mcs1_mcs_mat1_5_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[923]), .c ({new_AGEMA_signal_7110, mcs1_mcs_mat1_5_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[924]), .c ({new_AGEMA_signal_7526, mcs1_mcs_mat1_5_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_9769, mcs1_mcs_mat1_5_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_9543, mcs1_mcs_mat1_5_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_9990, mcs1_mcs_mat1_5_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_8918, mcs1_mcs_mat1_5_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_9272, mcs1_mcs_mat1_5_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_10451, mcs1_mcs_mat1_5_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_9770, mcs1_mcs_mat1_5_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_10709, mcs1_mcs_mat1_5_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9362, shiftr_out[9]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[925]), .c ({new_AGEMA_signal_9770, mcs1_mcs_mat1_5_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[926]), .c ({new_AGEMA_signal_8918, mcs1_mcs_mat1_5_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[927]), .c ({new_AGEMA_signal_9543, mcs1_mcs_mat1_5_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_8919, mcs1_mcs_mat1_5_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_8438, mcs1_mcs_mat1_5_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_9273, mcs1_mcs_mat1_5_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_7112, mcs1_mcs_mat1_5_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_8439, mcs1_mcs_mat1_5_mcs_out[29]}), .c ({new_AGEMA_signal_8919, mcs1_mcs_mat1_5_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_7111, mcs1_mcs_mat1_5_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_8438, mcs1_mcs_mat1_5_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_8920, mcs1_mcs_mat1_5_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_7963, mcs1_mcs_mat1_5_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_6610, shiftr_out[104]}), .c ({new_AGEMA_signal_8438, mcs1_mcs_mat1_5_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_8921, mcs1_mcs_mat1_5_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_7961, mcs1_mcs_mat1_5_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_9274, mcs1_mcs_mat1_5_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_8440, mcs1_mcs_mat1_5_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_7962, mcs1_mcs_mat1_5_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_8921, mcs1_mcs_mat1_5_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_7527, mcs1_mcs_mat1_5_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_7962, mcs1_mcs_mat1_5_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_7963, mcs1_mcs_mat1_5_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7112, mcs1_mcs_mat1_5_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_8440, mcs1_mcs_mat1_5_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[928]), .c ({new_AGEMA_signal_7963, mcs1_mcs_mat1_5_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[929]), .c ({new_AGEMA_signal_7112, mcs1_mcs_mat1_5_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[930]), .c ({new_AGEMA_signal_7527, mcs1_mcs_mat1_5_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_7964, mcs1_mcs_mat1_5_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_8441, mcs1_mcs_mat1_5_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_7528, mcs1_mcs_mat1_5_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7113, mcs1_mcs_mat1_5_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_7964, mcs1_mcs_mat1_5_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_8442, mcs1_mcs_mat1_5_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_8922, mcs1_mcs_mat1_5_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_7966, mcs1_mcs_mat1_5_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_7113, mcs1_mcs_mat1_5_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_8442, mcs1_mcs_mat1_5_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_8923, mcs1_mcs_mat1_5_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_6615, shiftr_out[72]}), .c ({new_AGEMA_signal_9275, mcs1_mcs_mat1_5_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_7966, mcs1_mcs_mat1_5_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8443, mcs1_mcs_mat1_5_mcs_out[24]}), .c ({new_AGEMA_signal_8923, mcs1_mcs_mat1_5_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_7965, mcs1_mcs_mat1_5_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_7229, shiftr_out[75]}), .c ({new_AGEMA_signal_8443, mcs1_mcs_mat1_5_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_7528, mcs1_mcs_mat1_5_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_6821, mcs1_mcs_mat1_5_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_7965, mcs1_mcs_mat1_5_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[931]), .c ({new_AGEMA_signal_7966, mcs1_mcs_mat1_5_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[932]), .c ({new_AGEMA_signal_7113, mcs1_mcs_mat1_5_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7229, shiftr_out[75]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[933]), .c ({new_AGEMA_signal_7528, mcs1_mcs_mat1_5_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_7967, mcs1_mcs_mat1_5_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_6689, shiftr_out[42]}), .c ({new_AGEMA_signal_8444, mcs1_mcs_mat1_5_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_7529, mcs1_mcs_mat1_5_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7114, mcs1_mcs_mat1_5_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_7967, mcs1_mcs_mat1_5_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_8445, mcs1_mcs_mat1_5_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_7301, shiftr_out[41]}), .c ({new_AGEMA_signal_8924, mcs1_mcs_mat1_5_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_7969, mcs1_mcs_mat1_5_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_7114, mcs1_mcs_mat1_5_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_8445, mcs1_mcs_mat1_5_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_8925, mcs1_mcs_mat1_5_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_6621, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_9276, mcs1_mcs_mat1_5_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_7969, mcs1_mcs_mat1_5_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8446, mcs1_mcs_mat1_5_mcs_out[20]}), .c ({new_AGEMA_signal_8925, mcs1_mcs_mat1_5_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_7968, mcs1_mcs_mat1_5_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_8446, mcs1_mcs_mat1_5_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_7529, mcs1_mcs_mat1_5_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_6822, mcs1_mcs_mat1_5_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_7968, mcs1_mcs_mat1_5_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7301, shiftr_out[41]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[934]), .c ({new_AGEMA_signal_7969, mcs1_mcs_mat1_5_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[935]), .c ({new_AGEMA_signal_7114, mcs1_mcs_mat1_5_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[936]), .c ({new_AGEMA_signal_7529, mcs1_mcs_mat1_5_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_9771, mcs1_mcs_mat1_5_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_9774, mcs1_mcs_mat1_5_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_9992, mcs1_mcs_mat1_5_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_9993, mcs1_mcs_mat1_5_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_8447, mcs1_mcs_mat1_5_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_10212, mcs1_mcs_mat1_5_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_10213, mcs1_mcs_mat1_5_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_8926, mcs1_mcs_mat1_5_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_10452, mcs1_mcs_mat1_5_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_7620, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_9993, mcs1_mcs_mat1_5_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_10213, mcs1_mcs_mat1_5_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_9772, mcs1_mcs_mat1_5_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_9362, shiftr_out[9]}), .c ({new_AGEMA_signal_9993, mcs1_mcs_mat1_5_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_9544, mcs1_mcs_mat1_5_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_9545, mcs1_mcs_mat1_5_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_9772, mcs1_mcs_mat1_5_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_9773, mcs1_mcs_mat1_5_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_8926, mcs1_mcs_mat1_5_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_9994, mcs1_mcs_mat1_5_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9362, shiftr_out[9]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[937]), .c ({new_AGEMA_signal_9774, mcs1_mcs_mat1_5_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[938]), .c ({new_AGEMA_signal_8926, mcs1_mcs_mat1_5_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[939]), .c ({new_AGEMA_signal_9545, mcs1_mcs_mat1_5_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_8929, mcs1_mcs_mat1_5_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_7267, mcs1_mcs_mat1_5_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_9277, mcs1_mcs_mat1_5_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_8450, mcs1_mcs_mat1_5_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_8448, mcs1_mcs_mat1_5_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_8927, mcs1_mcs_mat1_5_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_7971, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_7115, mcs1_mcs_mat1_5_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8448, mcs1_mcs_mat1_5_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_7267, mcs1_mcs_mat1_5_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_8449, mcs1_mcs_mat1_5_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_8928, mcs1_mcs_mat1_5_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_7970, mcs1_mcs_mat1_5_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_7971, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_8449, mcs1_mcs_mat1_5_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_6823, mcs1_mcs_mat1_5_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_7115, mcs1_mcs_mat1_5_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_7267, mcs1_mcs_mat1_5_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_9278, mcs1_mcs_mat1_5_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_9546, mcs1_mcs_mat1_5_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_8929, mcs1_mcs_mat1_5_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_7971, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_9278, mcs1_mcs_mat1_5_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_8450, mcs1_mcs_mat1_5_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_8929, mcs1_mcs_mat1_5_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_7970, mcs1_mcs_mat1_5_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_8450, mcs1_mcs_mat1_5_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_6610, shiftr_out[104]}), .b ({new_AGEMA_signal_7530, mcs1_mcs_mat1_5_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_7970, mcs1_mcs_mat1_5_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7290, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[940]), .c ({new_AGEMA_signal_7971, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6678, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[941]), .c ({new_AGEMA_signal_7115, mcs1_mcs_mat1_5_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7224, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[942]), .c ({new_AGEMA_signal_7530, mcs1_mcs_mat1_5_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_7268, mcs1_mcs_mat1_5_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_7229, shiftr_out[75]}), .c ({new_AGEMA_signal_7531, mcs1_mcs_mat1_5_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_8452, mcs1_mcs_mat1_5_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_8930, mcs1_mcs_mat1_5_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_7972, mcs1_mcs_mat1_5_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_8451, mcs1_mcs_mat1_5_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_7532, mcs1_mcs_mat1_5_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_7268, mcs1_mcs_mat1_5_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_7972, mcs1_mcs_mat1_5_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_6824, mcs1_mcs_mat1_5_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_7116, mcs1_mcs_mat1_5_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_7268, mcs1_mcs_mat1_5_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_8931, mcs1_mcs_mat1_5_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_6615, shiftr_out[72]}), .c ({new_AGEMA_signal_9279, mcs1_mcs_mat1_5_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_6824, mcs1_mcs_mat1_5_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8452, mcs1_mcs_mat1_5_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_8931, mcs1_mcs_mat1_5_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_7973, mcs1_mcs_mat1_5_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_7532, mcs1_mcs_mat1_5_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_8452, mcs1_mcs_mat1_5_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7295, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[943]), .c ({new_AGEMA_signal_7973, mcs1_mcs_mat1_5_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6683, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[944]), .c ({new_AGEMA_signal_7116, mcs1_mcs_mat1_5_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7229, shiftr_out[75]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[945]), .c ({new_AGEMA_signal_7532, mcs1_mcs_mat1_5_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_9547, mcs1_mcs_mat1_5_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_7534, mcs1_mcs_mat1_5_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_9775, mcs1_mcs_mat1_5_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_9280, mcs1_mcs_mat1_5_mcs_out[7]}), .b ({new_AGEMA_signal_6689, shiftr_out[42]}), .c ({new_AGEMA_signal_9547, mcs1_mcs_mat1_5_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_8932, mcs1_mcs_mat1_5_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_7301, shiftr_out[41]}), .c ({new_AGEMA_signal_9280, mcs1_mcs_mat1_5_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_8453, mcs1_mcs_mat1_5_mcs_out[6]}), .b ({new_AGEMA_signal_7118, mcs1_mcs_mat1_5_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_8932, mcs1_mcs_mat1_5_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_7117, mcs1_mcs_mat1_5_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_7974, mcs1_mcs_mat1_5_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_8453, mcs1_mcs_mat1_5_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7301, shiftr_out[41]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[946]), .c ({new_AGEMA_signal_7974, mcs1_mcs_mat1_5_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6689, shiftr_out[42]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[947]), .c ({new_AGEMA_signal_7118, mcs1_mcs_mat1_5_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7235, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[948]), .c ({new_AGEMA_signal_7534, mcs1_mcs_mat1_5_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_9548, mcs1_mcs_mat1_5_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_9776, mcs1_mcs_mat1_5_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_9996, mcs1_mcs_mat1_5_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_9362, shiftr_out[9]}), .b ({new_AGEMA_signal_9549, mcs1_mcs_mat1_5_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_9776, mcs1_mcs_mat1_5_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_9997, mcs1_mcs_mat1_5_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_8933, mcs1_mcs_mat1_5_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_10214, mcs1_mcs_mat1_5_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_9998, mcs1_mcs_mat1_5_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_9778, mcs1_mcs_mat1_5_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_10215, mcs1_mcs_mat1_5_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_9779, mcs1_mcs_mat1_5_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_8454, mcs1_mcs_mat1_5_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_9998, mcs1_mcs_mat1_5_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9362, shiftr_out[9]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[949]), .c ({new_AGEMA_signal_9779, mcs1_mcs_mat1_5_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8100, shiftr_out[10]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[950]), .c ({new_AGEMA_signal_8933, mcs1_mcs_mat1_5_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9058, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[951]), .c ({new_AGEMA_signal_9549, mcs1_mcs_mat1_5_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U96 ( .a ({new_AGEMA_signal_10710, mcs1_mcs_mat1_6_n128}), .b ({new_AGEMA_signal_9281, mcs1_mcs_mat1_6_n127}), .c ({temp_next_s1[69], temp_next_s0[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U95 ( .a ({new_AGEMA_signal_8969, mcs1_mcs_mat1_6_mcs_out[41]}), .b ({new_AGEMA_signal_8006, mcs1_mcs_mat1_6_mcs_out[45]}), .c ({new_AGEMA_signal_9281, mcs1_mcs_mat1_6_n127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U94 ( .a ({new_AGEMA_signal_7270, mcs1_mcs_mat1_6_mcs_out[33]}), .b ({new_AGEMA_signal_10475, mcs1_mcs_mat1_6_mcs_out[37]}), .c ({new_AGEMA_signal_10710, mcs1_mcs_mat1_6_n128}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U93 ( .a ({new_AGEMA_signal_10216, mcs1_mcs_mat1_6_n126}), .b ({new_AGEMA_signal_9780, mcs1_mcs_mat1_6_n125}), .c ({temp_next_s1[68], temp_next_s0[68]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U92 ( .a ({new_AGEMA_signal_8492, mcs1_mcs_mat1_6_mcs_out[40]}), .b ({new_AGEMA_signal_9574, mcs1_mcs_mat1_6_mcs_out[44]}), .c ({new_AGEMA_signal_9780, mcs1_mcs_mat1_6_n125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U91 ( .a ({new_AGEMA_signal_9578, mcs1_mcs_mat1_6_mcs_out[32]}), .b ({new_AGEMA_signal_10015, mcs1_mcs_mat1_6_mcs_out[36]}), .c ({new_AGEMA_signal_10216, mcs1_mcs_mat1_6_n126}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U90 ( .a ({new_AGEMA_signal_10217, mcs1_mcs_mat1_6_n124}), .b ({new_AGEMA_signal_9550, mcs1_mcs_mat1_6_n123}), .c ({temp_next_s1[39], temp_next_s0[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U89 ( .a ({new_AGEMA_signal_8499, mcs1_mcs_mat1_6_mcs_out[27]}), .b ({new_AGEMA_signal_9311, mcs1_mcs_mat1_6_mcs_out[31]}), .c ({new_AGEMA_signal_9550, mcs1_mcs_mat1_6_n123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U88 ( .a ({new_AGEMA_signal_8503, mcs1_mcs_mat1_6_mcs_out[19]}), .b ({new_AGEMA_signal_10016, mcs1_mcs_mat1_6_mcs_out[23]}), .c ({new_AGEMA_signal_10217, mcs1_mcs_mat1_6_n124}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U87 ( .a ({new_AGEMA_signal_10455, mcs1_mcs_mat1_6_n122}), .b ({new_AGEMA_signal_9282, mcs1_mcs_mat1_6_n121}), .c ({temp_next_s1[38], temp_next_s0[38]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U86 ( .a ({new_AGEMA_signal_8975, mcs1_mcs_mat1_6_mcs_out[26]}), .b ({new_AGEMA_signal_8973, mcs1_mcs_mat1_6_mcs_out[30]}), .c ({new_AGEMA_signal_9282, mcs1_mcs_mat1_6_n121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U85 ( .a ({new_AGEMA_signal_8978, mcs1_mcs_mat1_6_mcs_out[18]}), .b ({new_AGEMA_signal_10238, mcs1_mcs_mat1_6_mcs_out[22]}), .c ({new_AGEMA_signal_10455, mcs1_mcs_mat1_6_n122}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U84 ( .a ({new_AGEMA_signal_10712, mcs1_mcs_mat1_6_n120}), .b ({new_AGEMA_signal_9551, mcs1_mcs_mat1_6_n119}), .c ({temp_next_s1[37], temp_next_s0[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U83 ( .a ({new_AGEMA_signal_9313, mcs1_mcs_mat1_6_mcs_out[25]}), .b ({new_AGEMA_signal_8497, mcs1_mcs_mat1_6_mcs_out[29]}), .c ({new_AGEMA_signal_9551, mcs1_mcs_mat1_6_n119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U82 ( .a ({new_AGEMA_signal_9314, mcs1_mcs_mat1_6_mcs_out[17]}), .b ({new_AGEMA_signal_10476, mcs1_mcs_mat1_6_mcs_out[21]}), .c ({new_AGEMA_signal_10712, mcs1_mcs_mat1_6_n120}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U81 ( .a ({new_AGEMA_signal_10218, mcs1_mcs_mat1_6_n118}), .b ({new_AGEMA_signal_9552, mcs1_mcs_mat1_6_n117}), .c ({temp_next_s1[36], temp_next_s0[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U80 ( .a ({new_AGEMA_signal_8501, mcs1_mcs_mat1_6_mcs_out[24]}), .b ({new_AGEMA_signal_9312, mcs1_mcs_mat1_6_mcs_out[28]}), .c ({new_AGEMA_signal_9552, mcs1_mcs_mat1_6_n117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U79 ( .a ({new_AGEMA_signal_8505, mcs1_mcs_mat1_6_mcs_out[16]}), .b ({new_AGEMA_signal_10018, mcs1_mcs_mat1_6_mcs_out[20]}), .c ({new_AGEMA_signal_10218, mcs1_mcs_mat1_6_n118}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U78 ( .a ({new_AGEMA_signal_9553, mcs1_mcs_mat1_6_n116}), .b ({new_AGEMA_signal_10713, mcs1_mcs_mat1_6_n115}), .c ({temp_next_s1[7], temp_next_s0[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U77 ( .a ({new_AGEMA_signal_8512, mcs1_mcs_mat1_6_mcs_out[3]}), .b ({new_AGEMA_signal_10477, mcs1_mcs_mat1_6_mcs_out[7]}), .c ({new_AGEMA_signal_10713, mcs1_mcs_mat1_6_n115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U76 ( .a ({new_AGEMA_signal_7566, mcs1_mcs_mat1_6_mcs_out[11]}), .b ({new_AGEMA_signal_9315, mcs1_mcs_mat1_6_mcs_out[15]}), .c ({new_AGEMA_signal_9553, mcs1_mcs_mat1_6_n116}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U75 ( .a ({new_AGEMA_signal_10714, mcs1_mcs_mat1_6_n114}), .b ({new_AGEMA_signal_9554, mcs1_mcs_mat1_6_n113}), .c ({new_AGEMA_signal_10923, mcs_out[231]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U74 ( .a ({new_AGEMA_signal_9292, mcs1_mcs_mat1_6_mcs_out[123]}), .b ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_9554, mcs1_mcs_mat1_6_n113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U73 ( .a ({new_AGEMA_signal_8942, mcs1_mcs_mat1_6_mcs_out[115]}), .b ({new_AGEMA_signal_10468, mcs1_mcs_mat1_6_mcs_out[119]}), .c ({new_AGEMA_signal_10714, mcs1_mcs_mat1_6_n114}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U72 ( .a ({new_AGEMA_signal_10715, mcs1_mcs_mat1_6_n112}), .b ({new_AGEMA_signal_8455, mcs1_mcs_mat1_6_n111}), .c ({new_AGEMA_signal_10924, mcs_out[230]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U71 ( .a ({new_AGEMA_signal_7975, mcs1_mcs_mat1_6_mcs_out[122]}), .b ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_8455, mcs1_mcs_mat1_6_n111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U70 ( .a ({new_AGEMA_signal_8461, mcs1_mcs_mat1_6_mcs_out[114]}), .b ({new_AGEMA_signal_10469, mcs1_mcs_mat1_6_mcs_out[118]}), .c ({new_AGEMA_signal_10715, mcs1_mcs_mat1_6_n112}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U69 ( .a ({new_AGEMA_signal_9283, mcs1_mcs_mat1_6_n110}), .b ({new_AGEMA_signal_10219, mcs1_mcs_mat1_6_n109}), .c ({temp_next_s1[6], temp_next_s0[6]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U68 ( .a ({new_AGEMA_signal_8513, mcs1_mcs_mat1_6_mcs_out[2]}), .b ({new_AGEMA_signal_10019, mcs1_mcs_mat1_6_mcs_out[6]}), .c ({new_AGEMA_signal_10219, mcs1_mcs_mat1_6_n109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U67 ( .a ({new_AGEMA_signal_8983, mcs1_mcs_mat1_6_mcs_out[10]}), .b ({new_AGEMA_signal_8980, mcs1_mcs_mat1_6_mcs_out[14]}), .c ({new_AGEMA_signal_9283, mcs1_mcs_mat1_6_n110}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U66 ( .a ({new_AGEMA_signal_10458, mcs1_mcs_mat1_6_n108}), .b ({new_AGEMA_signal_9555, mcs1_mcs_mat1_6_n107}), .c ({new_AGEMA_signal_10716, mcs_out[229]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U65 ( .a ({new_AGEMA_signal_9293, mcs1_mcs_mat1_6_mcs_out[121]}), .b ({new_AGEMA_signal_7535, mcs1_mcs_mat1_6_mcs_out[125]}), .c ({new_AGEMA_signal_9555, mcs1_mcs_mat1_6_n107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U64 ( .a ({new_AGEMA_signal_7977, mcs1_mcs_mat1_6_mcs_out[113]}), .b ({new_AGEMA_signal_10228, mcs1_mcs_mat1_6_mcs_out[117]}), .c ({new_AGEMA_signal_10458, mcs1_mcs_mat1_6_n108}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U63 ( .a ({new_AGEMA_signal_10220, mcs1_mcs_mat1_6_n106}), .b ({new_AGEMA_signal_9284, mcs1_mcs_mat1_6_n105}), .c ({new_AGEMA_signal_10459, mcs_out[228]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U62 ( .a ({new_AGEMA_signal_8940, mcs1_mcs_mat1_6_mcs_out[120]}), .b ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_9284, mcs1_mcs_mat1_6_n105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U61 ( .a ({new_AGEMA_signal_9294, mcs1_mcs_mat1_6_mcs_out[112]}), .b ({new_AGEMA_signal_10005, mcs1_mcs_mat1_6_mcs_out[116]}), .c ({new_AGEMA_signal_10220, mcs1_mcs_mat1_6_n106}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U60 ( .a ({new_AGEMA_signal_10460, mcs1_mcs_mat1_6_n104}), .b ({new_AGEMA_signal_9556, mcs1_mcs_mat1_6_n103}), .c ({new_AGEMA_signal_10717, mcs_out[199]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U59 ( .a ({new_AGEMA_signal_9295, mcs1_mcs_mat1_6_mcs_out[111]}), .b ({new_AGEMA_signal_9300, mcs1_mcs_mat1_6_mcs_out[99]}), .c ({new_AGEMA_signal_9556, mcs1_mcs_mat1_6_n103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U58 ( .a ({new_AGEMA_signal_10229, mcs1_mcs_mat1_6_mcs_out[103]}), .b ({new_AGEMA_signal_8946, mcs1_mcs_mat1_6_mcs_out[107]}), .c ({new_AGEMA_signal_10460, mcs1_mcs_mat1_6_n104}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U57 ( .a ({new_AGEMA_signal_9999, mcs1_mcs_mat1_6_n102}), .b ({new_AGEMA_signal_9557, mcs1_mcs_mat1_6_n101}), .c ({new_AGEMA_signal_10221, mcs_out[198]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U56 ( .a ({new_AGEMA_signal_9296, mcs1_mcs_mat1_6_mcs_out[110]}), .b ({new_AGEMA_signal_8469, mcs1_mcs_mat1_6_mcs_out[98]}), .c ({new_AGEMA_signal_9557, mcs1_mcs_mat1_6_n101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U55 ( .a ({new_AGEMA_signal_9787, mcs1_mcs_mat1_6_mcs_out[102]}), .b ({new_AGEMA_signal_8947, mcs1_mcs_mat1_6_mcs_out[106]}), .c ({new_AGEMA_signal_9999, mcs1_mcs_mat1_6_n102}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U54 ( .a ({new_AGEMA_signal_10222, mcs1_mcs_mat1_6_n100}), .b ({new_AGEMA_signal_9558, mcs1_mcs_mat1_6_n99}), .c ({new_AGEMA_signal_10461, mcs_out[197]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U53 ( .a ({new_AGEMA_signal_9297, mcs1_mcs_mat1_6_mcs_out[109]}), .b ({new_AGEMA_signal_7543, mcs1_mcs_mat1_6_mcs_out[97]}), .c ({new_AGEMA_signal_9558, mcs1_mcs_mat1_6_n99}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U52 ( .a ({new_AGEMA_signal_10007, mcs1_mcs_mat1_6_mcs_out[101]}), .b ({new_AGEMA_signal_8948, mcs1_mcs_mat1_6_mcs_out[105]}), .c ({new_AGEMA_signal_10222, mcs1_mcs_mat1_6_n100}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U51 ( .a ({new_AGEMA_signal_10462, mcs1_mcs_mat1_6_n98}), .b ({new_AGEMA_signal_10000, mcs1_mcs_mat1_6_n97}), .c ({new_AGEMA_signal_10718, mcs_out[196]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U50 ( .a ({new_AGEMA_signal_9298, mcs1_mcs_mat1_6_mcs_out[108]}), .b ({new_AGEMA_signal_9791, mcs1_mcs_mat1_6_mcs_out[96]}), .c ({new_AGEMA_signal_10000, mcs1_mcs_mat1_6_n97}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U49 ( .a ({new_AGEMA_signal_10230, mcs1_mcs_mat1_6_mcs_out[100]}), .b ({new_AGEMA_signal_9299, mcs1_mcs_mat1_6_mcs_out[104]}), .c ({new_AGEMA_signal_10462, mcs1_mcs_mat1_6_n98}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U48 ( .a ({new_AGEMA_signal_10001, mcs1_mcs_mat1_6_n96}), .b ({new_AGEMA_signal_9285, mcs1_mcs_mat1_6_n95}), .c ({new_AGEMA_signal_10223, mcs_out[167]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U47 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_8952, mcs1_mcs_mat1_6_mcs_out[95]}), .c ({new_AGEMA_signal_9285, mcs1_mcs_mat1_6_n95}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U46 ( .a ({new_AGEMA_signal_8471, mcs1_mcs_mat1_6_mcs_out[83]}), .b ({new_AGEMA_signal_9792, mcs1_mcs_mat1_6_mcs_out[87]}), .c ({new_AGEMA_signal_10001, mcs1_mcs_mat1_6_n96}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U45 ( .a ({new_AGEMA_signal_8934, mcs1_mcs_mat1_6_n94}), .b ({new_AGEMA_signal_8456, mcs1_mcs_mat1_6_n93}), .c ({new_AGEMA_signal_9286, mcs_out[166]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U43 ( .a ({new_AGEMA_signal_8472, mcs1_mcs_mat1_6_mcs_out[82]}), .b ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_8934, mcs1_mcs_mat1_6_n94}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U42 ( .a ({new_AGEMA_signal_9559, mcs1_mcs_mat1_6_n92}), .b ({new_AGEMA_signal_8457, mcs1_mcs_mat1_6_n91}), .c ({new_AGEMA_signal_9781, mcs_out[165]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U41 ( .a ({new_AGEMA_signal_7549, mcs1_mcs_mat1_6_mcs_out[89]}), .b ({new_AGEMA_signal_7986, mcs1_mcs_mat1_6_mcs_out[93]}), .c ({new_AGEMA_signal_8457, mcs1_mcs_mat1_6_n91}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U40 ( .a ({new_AGEMA_signal_8473, mcs1_mcs_mat1_6_mcs_out[81]}), .b ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_9559, mcs1_mcs_mat1_6_n92}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U39 ( .a ({new_AGEMA_signal_10224, mcs1_mcs_mat1_6_n90}), .b ({new_AGEMA_signal_9560, mcs1_mcs_mat1_6_n89}), .c ({new_AGEMA_signal_10463, mcs_out[164]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U38 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_9301, mcs1_mcs_mat1_6_mcs_out[92]}), .c ({new_AGEMA_signal_9560, mcs1_mcs_mat1_6_n89}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U37 ( .a ({new_AGEMA_signal_8954, mcs1_mcs_mat1_6_mcs_out[80]}), .b ({new_AGEMA_signal_10009, mcs1_mcs_mat1_6_mcs_out[84]}), .c ({new_AGEMA_signal_10224, mcs1_mcs_mat1_6_n90}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U36 ( .a ({new_AGEMA_signal_9287, mcs1_mcs_mat1_6_n88}), .b ({new_AGEMA_signal_9782, mcs1_mcs_mat1_6_n87}), .c ({temp_next_s1[5], temp_next_s0[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U35 ( .a ({new_AGEMA_signal_9581, mcs1_mcs_mat1_6_mcs_out[5]}), .b ({new_AGEMA_signal_8509, mcs1_mcs_mat1_6_mcs_out[9]}), .c ({new_AGEMA_signal_9782, mcs1_mcs_mat1_6_n87}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U34 ( .a ({new_AGEMA_signal_8981, mcs1_mcs_mat1_6_mcs_out[13]}), .b ({new_AGEMA_signal_8987, mcs1_mcs_mat1_6_mcs_out[1]}), .c ({new_AGEMA_signal_9287, mcs1_mcs_mat1_6_n88}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U33 ( .a ({new_AGEMA_signal_10464, mcs1_mcs_mat1_6_n86}), .b ({new_AGEMA_signal_9288, mcs1_mcs_mat1_6_n85}), .c ({new_AGEMA_signal_10719, mcs_out[135]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U32 ( .a ({new_AGEMA_signal_7994, mcs1_mcs_mat1_6_mcs_out[75]}), .b ({new_AGEMA_signal_8955, mcs1_mcs_mat1_6_mcs_out[79]}), .c ({new_AGEMA_signal_9288, mcs1_mcs_mat1_6_n85}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U31 ( .a ({new_AGEMA_signal_9305, mcs1_mcs_mat1_6_mcs_out[67]}), .b ({new_AGEMA_signal_10231, mcs1_mcs_mat1_6_mcs_out[71]}), .c ({new_AGEMA_signal_10464, mcs1_mcs_mat1_6_n86}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U30 ( .a ({new_AGEMA_signal_10720, mcs1_mcs_mat1_6_n84}), .b ({new_AGEMA_signal_9561, mcs1_mcs_mat1_6_n83}), .c ({new_AGEMA_signal_10925, mcs_out[134]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U29 ( .a ({new_AGEMA_signal_9303, mcs1_mcs_mat1_6_mcs_out[74]}), .b ({new_AGEMA_signal_7129, mcs1_mcs_mat1_6_mcs_out[78]}), .c ({new_AGEMA_signal_9561, mcs1_mcs_mat1_6_n83}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U28 ( .a ({new_AGEMA_signal_8960, mcs1_mcs_mat1_6_mcs_out[66]}), .b ({new_AGEMA_signal_10470, mcs1_mcs_mat1_6_mcs_out[70]}), .c ({new_AGEMA_signal_10720, mcs1_mcs_mat1_6_n84}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U27 ( .a ({new_AGEMA_signal_10721, mcs1_mcs_mat1_6_n82}), .b ({new_AGEMA_signal_8935, mcs1_mcs_mat1_6_n81}), .c ({new_AGEMA_signal_10926, mcs_out[133]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U26 ( .a ({new_AGEMA_signal_8476, mcs1_mcs_mat1_6_mcs_out[73]}), .b ({new_AGEMA_signal_7992, mcs1_mcs_mat1_6_mcs_out[77]}), .c ({new_AGEMA_signal_8935, mcs1_mcs_mat1_6_n81}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U25 ( .a ({new_AGEMA_signal_7997, mcs1_mcs_mat1_6_mcs_out[65]}), .b ({new_AGEMA_signal_10471, mcs1_mcs_mat1_6_mcs_out[69]}), .c ({new_AGEMA_signal_10721, mcs1_mcs_mat1_6_n82}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U24 ( .a ({new_AGEMA_signal_10465, mcs1_mcs_mat1_6_n80}), .b ({new_AGEMA_signal_9562, mcs1_mcs_mat1_6_n79}), .c ({new_AGEMA_signal_10722, mcs_out[132]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U23 ( .a ({new_AGEMA_signal_9304, mcs1_mcs_mat1_6_mcs_out[72]}), .b ({new_AGEMA_signal_9302, mcs1_mcs_mat1_6_mcs_out[76]}), .c ({new_AGEMA_signal_9562, mcs1_mcs_mat1_6_n79}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U22 ( .a ({new_AGEMA_signal_9572, mcs1_mcs_mat1_6_mcs_out[64]}), .b ({new_AGEMA_signal_10233, mcs1_mcs_mat1_6_mcs_out[68]}), .c ({new_AGEMA_signal_10465, mcs1_mcs_mat1_6_n80}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U21 ( .a ({new_AGEMA_signal_10466, mcs1_mcs_mat1_6_n78}), .b ({new_AGEMA_signal_9289, mcs1_mcs_mat1_6_n77}), .c ({temp_next_s1[103], temp_next_s0[103]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U20 ( .a ({new_AGEMA_signal_8483, mcs1_mcs_mat1_6_mcs_out[59]}), .b ({new_AGEMA_signal_8962, mcs1_mcs_mat1_6_mcs_out[63]}), .c ({new_AGEMA_signal_9289, mcs1_mcs_mat1_6_n77}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U19 ( .a ({new_AGEMA_signal_8005, mcs1_mcs_mat1_6_mcs_out[51]}), .b ({new_AGEMA_signal_10234, mcs1_mcs_mat1_6_mcs_out[55]}), .c ({new_AGEMA_signal_10466, mcs1_mcs_mat1_6_n78}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U18 ( .a ({new_AGEMA_signal_10724, mcs1_mcs_mat1_6_n76}), .b ({new_AGEMA_signal_8936, mcs1_mcs_mat1_6_n75}), .c ({temp_next_s1[102], temp_next_s0[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U17 ( .a ({new_AGEMA_signal_8001, mcs1_mcs_mat1_6_mcs_out[58]}), .b ({new_AGEMA_signal_8480, mcs1_mcs_mat1_6_mcs_out[62]}), .c ({new_AGEMA_signal_8936, mcs1_mcs_mat1_6_n75}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U16 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_10472, mcs1_mcs_mat1_6_mcs_out[54]}), .c ({new_AGEMA_signal_10724, mcs1_mcs_mat1_6_n76}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U15 ( .a ({new_AGEMA_signal_10725, mcs1_mcs_mat1_6_n74}), .b ({new_AGEMA_signal_8937, mcs1_mcs_mat1_6_n73}), .c ({temp_next_s1[101], temp_next_s0[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U14 ( .a ({new_AGEMA_signal_8484, mcs1_mcs_mat1_6_mcs_out[57]}), .b ({new_AGEMA_signal_8481, mcs1_mcs_mat1_6_mcs_out[61]}), .c ({new_AGEMA_signal_8937, mcs1_mcs_mat1_6_n73}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U13 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_10473, mcs1_mcs_mat1_6_mcs_out[53]}), .c ({new_AGEMA_signal_10725, mcs1_mcs_mat1_6_n74}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U12 ( .a ({new_AGEMA_signal_10467, mcs1_mcs_mat1_6_n72}), .b ({new_AGEMA_signal_9563, mcs1_mcs_mat1_6_n71}), .c ({temp_next_s1[100], temp_next_s0[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U11 ( .a ({new_AGEMA_signal_8964, mcs1_mcs_mat1_6_mcs_out[56]}), .b ({new_AGEMA_signal_9307, mcs1_mcs_mat1_6_mcs_out[60]}), .c ({new_AGEMA_signal_9563, mcs1_mcs_mat1_6_n71}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U10 ( .a ({new_AGEMA_signal_8487, mcs1_mcs_mat1_6_mcs_out[48]}), .b ({new_AGEMA_signal_10236, mcs1_mcs_mat1_6_mcs_out[52]}), .c ({new_AGEMA_signal_10467, mcs1_mcs_mat1_6_n72}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U9 ( .a ({new_AGEMA_signal_10727, mcs1_mcs_mat1_6_n70}), .b ({new_AGEMA_signal_9290, mcs1_mcs_mat1_6_n69}), .c ({temp_next_s1[71], temp_next_s0[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U8 ( .a ({new_AGEMA_signal_8967, mcs1_mcs_mat1_6_mcs_out[43]}), .b ({new_AGEMA_signal_8966, mcs1_mcs_mat1_6_mcs_out[47]}), .c ({new_AGEMA_signal_9290, mcs1_mcs_mat1_6_n69}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U7 ( .a ({new_AGEMA_signal_8971, mcs1_mcs_mat1_6_mcs_out[35]}), .b ({new_AGEMA_signal_10474, mcs1_mcs_mat1_6_mcs_out[39]}), .c ({new_AGEMA_signal_10727, mcs1_mcs_mat1_6_n70}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U6 ( .a ({new_AGEMA_signal_10003, mcs1_mcs_mat1_6_n68}), .b ({new_AGEMA_signal_9291, mcs1_mcs_mat1_6_n67}), .c ({temp_next_s1[70], temp_next_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U5 ( .a ({new_AGEMA_signal_8968, mcs1_mcs_mat1_6_mcs_out[42]}), .b ({new_AGEMA_signal_7556, mcs1_mcs_mat1_6_mcs_out[46]}), .c ({new_AGEMA_signal_9291, mcs1_mcs_mat1_6_n67}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U4 ( .a ({new_AGEMA_signal_8494, mcs1_mcs_mat1_6_mcs_out[34]}), .b ({new_AGEMA_signal_9800, mcs1_mcs_mat1_6_mcs_out[38]}), .c ({new_AGEMA_signal_10003, mcs1_mcs_mat1_6_n68}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U3 ( .a ({new_AGEMA_signal_9783, mcs1_mcs_mat1_6_n66}), .b ({new_AGEMA_signal_11055, mcs1_mcs_mat1_6_n65}), .c ({temp_next_s1[4], temp_next_s0[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U2 ( .a ({new_AGEMA_signal_10930, mcs1_mcs_mat1_6_mcs_out[4]}), .b ({new_AGEMA_signal_9317, mcs1_mcs_mat1_6_mcs_out[8]}), .c ({new_AGEMA_signal_11055, mcs1_mcs_mat1_6_n65}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_U1 ( .a ({new_AGEMA_signal_8988, mcs1_mcs_mat1_6_mcs_out[0]}), .b ({new_AGEMA_signal_9580, mcs1_mcs_mat1_6_mcs_out[12]}), .c ({new_AGEMA_signal_9783, mcs1_mcs_mat1_6_n66}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_8938, mcs1_mcs_mat1_6_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_9292, mcs1_mcs_mat1_6_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_8458, mcs1_mcs_mat1_6_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_6826, mcs1_mcs_mat1_6_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8938, mcs1_mcs_mat1_6_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_7119, mcs1_mcs_mat1_6_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_7536, mcs1_mcs_mat1_6_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_7975, mcs1_mcs_mat1_6_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_7120, mcs1_mcs_mat1_6_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_7228, shiftr_out[71]}), .c ({new_AGEMA_signal_7536, mcs1_mcs_mat1_6_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_8939, mcs1_mcs_mat1_6_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_7228, shiftr_out[71]}), .c ({new_AGEMA_signal_9293, mcs1_mcs_mat1_6_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_8458, mcs1_mcs_mat1_6_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_8939, mcs1_mcs_mat1_6_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_7976, mcs1_mcs_mat1_6_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_7537, mcs1_mcs_mat1_6_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_8458, mcs1_mcs_mat1_6_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_8459, mcs1_mcs_mat1_6_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_8940, mcs1_mcs_mat1_6_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_7976, mcs1_mcs_mat1_6_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_7120, mcs1_mcs_mat1_6_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_8459, mcs1_mcs_mat1_6_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[952]), .c ({new_AGEMA_signal_7976, mcs1_mcs_mat1_6_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[953]), .c ({new_AGEMA_signal_7120, mcs1_mcs_mat1_6_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7228, shiftr_out[71]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[954]), .c ({new_AGEMA_signal_7537, mcs1_mcs_mat1_6_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_10226, mcs1_mcs_mat1_6_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_8098, shiftr_out[38]}), .c ({new_AGEMA_signal_10468, mcs1_mcs_mat1_6_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_10004, mcs1_mcs_mat1_6_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9566, mcs1_mcs_mat1_6_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_10226, mcs1_mcs_mat1_6_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_10227, mcs1_mcs_mat1_6_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_9785, mcs1_mcs_mat1_6_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_10469, mcs1_mcs_mat1_6_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_10004, mcs1_mcs_mat1_6_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9360, shiftr_out[37]}), .c ({new_AGEMA_signal_10227, mcs1_mcs_mat1_6_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_10004, mcs1_mcs_mat1_6_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9784, mcs1_mcs_mat1_6_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_10228, mcs1_mcs_mat1_6_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_9786, mcs1_mcs_mat1_6_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_8941, mcs1_mcs_mat1_6_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_10004, mcs1_mcs_mat1_6_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_9565, mcs1_mcs_mat1_6_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_9785, mcs1_mcs_mat1_6_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_10005, mcs1_mcs_mat1_6_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_8460, mcs1_mcs_mat1_6_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_9566, mcs1_mcs_mat1_6_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_9785, mcs1_mcs_mat1_6_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_8941, mcs1_mcs_mat1_6_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_9565, mcs1_mcs_mat1_6_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9360, shiftr_out[37]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[955]), .c ({new_AGEMA_signal_9786, mcs1_mcs_mat1_6_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[956]), .c ({new_AGEMA_signal_8941, mcs1_mcs_mat1_6_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[957]), .c ({new_AGEMA_signal_9566, mcs1_mcs_mat1_6_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_8462, mcs1_mcs_mat1_6_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_7121, mcs1_mcs_mat1_6_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_8942, mcs1_mcs_mat1_6_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_7538, mcs1_mcs_mat1_6_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_7539, mcs1_mcs_mat1_6_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_7977, mcs1_mcs_mat1_6_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_8463, mcs1_mcs_mat1_6_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_8943, mcs1_mcs_mat1_6_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_9294, mcs1_mcs_mat1_6_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_8462, mcs1_mcs_mat1_6_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_8943, mcs1_mcs_mat1_6_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_6827, mcs1_mcs_mat1_6_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_7979, mcs1_mcs_mat1_6_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_8462, mcs1_mcs_mat1_6_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_7122, mcs1_mcs_mat1_6_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_7978, mcs1_mcs_mat1_6_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8463, mcs1_mcs_mat1_6_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7307, shiftr_out[5]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[958]), .c ({new_AGEMA_signal_7979, mcs1_mcs_mat1_6_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[959]), .c ({new_AGEMA_signal_7122, mcs1_mcs_mat1_6_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[960]), .c ({new_AGEMA_signal_7539, mcs1_mcs_mat1_6_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({new_AGEMA_signal_8944, mcs1_mcs_mat1_6_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9295, mcs1_mcs_mat1_6_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({new_AGEMA_signal_8945, mcs1_mcs_mat1_6_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9296, mcs1_mcs_mat1_6_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_7540, mcs1_mcs_mat1_6_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_8944, mcs1_mcs_mat1_6_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9297, mcs1_mcs_mat1_6_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_7123, mcs1_mcs_mat1_6_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_8464, mcs1_mcs_mat1_6_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_8944, mcs1_mcs_mat1_6_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_7980, mcs1_mcs_mat1_6_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8945, mcs1_mcs_mat1_6_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9298, mcs1_mcs_mat1_6_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_8465, mcs1_mcs_mat1_6_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_8945, mcs1_mcs_mat1_6_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_7540, mcs1_mcs_mat1_6_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_7981, mcs1_mcs_mat1_6_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_8465, mcs1_mcs_mat1_6_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[961]), .c ({new_AGEMA_signal_7981, mcs1_mcs_mat1_6_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[962]), .c ({new_AGEMA_signal_7123, mcs1_mcs_mat1_6_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[963]), .c ({new_AGEMA_signal_7540, mcs1_mcs_mat1_6_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_8467, mcs1_mcs_mat1_6_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_8466, mcs1_mcs_mat1_6_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8946, mcs1_mcs_mat1_6_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_8466, mcs1_mcs_mat1_6_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_7541, mcs1_mcs_mat1_6_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_8947, mcs1_mcs_mat1_6_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_7124, mcs1_mcs_mat1_6_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7228, shiftr_out[71]}), .c ({new_AGEMA_signal_7541, mcs1_mcs_mat1_6_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_8466, mcs1_mcs_mat1_6_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_8948, mcs1_mcs_mat1_6_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_7983, mcs1_mcs_mat1_6_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_6829, mcs1_mcs_mat1_6_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_8466, mcs1_mcs_mat1_6_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_8949, mcs1_mcs_mat1_6_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_9299, mcs1_mcs_mat1_6_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_8467, mcs1_mcs_mat1_6_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_7983, mcs1_mcs_mat1_6_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_8949, mcs1_mcs_mat1_6_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_7982, mcs1_mcs_mat1_6_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_6614, shiftr_out[68]}), .c ({new_AGEMA_signal_8467, mcs1_mcs_mat1_6_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_7124, mcs1_mcs_mat1_6_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_7542, mcs1_mcs_mat1_6_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_7982, mcs1_mcs_mat1_6_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[964]), .c ({new_AGEMA_signal_7983, mcs1_mcs_mat1_6_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[965]), .c ({new_AGEMA_signal_7124, mcs1_mcs_mat1_6_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7228, shiftr_out[71]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[966]), .c ({new_AGEMA_signal_7542, mcs1_mcs_mat1_6_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_9567, mcs1_mcs_mat1_6_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_10006, mcs1_mcs_mat1_6_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_10229, mcs1_mcs_mat1_6_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_9790, mcs1_mcs_mat1_6_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_10006, mcs1_mcs_mat1_6_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_9788, mcs1_mcs_mat1_6_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_9568, mcs1_mcs_mat1_6_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_10007, mcs1_mcs_mat1_6_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_9789, mcs1_mcs_mat1_6_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_10008, mcs1_mcs_mat1_6_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_10230, mcs1_mcs_mat1_6_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_8468, mcs1_mcs_mat1_6_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_9790, mcs1_mcs_mat1_6_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_10008, mcs1_mcs_mat1_6_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_8950, mcs1_mcs_mat1_6_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_9360, shiftr_out[37]}), .c ({new_AGEMA_signal_9789, mcs1_mcs_mat1_6_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9360, shiftr_out[37]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[967]), .c ({new_AGEMA_signal_9790, mcs1_mcs_mat1_6_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[968]), .c ({new_AGEMA_signal_8950, mcs1_mcs_mat1_6_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[969]), .c ({new_AGEMA_signal_9568, mcs1_mcs_mat1_6_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_9569, mcs1_mcs_mat1_6_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_7544, mcs1_mcs_mat1_6_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_9791, mcs1_mcs_mat1_6_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_9300, mcs1_mcs_mat1_6_mcs_out[99]}), .b ({new_AGEMA_signal_6695, shiftr_out[6]}), .c ({new_AGEMA_signal_9569, mcs1_mcs_mat1_6_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_8951, mcs1_mcs_mat1_6_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_7307, shiftr_out[5]}), .c ({new_AGEMA_signal_9300, mcs1_mcs_mat1_6_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_8469, mcs1_mcs_mat1_6_mcs_out[98]}), .b ({new_AGEMA_signal_7126, mcs1_mcs_mat1_6_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_8951, mcs1_mcs_mat1_6_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_7125, mcs1_mcs_mat1_6_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_7984, mcs1_mcs_mat1_6_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_8469, mcs1_mcs_mat1_6_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7307, shiftr_out[5]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[970]), .c ({new_AGEMA_signal_7984, mcs1_mcs_mat1_6_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[971]), .c ({new_AGEMA_signal_7126, mcs1_mcs_mat1_6_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[972]), .c ({new_AGEMA_signal_7544, mcs1_mcs_mat1_6_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_8470, mcs1_mcs_mat1_6_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_8952, mcs1_mcs_mat1_6_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_7546, mcs1_mcs_mat1_6_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_7547, mcs1_mcs_mat1_6_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_7986, mcs1_mcs_mat1_6_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_8953, mcs1_mcs_mat1_6_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_7127, mcs1_mcs_mat1_6_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_9301, mcs1_mcs_mat1_6_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_8470, mcs1_mcs_mat1_6_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_8953, mcs1_mcs_mat1_6_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_6831, mcs1_mcs_mat1_6_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_7987, mcs1_mcs_mat1_6_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_8470, mcs1_mcs_mat1_6_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[973]), .c ({new_AGEMA_signal_7987, mcs1_mcs_mat1_6_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[974]), .c ({new_AGEMA_signal_7127, mcs1_mcs_mat1_6_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[975]), .c ({new_AGEMA_signal_7547, mcs1_mcs_mat1_6_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_7990, mcs1_mcs_mat1_6_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_7991, mcs1_mcs_mat1_6_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_8471, mcs1_mcs_mat1_6_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_7988, mcs1_mcs_mat1_6_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_6832, mcs1_mcs_mat1_6_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_8472, mcs1_mcs_mat1_6_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_7550, mcs1_mcs_mat1_6_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_7988, mcs1_mcs_mat1_6_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_7989, mcs1_mcs_mat1_6_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_8473, mcs1_mcs_mat1_6_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_7128, mcs1_mcs_mat1_6_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_7550, mcs1_mcs_mat1_6_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_7989, mcs1_mcs_mat1_6_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_8474, mcs1_mcs_mat1_6_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_6695, shiftr_out[6]}), .c ({new_AGEMA_signal_8954, mcs1_mcs_mat1_6_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_7990, mcs1_mcs_mat1_6_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_7128, mcs1_mcs_mat1_6_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_8474, mcs1_mcs_mat1_6_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7307, shiftr_out[5]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[976]), .c ({new_AGEMA_signal_7991, mcs1_mcs_mat1_6_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[977]), .c ({new_AGEMA_signal_7128, mcs1_mcs_mat1_6_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[978]), .c ({new_AGEMA_signal_7550, mcs1_mcs_mat1_6_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_8475, mcs1_mcs_mat1_6_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_8955, mcs1_mcs_mat1_6_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_7551, mcs1_mcs_mat1_6_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_7992, mcs1_mcs_mat1_6_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_8956, mcs1_mcs_mat1_6_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_7130, mcs1_mcs_mat1_6_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_9302, mcs1_mcs_mat1_6_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_8475, mcs1_mcs_mat1_6_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_6609, shiftr_out[100]}), .c ({new_AGEMA_signal_8956, mcs1_mcs_mat1_6_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_6833, mcs1_mcs_mat1_6_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7993, mcs1_mcs_mat1_6_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_8475, mcs1_mcs_mat1_6_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[979]), .c ({new_AGEMA_signal_7993, mcs1_mcs_mat1_6_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[980]), .c ({new_AGEMA_signal_7130, mcs1_mcs_mat1_6_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[981]), .c ({new_AGEMA_signal_7551, mcs1_mcs_mat1_6_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_8957, mcs1_mcs_mat1_6_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_9303, mcs1_mcs_mat1_6_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_8477, mcs1_mcs_mat1_6_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7995, mcs1_mcs_mat1_6_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_8957, mcs1_mcs_mat1_6_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_7269, mcs1_mcs_mat1_6_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_7994, mcs1_mcs_mat1_6_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_7995, mcs1_mcs_mat1_6_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_7269, mcs1_mcs_mat1_6_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_8476, mcs1_mcs_mat1_6_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_7131, mcs1_mcs_mat1_6_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_7132, mcs1_mcs_mat1_6_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_7269, mcs1_mcs_mat1_6_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_7552, mcs1_mcs_mat1_6_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_6614, shiftr_out[68]}), .c ({new_AGEMA_signal_7995, mcs1_mcs_mat1_6_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_8958, mcs1_mcs_mat1_6_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_7131, mcs1_mcs_mat1_6_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_9304, mcs1_mcs_mat1_6_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_8477, mcs1_mcs_mat1_6_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_7552, mcs1_mcs_mat1_6_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_8958, mcs1_mcs_mat1_6_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_7228, shiftr_out[71]}), .b ({new_AGEMA_signal_7996, mcs1_mcs_mat1_6_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_8477, mcs1_mcs_mat1_6_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[982]), .c ({new_AGEMA_signal_7996, mcs1_mcs_mat1_6_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[983]), .c ({new_AGEMA_signal_7132, mcs1_mcs_mat1_6_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7228, shiftr_out[71]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[984]), .c ({new_AGEMA_signal_7552, mcs1_mcs_mat1_6_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_10010, mcs1_mcs_mat1_6_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_9570, mcs1_mcs_mat1_6_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_10231, mcs1_mcs_mat1_6_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_9794, mcs1_mcs_mat1_6_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_10232, mcs1_mcs_mat1_6_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_10470, mcs1_mcs_mat1_6_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_10010, mcs1_mcs_mat1_6_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_10232, mcs1_mcs_mat1_6_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_10471, mcs1_mcs_mat1_6_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_9570, mcs1_mcs_mat1_6_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_10011, mcs1_mcs_mat1_6_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_10232, mcs1_mcs_mat1_6_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({new_AGEMA_signal_8959, mcs1_mcs_mat1_6_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_9570, mcs1_mcs_mat1_6_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_9793, mcs1_mcs_mat1_6_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_9360, shiftr_out[37]}), .c ({new_AGEMA_signal_10010, mcs1_mcs_mat1_6_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_9571, mcs1_mcs_mat1_6_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8478, mcs1_mcs_mat1_6_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_9793, mcs1_mcs_mat1_6_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_10011, mcs1_mcs_mat1_6_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_9794, mcs1_mcs_mat1_6_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_10233, mcs1_mcs_mat1_6_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_9571, mcs1_mcs_mat1_6_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_9794, mcs1_mcs_mat1_6_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({new_AGEMA_signal_9795, mcs1_mcs_mat1_6_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_10011, mcs1_mcs_mat1_6_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9360, shiftr_out[37]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[985]), .c ({new_AGEMA_signal_9795, mcs1_mcs_mat1_6_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[986]), .c ({new_AGEMA_signal_8959, mcs1_mcs_mat1_6_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[987]), .c ({new_AGEMA_signal_9571, mcs1_mcs_mat1_6_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_8961, mcs1_mcs_mat1_6_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_9305, mcs1_mcs_mat1_6_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({new_AGEMA_signal_8479, mcs1_mcs_mat1_6_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_8960, mcs1_mcs_mat1_6_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_9306, mcs1_mcs_mat1_6_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_7553, mcs1_mcs_mat1_6_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_9572, mcs1_mcs_mat1_6_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_8961, mcs1_mcs_mat1_6_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .c ({new_AGEMA_signal_9306, mcs1_mcs_mat1_6_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_7133, mcs1_mcs_mat1_6_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_8479, mcs1_mcs_mat1_6_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_8961, mcs1_mcs_mat1_6_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_6835, mcs1_mcs_mat1_6_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_7998, mcs1_mcs_mat1_6_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_8479, mcs1_mcs_mat1_6_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7307, shiftr_out[5]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[988]), .c ({new_AGEMA_signal_7998, mcs1_mcs_mat1_6_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[989]), .c ({new_AGEMA_signal_7133, mcs1_mcs_mat1_6_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[990]), .c ({new_AGEMA_signal_7553, mcs1_mcs_mat1_6_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_8482, mcs1_mcs_mat1_6_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7554, mcs1_mcs_mat1_6_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_8962, mcs1_mcs_mat1_6_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_7134, mcs1_mcs_mat1_6_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_7999, mcs1_mcs_mat1_6_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8480, mcs1_mcs_mat1_6_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({new_AGEMA_signal_8000, mcs1_mcs_mat1_6_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_8481, mcs1_mcs_mat1_6_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[991]), .c ({new_AGEMA_signal_8000, mcs1_mcs_mat1_6_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[992]), .c ({new_AGEMA_signal_7134, mcs1_mcs_mat1_6_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[993]), .c ({new_AGEMA_signal_7554, mcs1_mcs_mat1_6_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_7136, mcs1_mcs_mat1_6_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_7555, mcs1_mcs_mat1_6_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_8001, mcs1_mcs_mat1_6_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_7137, mcs1_mcs_mat1_6_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_8002, mcs1_mcs_mat1_6_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_8484, mcs1_mcs_mat1_6_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_8485, mcs1_mcs_mat1_6_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_8003, mcs1_mcs_mat1_6_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_8964, mcs1_mcs_mat1_6_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_8004, mcs1_mcs_mat1_6_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_8485, mcs1_mcs_mat1_6_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[994]), .c ({new_AGEMA_signal_8004, mcs1_mcs_mat1_6_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[995]), .c ({new_AGEMA_signal_7137, mcs1_mcs_mat1_6_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7228, shiftr_out[71]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[996]), .c ({new_AGEMA_signal_7555, mcs1_mcs_mat1_6_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_9797, mcs1_mcs_mat1_6_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_10012, mcs1_mcs_mat1_6_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_10234, mcs1_mcs_mat1_6_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_10235, mcs1_mcs_mat1_6_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_9796, mcs1_mcs_mat1_6_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_10472, mcs1_mcs_mat1_6_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_9573, mcs1_mcs_mat1_6_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_9796, mcs1_mcs_mat1_6_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({new_AGEMA_signal_10235, mcs1_mcs_mat1_6_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_10473, mcs1_mcs_mat1_6_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_8486, mcs1_mcs_mat1_6_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_10012, mcs1_mcs_mat1_6_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_10235, mcs1_mcs_mat1_6_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_8965, mcs1_mcs_mat1_6_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_9799, mcs1_mcs_mat1_6_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_10012, mcs1_mcs_mat1_6_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_9798, mcs1_mcs_mat1_6_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_10013, mcs1_mcs_mat1_6_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_10236, mcs1_mcs_mat1_6_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_9797, mcs1_mcs_mat1_6_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8965, mcs1_mcs_mat1_6_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_10013, mcs1_mcs_mat1_6_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_9573, mcs1_mcs_mat1_6_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_9797, mcs1_mcs_mat1_6_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9360, shiftr_out[37]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[997]), .c ({new_AGEMA_signal_9799, mcs1_mcs_mat1_6_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[998]), .c ({new_AGEMA_signal_8965, mcs1_mcs_mat1_6_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[999]), .c ({new_AGEMA_signal_9573, mcs1_mcs_mat1_6_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_7557, mcs1_mcs_mat1_6_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_8006, mcs1_mcs_mat1_6_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_9308, mcs1_mcs_mat1_6_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_7138, mcs1_mcs_mat1_6_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_9574, mcs1_mcs_mat1_6_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_8966, mcs1_mcs_mat1_6_mcs_out[47]}), .b ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_9308, mcs1_mcs_mat1_6_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_8488, mcs1_mcs_mat1_6_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_6609, shiftr_out[100]}), .c ({new_AGEMA_signal_8966, mcs1_mcs_mat1_6_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_6838, mcs1_mcs_mat1_6_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_8007, mcs1_mcs_mat1_6_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_8488, mcs1_mcs_mat1_6_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1000]), .c ({new_AGEMA_signal_8007, mcs1_mcs_mat1_6_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1001]), .c ({new_AGEMA_signal_7138, mcs1_mcs_mat1_6_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1002]), .c ({new_AGEMA_signal_7557, mcs1_mcs_mat1_6_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_8489, mcs1_mcs_mat1_6_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_7558, mcs1_mcs_mat1_6_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_8967, mcs1_mcs_mat1_6_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_8008, mcs1_mcs_mat1_6_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7139, mcs1_mcs_mat1_6_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_8489, mcs1_mcs_mat1_6_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_8490, mcs1_mcs_mat1_6_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_8010, mcs1_mcs_mat1_6_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_8968, mcs1_mcs_mat1_6_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_8491, mcs1_mcs_mat1_6_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_6839, mcs1_mcs_mat1_6_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_8969, mcs1_mcs_mat1_6_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_8008, mcs1_mcs_mat1_6_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7559, mcs1_mcs_mat1_6_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8491, mcs1_mcs_mat1_6_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_8009, mcs1_mcs_mat1_6_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_7559, mcs1_mcs_mat1_6_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_8492, mcs1_mcs_mat1_6_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1003]), .c ({new_AGEMA_signal_8010, mcs1_mcs_mat1_6_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1004]), .c ({new_AGEMA_signal_7139, mcs1_mcs_mat1_6_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7228, shiftr_out[71]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1005]), .c ({new_AGEMA_signal_7559, mcs1_mcs_mat1_6_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_10237, mcs1_mcs_mat1_6_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_8493, mcs1_mcs_mat1_6_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_10474, mcs1_mcs_mat1_6_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_9576, mcs1_mcs_mat1_6_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_9575, mcs1_mcs_mat1_6_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_9800, mcs1_mcs_mat1_6_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({new_AGEMA_signal_10237, mcs1_mcs_mat1_6_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_10475, mcs1_mcs_mat1_6_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_9801, mcs1_mcs_mat1_6_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_10014, mcs1_mcs_mat1_6_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_10237, mcs1_mcs_mat1_6_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_9802, mcs1_mcs_mat1_6_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9577, mcs1_mcs_mat1_6_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_10014, mcs1_mcs_mat1_6_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_9802, mcs1_mcs_mat1_6_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9576, mcs1_mcs_mat1_6_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_10015, mcs1_mcs_mat1_6_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_9309, mcs1_mcs_mat1_6_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_9576, mcs1_mcs_mat1_6_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({new_AGEMA_signal_8970, mcs1_mcs_mat1_6_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_9309, mcs1_mcs_mat1_6_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9360, shiftr_out[37]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1006]), .c ({new_AGEMA_signal_9802, mcs1_mcs_mat1_6_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1007]), .c ({new_AGEMA_signal_8970, mcs1_mcs_mat1_6_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1008]), .c ({new_AGEMA_signal_9577, mcs1_mcs_mat1_6_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_8011, mcs1_mcs_mat1_6_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7560, mcs1_mcs_mat1_6_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_8494, mcs1_mcs_mat1_6_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_7140, mcs1_mcs_mat1_6_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_7270, mcs1_mcs_mat1_6_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_9310, mcs1_mcs_mat1_6_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_8012, mcs1_mcs_mat1_6_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_9578, mcs1_mcs_mat1_6_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7307, shiftr_out[5]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1009]), .c ({new_AGEMA_signal_8012, mcs1_mcs_mat1_6_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1010]), .c ({new_AGEMA_signal_7140, mcs1_mcs_mat1_6_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1011]), .c ({new_AGEMA_signal_7560, mcs1_mcs_mat1_6_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_8972, mcs1_mcs_mat1_6_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_8496, mcs1_mcs_mat1_6_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_9311, mcs1_mcs_mat1_6_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_7142, mcs1_mcs_mat1_6_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_8497, mcs1_mcs_mat1_6_mcs_out[29]}), .c ({new_AGEMA_signal_8972, mcs1_mcs_mat1_6_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_7141, mcs1_mcs_mat1_6_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_8496, mcs1_mcs_mat1_6_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_8973, mcs1_mcs_mat1_6_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_8015, mcs1_mcs_mat1_6_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_6609, shiftr_out[100]}), .c ({new_AGEMA_signal_8496, mcs1_mcs_mat1_6_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_8974, mcs1_mcs_mat1_6_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_8013, mcs1_mcs_mat1_6_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_9312, mcs1_mcs_mat1_6_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_8498, mcs1_mcs_mat1_6_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_8014, mcs1_mcs_mat1_6_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_8974, mcs1_mcs_mat1_6_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_7561, mcs1_mcs_mat1_6_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_8014, mcs1_mcs_mat1_6_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_8015, mcs1_mcs_mat1_6_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7142, mcs1_mcs_mat1_6_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_8498, mcs1_mcs_mat1_6_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1012]), .c ({new_AGEMA_signal_8015, mcs1_mcs_mat1_6_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1013]), .c ({new_AGEMA_signal_7142, mcs1_mcs_mat1_6_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1014]), .c ({new_AGEMA_signal_7561, mcs1_mcs_mat1_6_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_8016, mcs1_mcs_mat1_6_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_8499, mcs1_mcs_mat1_6_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_7562, mcs1_mcs_mat1_6_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7143, mcs1_mcs_mat1_6_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_8016, mcs1_mcs_mat1_6_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_8500, mcs1_mcs_mat1_6_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_8975, mcs1_mcs_mat1_6_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_8018, mcs1_mcs_mat1_6_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_7143, mcs1_mcs_mat1_6_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_8500, mcs1_mcs_mat1_6_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_8976, mcs1_mcs_mat1_6_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_6614, shiftr_out[68]}), .c ({new_AGEMA_signal_9313, mcs1_mcs_mat1_6_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_8018, mcs1_mcs_mat1_6_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8501, mcs1_mcs_mat1_6_mcs_out[24]}), .c ({new_AGEMA_signal_8976, mcs1_mcs_mat1_6_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_8017, mcs1_mcs_mat1_6_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_7228, shiftr_out[71]}), .c ({new_AGEMA_signal_8501, mcs1_mcs_mat1_6_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_7562, mcs1_mcs_mat1_6_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_6842, mcs1_mcs_mat1_6_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_8017, mcs1_mcs_mat1_6_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1015]), .c ({new_AGEMA_signal_8018, mcs1_mcs_mat1_6_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1016]), .c ({new_AGEMA_signal_7143, mcs1_mcs_mat1_6_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7228, shiftr_out[71]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1017]), .c ({new_AGEMA_signal_7562, mcs1_mcs_mat1_6_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_9803, mcs1_mcs_mat1_6_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_8098, shiftr_out[38]}), .c ({new_AGEMA_signal_10016, mcs1_mcs_mat1_6_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_9579, mcs1_mcs_mat1_6_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8977, mcs1_mcs_mat1_6_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_9803, mcs1_mcs_mat1_6_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_10017, mcs1_mcs_mat1_6_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_9360, shiftr_out[37]}), .c ({new_AGEMA_signal_10238, mcs1_mcs_mat1_6_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_9805, mcs1_mcs_mat1_6_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8977, mcs1_mcs_mat1_6_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_10017, mcs1_mcs_mat1_6_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_10239, mcs1_mcs_mat1_6_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_7618, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_10476, mcs1_mcs_mat1_6_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_9805, mcs1_mcs_mat1_6_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_10018, mcs1_mcs_mat1_6_mcs_out[20]}), .c ({new_AGEMA_signal_10239, mcs1_mcs_mat1_6_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_9804, mcs1_mcs_mat1_6_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_10018, mcs1_mcs_mat1_6_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_9579, mcs1_mcs_mat1_6_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8502, mcs1_mcs_mat1_6_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_9804, mcs1_mcs_mat1_6_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9360, shiftr_out[37]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1018]), .c ({new_AGEMA_signal_9805, mcs1_mcs_mat1_6_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1019]), .c ({new_AGEMA_signal_8977, mcs1_mcs_mat1_6_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1020]), .c ({new_AGEMA_signal_9579, mcs1_mcs_mat1_6_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_8019, mcs1_mcs_mat1_6_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_8022, mcs1_mcs_mat1_6_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_8503, mcs1_mcs_mat1_6_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_8504, mcs1_mcs_mat1_6_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_6843, mcs1_mcs_mat1_6_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_8978, mcs1_mcs_mat1_6_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_8979, mcs1_mcs_mat1_6_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_7144, mcs1_mcs_mat1_6_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_9314, mcs1_mcs_mat1_6_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_6627, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_8504, mcs1_mcs_mat1_6_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_8979, mcs1_mcs_mat1_6_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_8020, mcs1_mcs_mat1_6_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_7307, shiftr_out[5]}), .c ({new_AGEMA_signal_8504, mcs1_mcs_mat1_6_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_7563, mcs1_mcs_mat1_6_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_7564, mcs1_mcs_mat1_6_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_8020, mcs1_mcs_mat1_6_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_8021, mcs1_mcs_mat1_6_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_7144, mcs1_mcs_mat1_6_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_8505, mcs1_mcs_mat1_6_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7307, shiftr_out[5]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1021]), .c ({new_AGEMA_signal_8022, mcs1_mcs_mat1_6_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1022]), .c ({new_AGEMA_signal_7144, mcs1_mcs_mat1_6_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1023]), .c ({new_AGEMA_signal_7564, mcs1_mcs_mat1_6_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_8982, mcs1_mcs_mat1_6_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_7271, mcs1_mcs_mat1_6_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_9315, mcs1_mcs_mat1_6_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_8508, mcs1_mcs_mat1_6_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_8506, mcs1_mcs_mat1_6_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_8980, mcs1_mcs_mat1_6_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_8024, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_7145, mcs1_mcs_mat1_6_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8506, mcs1_mcs_mat1_6_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_7271, mcs1_mcs_mat1_6_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_8507, mcs1_mcs_mat1_6_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_8981, mcs1_mcs_mat1_6_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_8023, mcs1_mcs_mat1_6_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_8024, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_8507, mcs1_mcs_mat1_6_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_6844, mcs1_mcs_mat1_6_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_7145, mcs1_mcs_mat1_6_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_7271, mcs1_mcs_mat1_6_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_9316, mcs1_mcs_mat1_6_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_9580, mcs1_mcs_mat1_6_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_8982, mcs1_mcs_mat1_6_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_8024, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_9316, mcs1_mcs_mat1_6_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_8508, mcs1_mcs_mat1_6_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_8982, mcs1_mcs_mat1_6_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_8023, mcs1_mcs_mat1_6_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_8508, mcs1_mcs_mat1_6_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_6609, shiftr_out[100]}), .b ({new_AGEMA_signal_7565, mcs1_mcs_mat1_6_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_8023, mcs1_mcs_mat1_6_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7289, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1024]), .c ({new_AGEMA_signal_8024, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6677, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1025]), .c ({new_AGEMA_signal_7145, mcs1_mcs_mat1_6_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7223, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1026]), .c ({new_AGEMA_signal_7565, mcs1_mcs_mat1_6_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_7272, mcs1_mcs_mat1_6_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_7228, shiftr_out[71]}), .c ({new_AGEMA_signal_7566, mcs1_mcs_mat1_6_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_8510, mcs1_mcs_mat1_6_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_8983, mcs1_mcs_mat1_6_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_8025, mcs1_mcs_mat1_6_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_8509, mcs1_mcs_mat1_6_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_7567, mcs1_mcs_mat1_6_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_7272, mcs1_mcs_mat1_6_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_8025, mcs1_mcs_mat1_6_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_6845, mcs1_mcs_mat1_6_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_7146, mcs1_mcs_mat1_6_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_7272, mcs1_mcs_mat1_6_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_8984, mcs1_mcs_mat1_6_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_6614, shiftr_out[68]}), .c ({new_AGEMA_signal_9317, mcs1_mcs_mat1_6_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_6845, mcs1_mcs_mat1_6_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8510, mcs1_mcs_mat1_6_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_8984, mcs1_mcs_mat1_6_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_8026, mcs1_mcs_mat1_6_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_7567, mcs1_mcs_mat1_6_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_8510, mcs1_mcs_mat1_6_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7294, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1027]), .c ({new_AGEMA_signal_8026, mcs1_mcs_mat1_6_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6682, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1028]), .c ({new_AGEMA_signal_7146, mcs1_mcs_mat1_6_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7228, shiftr_out[71]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1029]), .c ({new_AGEMA_signal_7567, mcs1_mcs_mat1_6_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_10728, mcs1_mcs_mat1_6_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_9582, mcs1_mcs_mat1_6_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_10930, mcs1_mcs_mat1_6_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_10477, mcs1_mcs_mat1_6_mcs_out[7]}), .b ({new_AGEMA_signal_8098, shiftr_out[38]}), .c ({new_AGEMA_signal_10728, mcs1_mcs_mat1_6_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_10240, mcs1_mcs_mat1_6_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_9360, shiftr_out[37]}), .c ({new_AGEMA_signal_10477, mcs1_mcs_mat1_6_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_10019, mcs1_mcs_mat1_6_mcs_out[6]}), .b ({new_AGEMA_signal_8986, mcs1_mcs_mat1_6_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_10240, mcs1_mcs_mat1_6_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_8985, mcs1_mcs_mat1_6_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_9806, mcs1_mcs_mat1_6_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_10019, mcs1_mcs_mat1_6_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9360, shiftr_out[37]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1030]), .c ({new_AGEMA_signal_9806, mcs1_mcs_mat1_6_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8098, shiftr_out[38]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1031]), .c ({new_AGEMA_signal_8986, mcs1_mcs_mat1_6_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1032]), .c ({new_AGEMA_signal_9582, mcs1_mcs_mat1_6_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_7568, mcs1_mcs_mat1_6_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_8027, mcs1_mcs_mat1_6_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_8513, mcs1_mcs_mat1_6_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_7307, shiftr_out[5]}), .b ({new_AGEMA_signal_7569, mcs1_mcs_mat1_6_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_8027, mcs1_mcs_mat1_6_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_8514, mcs1_mcs_mat1_6_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_7147, mcs1_mcs_mat1_6_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_8987, mcs1_mcs_mat1_6_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_8515, mcs1_mcs_mat1_6_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_8029, mcs1_mcs_mat1_6_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_8988, mcs1_mcs_mat1_6_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_8030, mcs1_mcs_mat1_6_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_6846, mcs1_mcs_mat1_6_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8515, mcs1_mcs_mat1_6_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7307, shiftr_out[5]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1033]), .c ({new_AGEMA_signal_8030, mcs1_mcs_mat1_6_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6695, shiftr_out[6]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1034]), .c ({new_AGEMA_signal_7147, mcs1_mcs_mat1_6_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7241, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1035]), .c ({new_AGEMA_signal_7569, mcs1_mcs_mat1_6_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U96 ( .a ({new_AGEMA_signal_9583, mcs1_mcs_mat1_7_n128}), .b ({new_AGEMA_signal_10478, mcs1_mcs_mat1_7_n127}), .c ({temp_next_s1[65], temp_next_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U95 ( .a ({new_AGEMA_signal_10263, mcs1_mcs_mat1_7_mcs_out[41]}), .b ({new_AGEMA_signal_8066, mcs1_mcs_mat1_7_mcs_out[45]}), .c ({new_AGEMA_signal_10478, mcs1_mcs_mat1_7_n127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U94 ( .a ({new_AGEMA_signal_7274, mcs1_mcs_mat1_7_mcs_out[33]}), .b ({new_AGEMA_signal_9344, mcs1_mcs_mat1_7_mcs_out[37]}), .c ({new_AGEMA_signal_9583, mcs1_mcs_mat1_7_n128}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U93 ( .a ({new_AGEMA_signal_9807, mcs1_mcs_mat1_7_n126}), .b ({new_AGEMA_signal_10241, mcs1_mcs_mat1_7_n125}), .c ({temp_next_s1[64], temp_next_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U92 ( .a ({new_AGEMA_signal_10040, mcs1_mcs_mat1_7_mcs_out[40]}), .b ({new_AGEMA_signal_9609, mcs1_mcs_mat1_7_mcs_out[44]}), .c ({new_AGEMA_signal_10241, mcs1_mcs_mat1_7_n125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U91 ( .a ({new_AGEMA_signal_9612, mcs1_mcs_mat1_7_mcs_out[32]}), .b ({new_AGEMA_signal_8550, mcs1_mcs_mat1_7_mcs_out[36]}), .c ({new_AGEMA_signal_9807, mcs1_mcs_mat1_7_n126}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U90 ( .a ({new_AGEMA_signal_8989, mcs1_mcs_mat1_7_n124}), .b ({new_AGEMA_signal_10242, mcs1_mcs_mat1_7_n123}), .c ({temp_next_s1[35], temp_next_s0[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U89 ( .a ({new_AGEMA_signal_10041, mcs1_mcs_mat1_7_mcs_out[27]}), .b ({new_AGEMA_signal_9346, mcs1_mcs_mat1_7_mcs_out[31]}), .c ({new_AGEMA_signal_10242, mcs1_mcs_mat1_7_n123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U88 ( .a ({new_AGEMA_signal_8560, mcs1_mcs_mat1_7_mcs_out[19]}), .b ({new_AGEMA_signal_8557, mcs1_mcs_mat1_7_mcs_out[23]}), .c ({new_AGEMA_signal_8989, mcs1_mcs_mat1_7_n124}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U87 ( .a ({new_AGEMA_signal_9318, mcs1_mcs_mat1_7_n122}), .b ({new_AGEMA_signal_10481, mcs1_mcs_mat1_7_n121}), .c ({temp_next_s1[34], temp_next_s0[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U86 ( .a ({new_AGEMA_signal_10264, mcs1_mcs_mat1_7_mcs_out[26]}), .b ({new_AGEMA_signal_9034, mcs1_mcs_mat1_7_mcs_out[30]}), .c ({new_AGEMA_signal_10481, mcs1_mcs_mat1_7_n121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U85 ( .a ({new_AGEMA_signal_9039, mcs1_mcs_mat1_7_mcs_out[18]}), .b ({new_AGEMA_signal_9037, mcs1_mcs_mat1_7_mcs_out[22]}), .c ({new_AGEMA_signal_9318, mcs1_mcs_mat1_7_n122}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U84 ( .a ({new_AGEMA_signal_9584, mcs1_mcs_mat1_7_n120}), .b ({new_AGEMA_signal_10731, mcs1_mcs_mat1_7_n119}), .c ({temp_next_s1[33], temp_next_s0[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U83 ( .a ({new_AGEMA_signal_10500, mcs1_mcs_mat1_7_mcs_out[25]}), .b ({new_AGEMA_signal_8554, mcs1_mcs_mat1_7_mcs_out[29]}), .c ({new_AGEMA_signal_10731, mcs1_mcs_mat1_7_n119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U82 ( .a ({new_AGEMA_signal_9349, mcs1_mcs_mat1_7_mcs_out[17]}), .b ({new_AGEMA_signal_9348, mcs1_mcs_mat1_7_mcs_out[21]}), .c ({new_AGEMA_signal_9584, mcs1_mcs_mat1_7_n120}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U81 ( .a ({new_AGEMA_signal_8990, mcs1_mcs_mat1_7_n118}), .b ({new_AGEMA_signal_10243, mcs1_mcs_mat1_7_n117}), .c ({temp_next_s1[32], temp_next_s0[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U80 ( .a ({new_AGEMA_signal_10043, mcs1_mcs_mat1_7_mcs_out[24]}), .b ({new_AGEMA_signal_9347, mcs1_mcs_mat1_7_mcs_out[28]}), .c ({new_AGEMA_signal_10243, mcs1_mcs_mat1_7_n117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U79 ( .a ({new_AGEMA_signal_8562, mcs1_mcs_mat1_7_mcs_out[16]}), .b ({new_AGEMA_signal_8559, mcs1_mcs_mat1_7_mcs_out[20]}), .c ({new_AGEMA_signal_8990, mcs1_mcs_mat1_7_n118}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U78 ( .a ({new_AGEMA_signal_9808, mcs1_mcs_mat1_7_n116}), .b ({new_AGEMA_signal_9585, mcs1_mcs_mat1_7_n115}), .c ({temp_next_s1[3], temp_next_s0[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U77 ( .a ({new_AGEMA_signal_8568, mcs1_mcs_mat1_7_mcs_out[3]}), .b ({new_AGEMA_signal_9353, mcs1_mcs_mat1_7_mcs_out[7]}), .c ({new_AGEMA_signal_9585, mcs1_mcs_mat1_7_n115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U76 ( .a ({new_AGEMA_signal_9615, mcs1_mcs_mat1_7_mcs_out[11]}), .b ({new_AGEMA_signal_9350, mcs1_mcs_mat1_7_mcs_out[15]}), .c ({new_AGEMA_signal_9808, mcs1_mcs_mat1_7_n116}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U75 ( .a ({new_AGEMA_signal_9586, mcs1_mcs_mat1_7_n114}), .b ({new_AGEMA_signal_10732, mcs1_mcs_mat1_7_n113}), .c ({new_AGEMA_signal_10932, mcs_out[227]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U74 ( .a ({new_AGEMA_signal_10495, mcs1_mcs_mat1_7_mcs_out[123]}), .b ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_10732, mcs1_mcs_mat1_7_n113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U73 ( .a ({new_AGEMA_signal_9001, mcs1_mcs_mat1_7_mcs_out[115]}), .b ({new_AGEMA_signal_9324, mcs1_mcs_mat1_7_mcs_out[119]}), .c ({new_AGEMA_signal_9586, mcs1_mcs_mat1_7_n114}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U72 ( .a ({new_AGEMA_signal_9587, mcs1_mcs_mat1_7_n112}), .b ({new_AGEMA_signal_10021, mcs1_mcs_mat1_7_n111}), .c ({new_AGEMA_signal_10244, mcs_out[226]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U71 ( .a ({new_AGEMA_signal_9815, mcs1_mcs_mat1_7_mcs_out[122]}), .b ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_10021, mcs1_mcs_mat1_7_n111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U70 ( .a ({new_AGEMA_signal_8519, mcs1_mcs_mat1_7_mcs_out[114]}), .b ({new_AGEMA_signal_9325, mcs1_mcs_mat1_7_mcs_out[118]}), .c ({new_AGEMA_signal_9587, mcs1_mcs_mat1_7_n112}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U69 ( .a ({new_AGEMA_signal_10483, mcs1_mcs_mat1_7_n110}), .b ({new_AGEMA_signal_8991, mcs1_mcs_mat1_7_n109}), .c ({temp_next_s1[2], temp_next_s0[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U68 ( .a ({new_AGEMA_signal_8569, mcs1_mcs_mat1_7_mcs_out[2]}), .b ({new_AGEMA_signal_8567, mcs1_mcs_mat1_7_mcs_out[6]}), .c ({new_AGEMA_signal_8991, mcs1_mcs_mat1_7_n109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U67 ( .a ({new_AGEMA_signal_10266, mcs1_mcs_mat1_7_mcs_out[10]}), .b ({new_AGEMA_signal_9041, mcs1_mcs_mat1_7_mcs_out[14]}), .c ({new_AGEMA_signal_10483, mcs1_mcs_mat1_7_n110}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U66 ( .a ({new_AGEMA_signal_9319, mcs1_mcs_mat1_7_n108}), .b ({new_AGEMA_signal_10734, mcs1_mcs_mat1_7_n107}), .c ({new_AGEMA_signal_10933, mcs_out[225]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U65 ( .a ({new_AGEMA_signal_10496, mcs1_mcs_mat1_7_mcs_out[121]}), .b ({new_AGEMA_signal_7570, mcs1_mcs_mat1_7_mcs_out[125]}), .c ({new_AGEMA_signal_10734, mcs1_mcs_mat1_7_n107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U64 ( .a ({new_AGEMA_signal_8034, mcs1_mcs_mat1_7_mcs_out[113]}), .b ({new_AGEMA_signal_9000, mcs1_mcs_mat1_7_mcs_out[117]}), .c ({new_AGEMA_signal_9319, mcs1_mcs_mat1_7_n108}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U63 ( .a ({new_AGEMA_signal_9588, mcs1_mcs_mat1_7_n106}), .b ({new_AGEMA_signal_10484, mcs1_mcs_mat1_7_n105}), .c ({new_AGEMA_signal_10735, mcs_out[224]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U62 ( .a ({new_AGEMA_signal_10253, mcs1_mcs_mat1_7_mcs_out[120]}), .b ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_10484, mcs1_mcs_mat1_7_n105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U61 ( .a ({new_AGEMA_signal_9326, mcs1_mcs_mat1_7_mcs_out[112]}), .b ({new_AGEMA_signal_8518, mcs1_mcs_mat1_7_mcs_out[116]}), .c ({new_AGEMA_signal_9588, mcs1_mcs_mat1_7_n106}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U60 ( .a ({new_AGEMA_signal_10485, mcs1_mcs_mat1_7_n104}), .b ({new_AGEMA_signal_9589, mcs1_mcs_mat1_7_n103}), .c ({new_AGEMA_signal_10736, mcs_out[195]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U59 ( .a ({new_AGEMA_signal_9327, mcs1_mcs_mat1_7_mcs_out[111]}), .b ({new_AGEMA_signal_9331, mcs1_mcs_mat1_7_mcs_out[99]}), .c ({new_AGEMA_signal_9589, mcs1_mcs_mat1_7_n103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U58 ( .a ({new_AGEMA_signal_9006, mcs1_mcs_mat1_7_mcs_out[103]}), .b ({new_AGEMA_signal_10254, mcs1_mcs_mat1_7_mcs_out[107]}), .c ({new_AGEMA_signal_10485, mcs1_mcs_mat1_7_n104}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U57 ( .a ({new_AGEMA_signal_10486, mcs1_mcs_mat1_7_n102}), .b ({new_AGEMA_signal_9590, mcs1_mcs_mat1_7_n101}), .c ({new_AGEMA_signal_10737, mcs_out[194]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U56 ( .a ({new_AGEMA_signal_9328, mcs1_mcs_mat1_7_mcs_out[110]}), .b ({new_AGEMA_signal_8528, mcs1_mcs_mat1_7_mcs_out[98]}), .c ({new_AGEMA_signal_9590, mcs1_mcs_mat1_7_n101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U55 ( .a ({new_AGEMA_signal_8039, mcs1_mcs_mat1_7_mcs_out[102]}), .b ({new_AGEMA_signal_10255, mcs1_mcs_mat1_7_mcs_out[106]}), .c ({new_AGEMA_signal_10486, mcs1_mcs_mat1_7_n102}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U54 ( .a ({new_AGEMA_signal_10487, mcs1_mcs_mat1_7_n100}), .b ({new_AGEMA_signal_9591, mcs1_mcs_mat1_7_n99}), .c ({new_AGEMA_signal_10738, mcs_out[193]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U53 ( .a ({new_AGEMA_signal_9329, mcs1_mcs_mat1_7_mcs_out[109]}), .b ({new_AGEMA_signal_7579, mcs1_mcs_mat1_7_mcs_out[97]}), .c ({new_AGEMA_signal_9591, mcs1_mcs_mat1_7_n99}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U52 ( .a ({new_AGEMA_signal_8526, mcs1_mcs_mat1_7_mcs_out[101]}), .b ({new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[105]}), .c ({new_AGEMA_signal_10487, mcs1_mcs_mat1_7_n100}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U51 ( .a ({new_AGEMA_signal_10739, mcs1_mcs_mat1_7_n98}), .b ({new_AGEMA_signal_10022, mcs1_mcs_mat1_7_n97}), .c ({new_AGEMA_signal_10934, mcs_out[192]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U50 ( .a ({new_AGEMA_signal_9330, mcs1_mcs_mat1_7_mcs_out[108]}), .b ({new_AGEMA_signal_9819, mcs1_mcs_mat1_7_mcs_out[96]}), .c ({new_AGEMA_signal_10022, mcs1_mcs_mat1_7_n97}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U49 ( .a ({new_AGEMA_signal_9007, mcs1_mcs_mat1_7_mcs_out[100]}), .b ({new_AGEMA_signal_10497, mcs1_mcs_mat1_7_mcs_out[104]}), .c ({new_AGEMA_signal_10739, mcs1_mcs_mat1_7_n98}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U48 ( .a ({new_AGEMA_signal_8992, mcs1_mcs_mat1_7_n96}), .b ({new_AGEMA_signal_9809, mcs1_mcs_mat1_7_n95}), .c ({new_AGEMA_signal_10023, mcs_out[163]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U47 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_9009, mcs1_mcs_mat1_7_mcs_out[95]}), .c ({new_AGEMA_signal_9809, mcs1_mcs_mat1_7_n95}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U46 ( .a ({new_AGEMA_signal_8531, mcs1_mcs_mat1_7_mcs_out[83]}), .b ({new_AGEMA_signal_8047, mcs1_mcs_mat1_7_mcs_out[87]}), .c ({new_AGEMA_signal_8992, mcs1_mcs_mat1_7_n96}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U45 ( .a ({new_AGEMA_signal_8993, mcs1_mcs_mat1_7_n94}), .b ({new_AGEMA_signal_9810, mcs1_mcs_mat1_7_n93}), .c ({new_AGEMA_signal_10024, mcs_out[162]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U43 ( .a ({new_AGEMA_signal_8532, mcs1_mcs_mat1_7_mcs_out[82]}), .b ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_8993, mcs1_mcs_mat1_7_n94}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U42 ( .a ({new_AGEMA_signal_8994, mcs1_mcs_mat1_7_n92}), .b ({new_AGEMA_signal_9811, mcs1_mcs_mat1_7_n91}), .c ({new_AGEMA_signal_10025, mcs_out[161]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U41 ( .a ({new_AGEMA_signal_9605, mcs1_mcs_mat1_7_mcs_out[89]}), .b ({new_AGEMA_signal_8045, mcs1_mcs_mat1_7_mcs_out[93]}), .c ({new_AGEMA_signal_9811, mcs1_mcs_mat1_7_n91}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U40 ( .a ({new_AGEMA_signal_8533, mcs1_mcs_mat1_7_mcs_out[81]}), .b ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_8994, mcs1_mcs_mat1_7_n92}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U39 ( .a ({new_AGEMA_signal_9320, mcs1_mcs_mat1_7_n90}), .b ({new_AGEMA_signal_9592, mcs1_mcs_mat1_7_n89}), .c ({new_AGEMA_signal_9812, mcs_out[160]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U38 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_9332, mcs1_mcs_mat1_7_mcs_out[92]}), .c ({new_AGEMA_signal_9592, mcs1_mcs_mat1_7_n89}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U37 ( .a ({new_AGEMA_signal_9011, mcs1_mcs_mat1_7_mcs_out[80]}), .b ({new_AGEMA_signal_8530, mcs1_mcs_mat1_7_mcs_out[84]}), .c ({new_AGEMA_signal_9320, mcs1_mcs_mat1_7_n90}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U36 ( .a ({new_AGEMA_signal_9321, mcs1_mcs_mat1_7_n88}), .b ({new_AGEMA_signal_10245, mcs1_mcs_mat1_7_n87}), .c ({temp_next_s1[1], temp_next_s0[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U35 ( .a ({new_AGEMA_signal_7602, mcs1_mcs_mat1_7_mcs_out[5]}), .b ({new_AGEMA_signal_10044, mcs1_mcs_mat1_7_mcs_out[9]}), .c ({new_AGEMA_signal_10245, mcs1_mcs_mat1_7_n87}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U34 ( .a ({new_AGEMA_signal_9042, mcs1_mcs_mat1_7_mcs_out[13]}), .b ({new_AGEMA_signal_9046, mcs1_mcs_mat1_7_mcs_out[1]}), .c ({new_AGEMA_signal_9321, mcs1_mcs_mat1_7_n88}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U33 ( .a ({new_AGEMA_signal_9593, mcs1_mcs_mat1_7_n86}), .b ({new_AGEMA_signal_10026, mcs1_mcs_mat1_7_n85}), .c ({new_AGEMA_signal_10246, mcs_out[131]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U32 ( .a ({new_AGEMA_signal_9820, mcs1_mcs_mat1_7_mcs_out[75]}), .b ({new_AGEMA_signal_9012, mcs1_mcs_mat1_7_mcs_out[79]}), .c ({new_AGEMA_signal_10026, mcs1_mcs_mat1_7_n85}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U31 ( .a ({new_AGEMA_signal_9337, mcs1_mcs_mat1_7_mcs_out[67]}), .b ({new_AGEMA_signal_9016, mcs1_mcs_mat1_7_mcs_out[71]}), .c ({new_AGEMA_signal_9593, mcs1_mcs_mat1_7_n86}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U30 ( .a ({new_AGEMA_signal_9594, mcs1_mcs_mat1_7_n84}), .b ({new_AGEMA_signal_10740, mcs1_mcs_mat1_7_n83}), .c ({new_AGEMA_signal_10935, mcs_out[130]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U29 ( .a ({new_AGEMA_signal_10498, mcs1_mcs_mat1_7_mcs_out[74]}), .b ({new_AGEMA_signal_7157, mcs1_mcs_mat1_7_mcs_out[78]}), .c ({new_AGEMA_signal_10740, mcs1_mcs_mat1_7_n83}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U28 ( .a ({new_AGEMA_signal_9019, mcs1_mcs_mat1_7_mcs_out[66]}), .b ({new_AGEMA_signal_9335, mcs1_mcs_mat1_7_mcs_out[70]}), .c ({new_AGEMA_signal_9594, mcs1_mcs_mat1_7_n84}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U27 ( .a ({new_AGEMA_signal_9595, mcs1_mcs_mat1_7_n82}), .b ({new_AGEMA_signal_10247, mcs1_mcs_mat1_7_n81}), .c ({new_AGEMA_signal_10489, mcs_out[129]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U26 ( .a ({new_AGEMA_signal_10032, mcs1_mcs_mat1_7_mcs_out[73]}), .b ({new_AGEMA_signal_8052, mcs1_mcs_mat1_7_mcs_out[77]}), .c ({new_AGEMA_signal_10247, mcs1_mcs_mat1_7_n81}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U25 ( .a ({new_AGEMA_signal_8057, mcs1_mcs_mat1_7_mcs_out[65]}), .b ({new_AGEMA_signal_9336, mcs1_mcs_mat1_7_mcs_out[69]}), .c ({new_AGEMA_signal_9595, mcs1_mcs_mat1_7_n82}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U24 ( .a ({new_AGEMA_signal_9813, mcs1_mcs_mat1_7_n80}), .b ({new_AGEMA_signal_10741, mcs1_mcs_mat1_7_n79}), .c ({new_AGEMA_signal_10936, mcs_out[128]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U23 ( .a ({new_AGEMA_signal_10499, mcs1_mcs_mat1_7_mcs_out[72]}), .b ({new_AGEMA_signal_9333, mcs1_mcs_mat1_7_mcs_out[76]}), .c ({new_AGEMA_signal_10741, mcs1_mcs_mat1_7_n79}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U22 ( .a ({new_AGEMA_signal_9607, mcs1_mcs_mat1_7_mcs_out[64]}), .b ({new_AGEMA_signal_9018, mcs1_mcs_mat1_7_mcs_out[68]}), .c ({new_AGEMA_signal_9813, mcs1_mcs_mat1_7_n80}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U21 ( .a ({new_AGEMA_signal_9322, mcs1_mcs_mat1_7_n78}), .b ({new_AGEMA_signal_10248, mcs1_mcs_mat1_7_n77}), .c ({temp_next_s1[99], temp_next_s0[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U20 ( .a ({new_AGEMA_signal_10034, mcs1_mcs_mat1_7_mcs_out[59]}), .b ({new_AGEMA_signal_9021, mcs1_mcs_mat1_7_mcs_out[63]}), .c ({new_AGEMA_signal_10248, mcs1_mcs_mat1_7_n77}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U19 ( .a ({new_AGEMA_signal_8065, mcs1_mcs_mat1_7_mcs_out[51]}), .b ({new_AGEMA_signal_9026, mcs1_mcs_mat1_7_mcs_out[55]}), .c ({new_AGEMA_signal_9322, mcs1_mcs_mat1_7_n78}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U18 ( .a ({new_AGEMA_signal_9596, mcs1_mcs_mat1_7_n76}), .b ({new_AGEMA_signal_10027, mcs1_mcs_mat1_7_n75}), .c ({temp_next_s1[98], temp_next_s0[98]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U17 ( .a ({new_AGEMA_signal_9823, mcs1_mcs_mat1_7_mcs_out[58]}), .b ({new_AGEMA_signal_8540, mcs1_mcs_mat1_7_mcs_out[62]}), .c ({new_AGEMA_signal_10027, mcs1_mcs_mat1_7_n75}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U16 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_9340, mcs1_mcs_mat1_7_mcs_out[54]}), .c ({new_AGEMA_signal_9596, mcs1_mcs_mat1_7_n76}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U15 ( .a ({new_AGEMA_signal_9597, mcs1_mcs_mat1_7_n74}), .b ({new_AGEMA_signal_10250, mcs1_mcs_mat1_7_n73}), .c ({temp_next_s1[97], temp_next_s0[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U14 ( .a ({new_AGEMA_signal_10035, mcs1_mcs_mat1_7_mcs_out[57]}), .b ({new_AGEMA_signal_8541, mcs1_mcs_mat1_7_mcs_out[61]}), .c ({new_AGEMA_signal_10250, mcs1_mcs_mat1_7_n73}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U13 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_9341, mcs1_mcs_mat1_7_mcs_out[53]}), .c ({new_AGEMA_signal_9597, mcs1_mcs_mat1_7_n74}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U12 ( .a ({new_AGEMA_signal_9323, mcs1_mcs_mat1_7_n72}), .b ({new_AGEMA_signal_10492, mcs1_mcs_mat1_7_n71}), .c ({temp_next_s1[96], temp_next_s0[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U11 ( .a ({new_AGEMA_signal_10260, mcs1_mcs_mat1_7_mcs_out[56]}), .b ({new_AGEMA_signal_9339, mcs1_mcs_mat1_7_mcs_out[60]}), .c ({new_AGEMA_signal_10492, mcs1_mcs_mat1_7_n71}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U10 ( .a ({new_AGEMA_signal_8546, mcs1_mcs_mat1_7_mcs_out[48]}), .b ({new_AGEMA_signal_9028, mcs1_mcs_mat1_7_mcs_out[52]}), .c ({new_AGEMA_signal_9323, mcs1_mcs_mat1_7_n72}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U9 ( .a ({new_AGEMA_signal_9598, mcs1_mcs_mat1_7_n70}), .b ({new_AGEMA_signal_10493, mcs1_mcs_mat1_7_n69}), .c ({temp_next_s1[67], temp_next_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U8 ( .a ({new_AGEMA_signal_10261, mcs1_mcs_mat1_7_mcs_out[43]}), .b ({new_AGEMA_signal_9029, mcs1_mcs_mat1_7_mcs_out[47]}), .c ({new_AGEMA_signal_10493, mcs1_mcs_mat1_7_n69}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U7 ( .a ({new_AGEMA_signal_9032, mcs1_mcs_mat1_7_mcs_out[35]}), .b ({new_AGEMA_signal_9343, mcs1_mcs_mat1_7_mcs_out[39]}), .c ({new_AGEMA_signal_9598, mcs1_mcs_mat1_7_n70}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U6 ( .a ({new_AGEMA_signal_8995, mcs1_mcs_mat1_7_n68}), .b ({new_AGEMA_signal_10494, mcs1_mcs_mat1_7_n67}), .c ({temp_next_s1[66], temp_next_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U5 ( .a ({new_AGEMA_signal_10262, mcs1_mcs_mat1_7_mcs_out[42]}), .b ({new_AGEMA_signal_7591, mcs1_mcs_mat1_7_mcs_out[46]}), .c ({new_AGEMA_signal_10494, mcs1_mcs_mat1_7_n67}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U4 ( .a ({new_AGEMA_signal_8551, mcs1_mcs_mat1_7_mcs_out[34]}), .b ({new_AGEMA_signal_8068, mcs1_mcs_mat1_7_mcs_out[38]}), .c ({new_AGEMA_signal_8995, mcs1_mcs_mat1_7_n68}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U3 ( .a ({new_AGEMA_signal_9814, mcs1_mcs_mat1_7_n66}), .b ({new_AGEMA_signal_10745, mcs1_mcs_mat1_7_n65}), .c ({temp_next_s1[0], temp_next_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U2 ( .a ({new_AGEMA_signal_9835, mcs1_mcs_mat1_7_mcs_out[4]}), .b ({new_AGEMA_signal_10501, mcs1_mcs_mat1_7_mcs_out[8]}), .c ({new_AGEMA_signal_10745, mcs1_mcs_mat1_7_n65}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_U1 ( .a ({new_AGEMA_signal_9047, mcs1_mcs_mat1_7_mcs_out[0]}), .b ({new_AGEMA_signal_9614, mcs1_mcs_mat1_7_mcs_out[12]}), .c ({new_AGEMA_signal_9814, mcs1_mcs_mat1_7_n66}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_10251, mcs1_mcs_mat1_7_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_10495, mcs1_mcs_mat1_7_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_10028, mcs1_mcs_mat1_7_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_8516, mcs1_mcs_mat1_7_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_10251, mcs1_mcs_mat1_7_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_8996, mcs1_mcs_mat1_7_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_9599, mcs1_mcs_mat1_7_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_9815, mcs1_mcs_mat1_7_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_8997, mcs1_mcs_mat1_7_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_9054, shiftr_out[67]}), .c ({new_AGEMA_signal_9599, mcs1_mcs_mat1_7_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_10252, mcs1_mcs_mat1_7_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_9054, shiftr_out[67]}), .c ({new_AGEMA_signal_10496, mcs1_mcs_mat1_7_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_10028, mcs1_mcs_mat1_7_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_10252, mcs1_mcs_mat1_7_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_9816, mcs1_mcs_mat1_7_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9600, mcs1_mcs_mat1_7_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_10028, mcs1_mcs_mat1_7_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_10029, mcs1_mcs_mat1_7_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_10253, mcs1_mcs_mat1_7_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_9816, mcs1_mcs_mat1_7_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_8997, mcs1_mcs_mat1_7_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_10029, mcs1_mcs_mat1_7_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1036]), .c ({new_AGEMA_signal_9816, mcs1_mcs_mat1_7_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1037]), .c ({new_AGEMA_signal_8997, mcs1_mcs_mat1_7_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9054, shiftr_out[67]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1038]), .c ({new_AGEMA_signal_9600, mcs1_mcs_mat1_7_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_8998, mcs1_mcs_mat1_7_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_6688, shiftr_out[34]}), .c ({new_AGEMA_signal_9324, mcs1_mcs_mat1_7_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_8517, mcs1_mcs_mat1_7_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7573, mcs1_mcs_mat1_7_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_8998, mcs1_mcs_mat1_7_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_8999, mcs1_mcs_mat1_7_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_8032, mcs1_mcs_mat1_7_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_9325, mcs1_mcs_mat1_7_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_8517, mcs1_mcs_mat1_7_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_7300, shiftr_out[33]}), .c ({new_AGEMA_signal_8999, mcs1_mcs_mat1_7_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_8517, mcs1_mcs_mat1_7_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_8031, mcs1_mcs_mat1_7_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_9000, mcs1_mcs_mat1_7_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_8033, mcs1_mcs_mat1_7_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_7148, mcs1_mcs_mat1_7_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_8517, mcs1_mcs_mat1_7_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_7572, mcs1_mcs_mat1_7_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_8032, mcs1_mcs_mat1_7_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_8518, mcs1_mcs_mat1_7_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_6847, mcs1_mcs_mat1_7_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_7573, mcs1_mcs_mat1_7_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_8032, mcs1_mcs_mat1_7_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_7148, mcs1_mcs_mat1_7_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_7572, mcs1_mcs_mat1_7_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7300, shiftr_out[33]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1039]), .c ({new_AGEMA_signal_8033, mcs1_mcs_mat1_7_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1040]), .c ({new_AGEMA_signal_7148, mcs1_mcs_mat1_7_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1041]), .c ({new_AGEMA_signal_7573, mcs1_mcs_mat1_7_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_8520, mcs1_mcs_mat1_7_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_7149, mcs1_mcs_mat1_7_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_9001, mcs1_mcs_mat1_7_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_7574, mcs1_mcs_mat1_7_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_7575, mcs1_mcs_mat1_7_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_8034, mcs1_mcs_mat1_7_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_8521, mcs1_mcs_mat1_7_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_9002, mcs1_mcs_mat1_7_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_9326, mcs1_mcs_mat1_7_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_8520, mcs1_mcs_mat1_7_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_9002, mcs1_mcs_mat1_7_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_6848, mcs1_mcs_mat1_7_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_8036, mcs1_mcs_mat1_7_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_8520, mcs1_mcs_mat1_7_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_7150, mcs1_mcs_mat1_7_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_8035, mcs1_mcs_mat1_7_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_8521, mcs1_mcs_mat1_7_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7306, shiftr_out[1]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1042]), .c ({new_AGEMA_signal_8036, mcs1_mcs_mat1_7_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1043]), .c ({new_AGEMA_signal_7150, mcs1_mcs_mat1_7_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1044]), .c ({new_AGEMA_signal_7575, mcs1_mcs_mat1_7_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({new_AGEMA_signal_9003, mcs1_mcs_mat1_7_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9327, mcs1_mcs_mat1_7_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({new_AGEMA_signal_9004, mcs1_mcs_mat1_7_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9328, mcs1_mcs_mat1_7_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_7576, mcs1_mcs_mat1_7_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_9003, mcs1_mcs_mat1_7_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_9329, mcs1_mcs_mat1_7_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_7151, mcs1_mcs_mat1_7_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_8522, mcs1_mcs_mat1_7_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_9003, mcs1_mcs_mat1_7_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_8037, mcs1_mcs_mat1_7_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_9004, mcs1_mcs_mat1_7_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_9330, mcs1_mcs_mat1_7_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_8523, mcs1_mcs_mat1_7_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_9004, mcs1_mcs_mat1_7_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_7576, mcs1_mcs_mat1_7_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_8038, mcs1_mcs_mat1_7_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_8523, mcs1_mcs_mat1_7_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1045]), .c ({new_AGEMA_signal_8038, mcs1_mcs_mat1_7_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1046]), .c ({new_AGEMA_signal_7151, mcs1_mcs_mat1_7_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1047]), .c ({new_AGEMA_signal_7576, mcs1_mcs_mat1_7_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_10031, mcs1_mcs_mat1_7_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_10030, mcs1_mcs_mat1_7_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_10254, mcs1_mcs_mat1_7_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_10030, mcs1_mcs_mat1_7_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_9601, mcs1_mcs_mat1_7_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_10255, mcs1_mcs_mat1_7_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_9005, mcs1_mcs_mat1_7_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_9054, shiftr_out[67]}), .c ({new_AGEMA_signal_9601, mcs1_mcs_mat1_7_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_10030, mcs1_mcs_mat1_7_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_9818, mcs1_mcs_mat1_7_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_8524, mcs1_mcs_mat1_7_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_10030, mcs1_mcs_mat1_7_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_10257, mcs1_mcs_mat1_7_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_10497, mcs1_mcs_mat1_7_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_10031, mcs1_mcs_mat1_7_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_9818, mcs1_mcs_mat1_7_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_10257, mcs1_mcs_mat1_7_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_9817, mcs1_mcs_mat1_7_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_7616, shiftr_out[64]}), .c ({new_AGEMA_signal_10031, mcs1_mcs_mat1_7_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_9005, mcs1_mcs_mat1_7_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_9602, mcs1_mcs_mat1_7_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_9817, mcs1_mcs_mat1_7_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1048]), .c ({new_AGEMA_signal_9818, mcs1_mcs_mat1_7_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1049]), .c ({new_AGEMA_signal_9005, mcs1_mcs_mat1_7_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9054, shiftr_out[67]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1050]), .c ({new_AGEMA_signal_9602, mcs1_mcs_mat1_7_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_7577, mcs1_mcs_mat1_7_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_8525, mcs1_mcs_mat1_7_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_9006, mcs1_mcs_mat1_7_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_8042, mcs1_mcs_mat1_7_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_8525, mcs1_mcs_mat1_7_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_8040, mcs1_mcs_mat1_7_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_7578, mcs1_mcs_mat1_7_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_8526, mcs1_mcs_mat1_7_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_8041, mcs1_mcs_mat1_7_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_8527, mcs1_mcs_mat1_7_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_9007, mcs1_mcs_mat1_7_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_6850, mcs1_mcs_mat1_7_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_8042, mcs1_mcs_mat1_7_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_8527, mcs1_mcs_mat1_7_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_7152, mcs1_mcs_mat1_7_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_7300, shiftr_out[33]}), .c ({new_AGEMA_signal_8041, mcs1_mcs_mat1_7_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7300, shiftr_out[33]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1051]), .c ({new_AGEMA_signal_8042, mcs1_mcs_mat1_7_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1052]), .c ({new_AGEMA_signal_7152, mcs1_mcs_mat1_7_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1053]), .c ({new_AGEMA_signal_7578, mcs1_mcs_mat1_7_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_9603, mcs1_mcs_mat1_7_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_7580, mcs1_mcs_mat1_7_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_9819, mcs1_mcs_mat1_7_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_9331, mcs1_mcs_mat1_7_mcs_out[99]}), .b ({new_AGEMA_signal_6694, shiftr_out[2]}), .c ({new_AGEMA_signal_9603, mcs1_mcs_mat1_7_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_9008, mcs1_mcs_mat1_7_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_7306, shiftr_out[1]}), .c ({new_AGEMA_signal_9331, mcs1_mcs_mat1_7_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_8528, mcs1_mcs_mat1_7_mcs_out[98]}), .b ({new_AGEMA_signal_7154, mcs1_mcs_mat1_7_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_9008, mcs1_mcs_mat1_7_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_7153, mcs1_mcs_mat1_7_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_8043, mcs1_mcs_mat1_7_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_8528, mcs1_mcs_mat1_7_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7306, shiftr_out[1]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1054]), .c ({new_AGEMA_signal_8043, mcs1_mcs_mat1_7_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1055]), .c ({new_AGEMA_signal_7154, mcs1_mcs_mat1_7_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1056]), .c ({new_AGEMA_signal_7580, mcs1_mcs_mat1_7_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_8529, mcs1_mcs_mat1_7_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_9009, mcs1_mcs_mat1_7_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_7582, mcs1_mcs_mat1_7_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_7583, mcs1_mcs_mat1_7_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_8045, mcs1_mcs_mat1_7_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_9010, mcs1_mcs_mat1_7_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_7155, mcs1_mcs_mat1_7_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_9332, mcs1_mcs_mat1_7_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_8529, mcs1_mcs_mat1_7_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_9010, mcs1_mcs_mat1_7_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_6852, mcs1_mcs_mat1_7_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_8046, mcs1_mcs_mat1_7_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_8529, mcs1_mcs_mat1_7_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1057]), .c ({new_AGEMA_signal_8046, mcs1_mcs_mat1_7_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1058]), .c ({new_AGEMA_signal_7155, mcs1_mcs_mat1_7_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1059]), .c ({new_AGEMA_signal_7583, mcs1_mcs_mat1_7_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_8050, mcs1_mcs_mat1_7_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_8051, mcs1_mcs_mat1_7_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_8531, mcs1_mcs_mat1_7_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_8048, mcs1_mcs_mat1_7_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_6853, mcs1_mcs_mat1_7_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_8532, mcs1_mcs_mat1_7_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_7584, mcs1_mcs_mat1_7_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_8048, mcs1_mcs_mat1_7_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_8049, mcs1_mcs_mat1_7_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_8533, mcs1_mcs_mat1_7_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_7156, mcs1_mcs_mat1_7_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_7584, mcs1_mcs_mat1_7_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_8049, mcs1_mcs_mat1_7_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_8534, mcs1_mcs_mat1_7_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_6694, shiftr_out[2]}), .c ({new_AGEMA_signal_9011, mcs1_mcs_mat1_7_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_8050, mcs1_mcs_mat1_7_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_7156, mcs1_mcs_mat1_7_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_8534, mcs1_mcs_mat1_7_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7306, shiftr_out[1]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1060]), .c ({new_AGEMA_signal_8051, mcs1_mcs_mat1_7_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1061]), .c ({new_AGEMA_signal_7156, mcs1_mcs_mat1_7_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1062]), .c ({new_AGEMA_signal_7584, mcs1_mcs_mat1_7_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_8535, mcs1_mcs_mat1_7_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_9012, mcs1_mcs_mat1_7_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_7585, mcs1_mcs_mat1_7_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_8052, mcs1_mcs_mat1_7_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_9013, mcs1_mcs_mat1_7_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_7158, mcs1_mcs_mat1_7_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_9333, mcs1_mcs_mat1_7_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_8535, mcs1_mcs_mat1_7_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_6608, shiftr_out[96]}), .c ({new_AGEMA_signal_9013, mcs1_mcs_mat1_7_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_6854, mcs1_mcs_mat1_7_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_8053, mcs1_mcs_mat1_7_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_8535, mcs1_mcs_mat1_7_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1063]), .c ({new_AGEMA_signal_8053, mcs1_mcs_mat1_7_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1064]), .c ({new_AGEMA_signal_7158, mcs1_mcs_mat1_7_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1065]), .c ({new_AGEMA_signal_7585, mcs1_mcs_mat1_7_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_10258, mcs1_mcs_mat1_7_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_10498, mcs1_mcs_mat1_7_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_10033, mcs1_mcs_mat1_7_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9821, mcs1_mcs_mat1_7_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_10258, mcs1_mcs_mat1_7_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_9334, mcs1_mcs_mat1_7_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_9820, mcs1_mcs_mat1_7_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_9821, mcs1_mcs_mat1_7_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_9334, mcs1_mcs_mat1_7_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_10032, mcs1_mcs_mat1_7_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_9014, mcs1_mcs_mat1_7_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_9015, mcs1_mcs_mat1_7_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_9334, mcs1_mcs_mat1_7_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_9606, mcs1_mcs_mat1_7_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_7616, shiftr_out[64]}), .c ({new_AGEMA_signal_9821, mcs1_mcs_mat1_7_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_10259, mcs1_mcs_mat1_7_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_9014, mcs1_mcs_mat1_7_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_10499, mcs1_mcs_mat1_7_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_10033, mcs1_mcs_mat1_7_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9606, mcs1_mcs_mat1_7_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_10259, mcs1_mcs_mat1_7_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_9054, shiftr_out[67]}), .b ({new_AGEMA_signal_9822, mcs1_mcs_mat1_7_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_10033, mcs1_mcs_mat1_7_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1066]), .c ({new_AGEMA_signal_9822, mcs1_mcs_mat1_7_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1067]), .c ({new_AGEMA_signal_9015, mcs1_mcs_mat1_7_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9054, shiftr_out[67]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1068]), .c ({new_AGEMA_signal_9606, mcs1_mcs_mat1_7_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_8537, mcs1_mcs_mat1_7_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_7586, mcs1_mcs_mat1_7_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_9016, mcs1_mcs_mat1_7_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_8055, mcs1_mcs_mat1_7_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_9017, mcs1_mcs_mat1_7_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9335, mcs1_mcs_mat1_7_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_8537, mcs1_mcs_mat1_7_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_9017, mcs1_mcs_mat1_7_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_9336, mcs1_mcs_mat1_7_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_7586, mcs1_mcs_mat1_7_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_8538, mcs1_mcs_mat1_7_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_9017, mcs1_mcs_mat1_7_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({new_AGEMA_signal_7159, mcs1_mcs_mat1_7_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_7586, mcs1_mcs_mat1_7_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_8054, mcs1_mcs_mat1_7_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_7300, shiftr_out[33]}), .c ({new_AGEMA_signal_8537, mcs1_mcs_mat1_7_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_7587, mcs1_mcs_mat1_7_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6855, mcs1_mcs_mat1_7_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_8054, mcs1_mcs_mat1_7_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_8538, mcs1_mcs_mat1_7_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_8055, mcs1_mcs_mat1_7_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_9018, mcs1_mcs_mat1_7_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_7587, mcs1_mcs_mat1_7_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_8055, mcs1_mcs_mat1_7_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({new_AGEMA_signal_8056, mcs1_mcs_mat1_7_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_8538, mcs1_mcs_mat1_7_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7300, shiftr_out[33]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1069]), .c ({new_AGEMA_signal_8056, mcs1_mcs_mat1_7_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1070]), .c ({new_AGEMA_signal_7159, mcs1_mcs_mat1_7_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1071]), .c ({new_AGEMA_signal_7587, mcs1_mcs_mat1_7_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_9020, mcs1_mcs_mat1_7_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_9337, mcs1_mcs_mat1_7_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({new_AGEMA_signal_8539, mcs1_mcs_mat1_7_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_9019, mcs1_mcs_mat1_7_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_9338, mcs1_mcs_mat1_7_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_7588, mcs1_mcs_mat1_7_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_9607, mcs1_mcs_mat1_7_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_9020, mcs1_mcs_mat1_7_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .c ({new_AGEMA_signal_9338, mcs1_mcs_mat1_7_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_7160, mcs1_mcs_mat1_7_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_8539, mcs1_mcs_mat1_7_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_9020, mcs1_mcs_mat1_7_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_6856, mcs1_mcs_mat1_7_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_8058, mcs1_mcs_mat1_7_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_8539, mcs1_mcs_mat1_7_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7306, shiftr_out[1]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1072]), .c ({new_AGEMA_signal_8058, mcs1_mcs_mat1_7_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1073]), .c ({new_AGEMA_signal_7160, mcs1_mcs_mat1_7_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1074]), .c ({new_AGEMA_signal_7588, mcs1_mcs_mat1_7_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_8542, mcs1_mcs_mat1_7_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_7589, mcs1_mcs_mat1_7_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_9021, mcs1_mcs_mat1_7_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_7161, mcs1_mcs_mat1_7_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_8059, mcs1_mcs_mat1_7_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_8540, mcs1_mcs_mat1_7_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({new_AGEMA_signal_8060, mcs1_mcs_mat1_7_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_8541, mcs1_mcs_mat1_7_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1075]), .c ({new_AGEMA_signal_8060, mcs1_mcs_mat1_7_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1076]), .c ({new_AGEMA_signal_7161, mcs1_mcs_mat1_7_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1077]), .c ({new_AGEMA_signal_7589, mcs1_mcs_mat1_7_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_9024, mcs1_mcs_mat1_7_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_9608, mcs1_mcs_mat1_7_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_9823, mcs1_mcs_mat1_7_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_9025, mcs1_mcs_mat1_7_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_9824, mcs1_mcs_mat1_7_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_10035, mcs1_mcs_mat1_7_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_10036, mcs1_mcs_mat1_7_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_9825, mcs1_mcs_mat1_7_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_10260, mcs1_mcs_mat1_7_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_9826, mcs1_mcs_mat1_7_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_10036, mcs1_mcs_mat1_7_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1078]), .c ({new_AGEMA_signal_9826, mcs1_mcs_mat1_7_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1079]), .c ({new_AGEMA_signal_9025, mcs1_mcs_mat1_7_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9054, shiftr_out[67]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1080]), .c ({new_AGEMA_signal_9608, mcs1_mcs_mat1_7_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_8062, mcs1_mcs_mat1_7_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8544, mcs1_mcs_mat1_7_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_9026, mcs1_mcs_mat1_7_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_9027, mcs1_mcs_mat1_7_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_8061, mcs1_mcs_mat1_7_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_9340, mcs1_mcs_mat1_7_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_7590, mcs1_mcs_mat1_7_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_8061, mcs1_mcs_mat1_7_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({new_AGEMA_signal_9027, mcs1_mcs_mat1_7_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_9341, mcs1_mcs_mat1_7_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_6858, mcs1_mcs_mat1_7_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_8544, mcs1_mcs_mat1_7_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_9027, mcs1_mcs_mat1_7_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_7162, mcs1_mcs_mat1_7_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_8064, mcs1_mcs_mat1_7_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_8544, mcs1_mcs_mat1_7_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_8063, mcs1_mcs_mat1_7_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_8545, mcs1_mcs_mat1_7_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_9028, mcs1_mcs_mat1_7_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_8062, mcs1_mcs_mat1_7_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_7162, mcs1_mcs_mat1_7_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_8545, mcs1_mcs_mat1_7_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_7590, mcs1_mcs_mat1_7_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_8062, mcs1_mcs_mat1_7_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7300, shiftr_out[33]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1081]), .c ({new_AGEMA_signal_8064, mcs1_mcs_mat1_7_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1082]), .c ({new_AGEMA_signal_7162, mcs1_mcs_mat1_7_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1083]), .c ({new_AGEMA_signal_7590, mcs1_mcs_mat1_7_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_7592, mcs1_mcs_mat1_7_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_8066, mcs1_mcs_mat1_7_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_9342, mcs1_mcs_mat1_7_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_7163, mcs1_mcs_mat1_7_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_9609, mcs1_mcs_mat1_7_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_9029, mcs1_mcs_mat1_7_mcs_out[47]}), .b ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_9342, mcs1_mcs_mat1_7_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_8547, mcs1_mcs_mat1_7_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_6608, shiftr_out[96]}), .c ({new_AGEMA_signal_9029, mcs1_mcs_mat1_7_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_6859, mcs1_mcs_mat1_7_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_8067, mcs1_mcs_mat1_7_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_8547, mcs1_mcs_mat1_7_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1084]), .c ({new_AGEMA_signal_8067, mcs1_mcs_mat1_7_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1085]), .c ({new_AGEMA_signal_7163, mcs1_mcs_mat1_7_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1086]), .c ({new_AGEMA_signal_7592, mcs1_mcs_mat1_7_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_10037, mcs1_mcs_mat1_7_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_9610, mcs1_mcs_mat1_7_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_10261, mcs1_mcs_mat1_7_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_9827, mcs1_mcs_mat1_7_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9030, mcs1_mcs_mat1_7_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_10037, mcs1_mcs_mat1_7_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_10038, mcs1_mcs_mat1_7_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_9829, mcs1_mcs_mat1_7_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_10262, mcs1_mcs_mat1_7_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_10039, mcs1_mcs_mat1_7_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_8548, mcs1_mcs_mat1_7_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_10263, mcs1_mcs_mat1_7_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_9827, mcs1_mcs_mat1_7_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9611, mcs1_mcs_mat1_7_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_10039, mcs1_mcs_mat1_7_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_9828, mcs1_mcs_mat1_7_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_9611, mcs1_mcs_mat1_7_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_10040, mcs1_mcs_mat1_7_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1087]), .c ({new_AGEMA_signal_9829, mcs1_mcs_mat1_7_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1088]), .c ({new_AGEMA_signal_9030, mcs1_mcs_mat1_7_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9054, shiftr_out[67]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1089]), .c ({new_AGEMA_signal_9611, mcs1_mcs_mat1_7_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_9031, mcs1_mcs_mat1_7_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_6860, mcs1_mcs_mat1_7_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9343, mcs1_mcs_mat1_7_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_7594, mcs1_mcs_mat1_7_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_7593, mcs1_mcs_mat1_7_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_8068, mcs1_mcs_mat1_7_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({new_AGEMA_signal_9031, mcs1_mcs_mat1_7_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_9344, mcs1_mcs_mat1_7_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_8069, mcs1_mcs_mat1_7_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_8549, mcs1_mcs_mat1_7_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_9031, mcs1_mcs_mat1_7_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_8070, mcs1_mcs_mat1_7_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7595, mcs1_mcs_mat1_7_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_8549, mcs1_mcs_mat1_7_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_8070, mcs1_mcs_mat1_7_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_7594, mcs1_mcs_mat1_7_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_8550, mcs1_mcs_mat1_7_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_7273, mcs1_mcs_mat1_7_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_7594, mcs1_mcs_mat1_7_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({new_AGEMA_signal_7164, mcs1_mcs_mat1_7_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_7273, mcs1_mcs_mat1_7_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7300, shiftr_out[33]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1090]), .c ({new_AGEMA_signal_8070, mcs1_mcs_mat1_7_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1091]), .c ({new_AGEMA_signal_7164, mcs1_mcs_mat1_7_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1092]), .c ({new_AGEMA_signal_7595, mcs1_mcs_mat1_7_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_8071, mcs1_mcs_mat1_7_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7596, mcs1_mcs_mat1_7_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_8551, mcs1_mcs_mat1_7_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_7165, mcs1_mcs_mat1_7_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_7274, mcs1_mcs_mat1_7_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_9345, mcs1_mcs_mat1_7_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_8072, mcs1_mcs_mat1_7_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_9612, mcs1_mcs_mat1_7_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7306, shiftr_out[1]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1093]), .c ({new_AGEMA_signal_8072, mcs1_mcs_mat1_7_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1094]), .c ({new_AGEMA_signal_7165, mcs1_mcs_mat1_7_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1095]), .c ({new_AGEMA_signal_7596, mcs1_mcs_mat1_7_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_9033, mcs1_mcs_mat1_7_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_8553, mcs1_mcs_mat1_7_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_9346, mcs1_mcs_mat1_7_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_7167, mcs1_mcs_mat1_7_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_8554, mcs1_mcs_mat1_7_mcs_out[29]}), .c ({new_AGEMA_signal_9033, mcs1_mcs_mat1_7_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_7166, mcs1_mcs_mat1_7_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_8553, mcs1_mcs_mat1_7_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_9034, mcs1_mcs_mat1_7_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_8075, mcs1_mcs_mat1_7_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_6608, shiftr_out[96]}), .c ({new_AGEMA_signal_8553, mcs1_mcs_mat1_7_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_9035, mcs1_mcs_mat1_7_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_8073, mcs1_mcs_mat1_7_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_9347, mcs1_mcs_mat1_7_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_8555, mcs1_mcs_mat1_7_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_8074, mcs1_mcs_mat1_7_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_9035, mcs1_mcs_mat1_7_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_7597, mcs1_mcs_mat1_7_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_8074, mcs1_mcs_mat1_7_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_8075, mcs1_mcs_mat1_7_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7167, mcs1_mcs_mat1_7_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_8555, mcs1_mcs_mat1_7_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1096]), .c ({new_AGEMA_signal_8075, mcs1_mcs_mat1_7_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1097]), .c ({new_AGEMA_signal_7167, mcs1_mcs_mat1_7_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1098]), .c ({new_AGEMA_signal_7597, mcs1_mcs_mat1_7_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_9830, mcs1_mcs_mat1_7_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_10041, mcs1_mcs_mat1_7_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_9613, mcs1_mcs_mat1_7_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_9036, mcs1_mcs_mat1_7_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_9830, mcs1_mcs_mat1_7_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_10042, mcs1_mcs_mat1_7_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_10264, mcs1_mcs_mat1_7_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_9832, mcs1_mcs_mat1_7_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_9036, mcs1_mcs_mat1_7_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_10042, mcs1_mcs_mat1_7_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_10265, mcs1_mcs_mat1_7_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_7616, shiftr_out[64]}), .c ({new_AGEMA_signal_10500, mcs1_mcs_mat1_7_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_9832, mcs1_mcs_mat1_7_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_10043, mcs1_mcs_mat1_7_mcs_out[24]}), .c ({new_AGEMA_signal_10265, mcs1_mcs_mat1_7_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_9831, mcs1_mcs_mat1_7_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_9054, shiftr_out[67]}), .c ({new_AGEMA_signal_10043, mcs1_mcs_mat1_7_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_9613, mcs1_mcs_mat1_7_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8556, mcs1_mcs_mat1_7_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_9831, mcs1_mcs_mat1_7_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1099]), .c ({new_AGEMA_signal_9832, mcs1_mcs_mat1_7_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1100]), .c ({new_AGEMA_signal_9036, mcs1_mcs_mat1_7_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9054, shiftr_out[67]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1101]), .c ({new_AGEMA_signal_9613, mcs1_mcs_mat1_7_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_8076, mcs1_mcs_mat1_7_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_6688, shiftr_out[34]}), .c ({new_AGEMA_signal_8557, mcs1_mcs_mat1_7_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_7598, mcs1_mcs_mat1_7_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7168, mcs1_mcs_mat1_7_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_8076, mcs1_mcs_mat1_7_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_8558, mcs1_mcs_mat1_7_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_7300, shiftr_out[33]}), .c ({new_AGEMA_signal_9037, mcs1_mcs_mat1_7_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_8078, mcs1_mcs_mat1_7_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_7168, mcs1_mcs_mat1_7_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_8558, mcs1_mcs_mat1_7_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_9038, mcs1_mcs_mat1_7_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_6620, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_9348, mcs1_mcs_mat1_7_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_8078, mcs1_mcs_mat1_7_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8559, mcs1_mcs_mat1_7_mcs_out[20]}), .c ({new_AGEMA_signal_9038, mcs1_mcs_mat1_7_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_8077, mcs1_mcs_mat1_7_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_8559, mcs1_mcs_mat1_7_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_7598, mcs1_mcs_mat1_7_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_6863, mcs1_mcs_mat1_7_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_8077, mcs1_mcs_mat1_7_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7300, shiftr_out[33]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1102]), .c ({new_AGEMA_signal_8078, mcs1_mcs_mat1_7_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1103]), .c ({new_AGEMA_signal_7168, mcs1_mcs_mat1_7_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1104]), .c ({new_AGEMA_signal_7598, mcs1_mcs_mat1_7_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_8079, mcs1_mcs_mat1_7_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_8082, mcs1_mcs_mat1_7_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_8560, mcs1_mcs_mat1_7_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_8561, mcs1_mcs_mat1_7_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_6864, mcs1_mcs_mat1_7_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_9039, mcs1_mcs_mat1_7_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_9040, mcs1_mcs_mat1_7_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_7169, mcs1_mcs_mat1_7_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_9349, mcs1_mcs_mat1_7_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_6626, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_8561, mcs1_mcs_mat1_7_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_9040, mcs1_mcs_mat1_7_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_8080, mcs1_mcs_mat1_7_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_7306, shiftr_out[1]}), .c ({new_AGEMA_signal_8561, mcs1_mcs_mat1_7_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_7599, mcs1_mcs_mat1_7_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_7600, mcs1_mcs_mat1_7_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_8080, mcs1_mcs_mat1_7_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_8081, mcs1_mcs_mat1_7_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_7169, mcs1_mcs_mat1_7_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_8562, mcs1_mcs_mat1_7_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7306, shiftr_out[1]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1105]), .c ({new_AGEMA_signal_8082, mcs1_mcs_mat1_7_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1106]), .c ({new_AGEMA_signal_7169, mcs1_mcs_mat1_7_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1107]), .c ({new_AGEMA_signal_7600, mcs1_mcs_mat1_7_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_9043, mcs1_mcs_mat1_7_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_7275, mcs1_mcs_mat1_7_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_9350, mcs1_mcs_mat1_7_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_8565, mcs1_mcs_mat1_7_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_8563, mcs1_mcs_mat1_7_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_9041, mcs1_mcs_mat1_7_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_8084, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_7170, mcs1_mcs_mat1_7_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8563, mcs1_mcs_mat1_7_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_7275, mcs1_mcs_mat1_7_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_9042, mcs1_mcs_mat1_7_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_8083, mcs1_mcs_mat1_7_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_8084, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_6865, mcs1_mcs_mat1_7_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_7170, mcs1_mcs_mat1_7_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_7275, mcs1_mcs_mat1_7_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_9351, mcs1_mcs_mat1_7_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_9614, mcs1_mcs_mat1_7_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_9043, mcs1_mcs_mat1_7_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_8084, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_9351, mcs1_mcs_mat1_7_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_8565, mcs1_mcs_mat1_7_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_9043, mcs1_mcs_mat1_7_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_8083, mcs1_mcs_mat1_7_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_8565, mcs1_mcs_mat1_7_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_6608, shiftr_out[96]}), .b ({new_AGEMA_signal_7601, mcs1_mcs_mat1_7_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_8083, mcs1_mcs_mat1_7_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7288, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1108]), .c ({new_AGEMA_signal_8084, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6676, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1109]), .c ({new_AGEMA_signal_7170, mcs1_mcs_mat1_7_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7222, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1110]), .c ({new_AGEMA_signal_7601, mcs1_mcs_mat1_7_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_9352, mcs1_mcs_mat1_7_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_9054, shiftr_out[67]}), .c ({new_AGEMA_signal_9615, mcs1_mcs_mat1_7_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_10045, mcs1_mcs_mat1_7_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_10266, mcs1_mcs_mat1_7_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_9833, mcs1_mcs_mat1_7_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_10044, mcs1_mcs_mat1_7_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_9616, mcs1_mcs_mat1_7_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_9352, mcs1_mcs_mat1_7_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_9833, mcs1_mcs_mat1_7_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_8566, mcs1_mcs_mat1_7_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_9044, mcs1_mcs_mat1_7_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_9352, mcs1_mcs_mat1_7_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_10267, mcs1_mcs_mat1_7_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_7616, shiftr_out[64]}), .c ({new_AGEMA_signal_10501, mcs1_mcs_mat1_7_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_8566, mcs1_mcs_mat1_7_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_10045, mcs1_mcs_mat1_7_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_10267, mcs1_mcs_mat1_7_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_9834, mcs1_mcs_mat1_7_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_9616, mcs1_mcs_mat1_7_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_10045, mcs1_mcs_mat1_7_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_9358, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1111]), .c ({new_AGEMA_signal_9834, mcs1_mcs_mat1_7_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8096, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1112]), .c ({new_AGEMA_signal_9044, mcs1_mcs_mat1_7_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_9054, shiftr_out[67]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1113]), .c ({new_AGEMA_signal_9616, mcs1_mcs_mat1_7_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_9617, mcs1_mcs_mat1_7_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_7603, mcs1_mcs_mat1_7_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_9835, mcs1_mcs_mat1_7_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_9353, mcs1_mcs_mat1_7_mcs_out[7]}), .b ({new_AGEMA_signal_6688, shiftr_out[34]}), .c ({new_AGEMA_signal_9617, mcs1_mcs_mat1_7_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_9045, mcs1_mcs_mat1_7_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_7300, shiftr_out[33]}), .c ({new_AGEMA_signal_9353, mcs1_mcs_mat1_7_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_8567, mcs1_mcs_mat1_7_mcs_out[6]}), .b ({new_AGEMA_signal_7172, mcs1_mcs_mat1_7_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_9045, mcs1_mcs_mat1_7_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_7171, mcs1_mcs_mat1_7_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_8085, mcs1_mcs_mat1_7_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_8567, mcs1_mcs_mat1_7_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7300, shiftr_out[33]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1114]), .c ({new_AGEMA_signal_8085, mcs1_mcs_mat1_7_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6688, shiftr_out[34]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1115]), .c ({new_AGEMA_signal_7172, mcs1_mcs_mat1_7_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7234, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1116]), .c ({new_AGEMA_signal_7603, mcs1_mcs_mat1_7_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_7604, mcs1_mcs_mat1_7_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_8086, mcs1_mcs_mat1_7_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_8569, mcs1_mcs_mat1_7_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_7306, shiftr_out[1]}), .b ({new_AGEMA_signal_7605, mcs1_mcs_mat1_7_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_8086, mcs1_mcs_mat1_7_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_8570, mcs1_mcs_mat1_7_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_7173, mcs1_mcs_mat1_7_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_9046, mcs1_mcs_mat1_7_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_8571, mcs1_mcs_mat1_7_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_8088, mcs1_mcs_mat1_7_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_9047, mcs1_mcs_mat1_7_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_8089, mcs1_mcs_mat1_7_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_6867, mcs1_mcs_mat1_7_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_8571, mcs1_mcs_mat1_7_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_7306, shiftr_out[1]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1117]), .c ({new_AGEMA_signal_8089, mcs1_mcs_mat1_7_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_6694, shiftr_out[2]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1118]), .c ({new_AGEMA_signal_7173, mcs1_mcs_mat1_7_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_7240, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, p256_sel}), .clk (clk), .r (Fresh[1119]), .c ({new_AGEMA_signal_7605, mcs1_mcs_mat1_7_mcs_rom0_31_x3x4}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10936, mcs_out[128]}), .a ({new_AGEMA_signal_10956, y0_1[0]}), .c ({y0_s1[0], y0_s0[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10489, mcs_out[129]}), .a ({new_AGEMA_signal_10519, y0_1[1]}), .c ({y0_s1[1], y0_s0[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10935, mcs_out[130]}), .a ({new_AGEMA_signal_10973, y0_1[2]}), .c ({y0_s1[2], y0_s0[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10246, mcs_out[131]}), .a ({new_AGEMA_signal_10286, y0_1[3]}), .c ({y0_s1[3], y0_s0[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10722, mcs_out[132]}), .a ({new_AGEMA_signal_10777, y0_1[4]}), .c ({y0_s1[4], y0_s0[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10926, mcs_out[133]}), .a ({new_AGEMA_signal_10975, y0_1[5]}), .c ({y0_s1[5], y0_s0[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10925, mcs_out[134]}), .a ({new_AGEMA_signal_10978, y0_1[6]}), .c ({y0_s1[6], y0_s0[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10719, mcs_out[135]}), .a ({new_AGEMA_signal_10785, y0_1[7]}), .c ({y0_s1[7], y0_s0[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11054, mcs_out[136]}), .a ({new_AGEMA_signal_11085, y0_1[8]}), .c ({y0_s1[8], y0_s0[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10201, mcs_out[137]}), .a ({new_AGEMA_signal_10295, y0_1[9]}), .c ({y0_s1[9], y0_s0[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10704, mcs_out[138]}), .a ({new_AGEMA_signal_10766, y0_1[10]}), .c ({y0_s1[10], y0_s0[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10917, mcs_out[139]}), .a ({new_AGEMA_signal_10964, y0_1[11]}), .c ({y0_s1[11], y0_s0[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10910, mcs_out[140]}), .a ({new_AGEMA_signal_10966, y0_1[12]}), .c ({y0_s1[12], y0_s0[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10173, mcs_out[141]}), .a ({new_AGEMA_signal_10281, y0_1[13]}), .c ({y0_s1[13], y0_s0[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9732, mcs_out[142]}), .a ({new_AGEMA_signal_9842, y0_1[14]}), .c ({y0_s1[14], y0_s0[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10689, mcs_out[143]}), .a ({new_AGEMA_signal_10770, y0_1[15]}), .c ({y0_s1[15], y0_s0[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10899, mcs_out[144]}), .a ({new_AGEMA_signal_10967, y0_1[16]}), .c ({y0_s1[16], y0_s0[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10394, mcs_out[145]}), .a ({new_AGEMA_signal_10518, y0_1[17]}), .c ({y0_s1[17], y0_s0[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10898, mcs_out[146]}), .a ({new_AGEMA_signal_10968, y0_1[18]}), .c ({y0_s1[18], y0_s0[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10147, mcs_out[147]}), .a ({new_AGEMA_signal_10282, y0_1[19]}), .c ({y0_s1[19], y0_s0[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10653, mcs_out[148]}), .a ({new_AGEMA_signal_10771, y0_1[20]}), .c ({y0_s1[20], y0_s0[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10889, mcs_out[149]}), .a ({new_AGEMA_signal_10969, y0_1[21]}), .c ({y0_s1[21], y0_s0[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10888, mcs_out[150]}), .a ({new_AGEMA_signal_10970, y0_1[22]}), .c ({y0_s1[22], y0_s0[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10650, mcs_out[151]}), .a ({new_AGEMA_signal_10772, y0_1[23]}), .c ({y0_s1[23], y0_s0[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11048, mcs_out[152]}), .a ({new_AGEMA_signal_11084, y0_1[24]}), .c ({y0_s1[24], y0_s0[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10102, mcs_out[153]}), .a ({new_AGEMA_signal_10283, y0_1[25]}), .c ({y0_s1[25], y0_s0[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10635, mcs_out[154]}), .a ({new_AGEMA_signal_10773, y0_1[26]}), .c ({y0_s1[26], y0_s0[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10880, mcs_out[155]}), .a ({new_AGEMA_signal_10971, y0_1[27]}), .c ({y0_s1[27], y0_s0[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10873, mcs_out[156]}), .a ({new_AGEMA_signal_10972, y0_1[28]}), .c ({y0_s1[28], y0_s0[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10074, mcs_out[157]}), .a ({new_AGEMA_signal_10284, y0_1[29]}), .c ({y0_s1[29], y0_s0[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9623, mcs_out[158]}), .a ({new_AGEMA_signal_9843, y0_1[30]}), .c ({y0_s1[30], y0_s0[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10620, mcs_out[159]}), .a ({new_AGEMA_signal_10774, y0_1[31]}), .c ({y0_s1[31], y0_s0[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_32_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9812, mcs_out[160]}), .a ({new_AGEMA_signal_9844, y0_1[32]}), .c ({y0_s1[32], y0_s0[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_33_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10025, mcs_out[161]}), .a ({new_AGEMA_signal_10050, y0_1[33]}), .c ({y0_s1[33], y0_s0[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_34_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10024, mcs_out[162]}), .a ({new_AGEMA_signal_10051, y0_1[34]}), .c ({y0_s1[34], y0_s0[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_35_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10023, mcs_out[163]}), .a ({new_AGEMA_signal_10052, y0_1[35]}), .c ({y0_s1[35], y0_s0[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_36_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10463, mcs_out[164]}), .a ({new_AGEMA_signal_10520, y0_1[36]}), .c ({y0_s1[36], y0_s0[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_37_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9781, mcs_out[165]}), .a ({new_AGEMA_signal_9845, y0_1[37]}), .c ({y0_s1[37], y0_s0[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_38_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9286, mcs_out[166]}), .a ({new_AGEMA_signal_9354, y0_1[38]}), .c ({y0_s1[38], y0_s0[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_39_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10223, mcs_out[167]}), .a ({new_AGEMA_signal_10285, y0_1[39]}), .c ({y0_s1[39], y0_s0[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_40_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10701, mcs_out[168]}), .a ({new_AGEMA_signal_10775, y0_1[40]}), .c ({y0_s1[40], y0_s0[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_41_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10439, mcs_out[169]}), .a ({new_AGEMA_signal_10521, y0_1[41]}), .c ({y0_s1[41], y0_s0[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_42_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10438, mcs_out[170]}), .a ({new_AGEMA_signal_10522, y0_1[42]}), .c ({y0_s1[42], y0_s0[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_43_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10437, mcs_out[171]}), .a ({new_AGEMA_signal_10523, y0_1[43]}), .c ({y0_s1[43], y0_s0[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_44_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10909, mcs_out[172]}), .a ({new_AGEMA_signal_10974, y0_1[44]}), .c ({y0_s1[44], y0_s0[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_45_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10172, mcs_out[173]}), .a ({new_AGEMA_signal_10287, y0_1[45]}), .c ({y0_s1[45], y0_s0[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_46_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10171, mcs_out[174]}), .a ({new_AGEMA_signal_10288, y0_1[46]}), .c ({y0_s1[46], y0_s0[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_47_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10686, mcs_out[175]}), .a ({new_AGEMA_signal_10776, y0_1[47]}), .c ({y0_s1[47], y0_s0[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_48_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9703, mcs_out[176]}), .a ({new_AGEMA_signal_9846, y0_1[48]}), .c ({y0_s1[48], y0_s0[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_49_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9932, mcs_out[177]}), .a ({new_AGEMA_signal_10053, y0_1[49]}), .c ({y0_s1[49], y0_s0[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_50_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9931, mcs_out[178]}), .a ({new_AGEMA_signal_10054, y0_1[50]}), .c ({y0_s1[50], y0_s0[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_51_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9930, mcs_out[179]}), .a ({new_AGEMA_signal_10055, y0_1[51]}), .c ({y0_s1[51], y0_s0[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_52_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10368, mcs_out[180]}), .a ({new_AGEMA_signal_10524, y0_1[52]}), .c ({y0_s1[52], y0_s0[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_53_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9672, mcs_out[181]}), .a ({new_AGEMA_signal_9847, y0_1[53]}), .c ({y0_s1[53], y0_s0[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_54_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9139, mcs_out[182]}), .a ({new_AGEMA_signal_9355, y0_1[54]}), .c ({y0_s1[54], y0_s0[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_55_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10124, mcs_out[183]}), .a ({new_AGEMA_signal_10289, y0_1[55]}), .c ({y0_s1[55], y0_s0[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_56_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10632, mcs_out[184]}), .a ({new_AGEMA_signal_10778, y0_1[56]}), .c ({y0_s1[56], y0_s0[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_57_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10344, mcs_out[185]}), .a ({new_AGEMA_signal_10525, y0_1[57]}), .c ({y0_s1[57], y0_s0[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_58_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10343, mcs_out[186]}), .a ({new_AGEMA_signal_10526, y0_1[58]}), .c ({y0_s1[58], y0_s0[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_59_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10342, mcs_out[187]}), .a ({new_AGEMA_signal_10527, y0_1[59]}), .c ({y0_s1[59], y0_s0[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_60_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10872, mcs_out[188]}), .a ({new_AGEMA_signal_10976, y0_1[60]}), .c ({y0_s1[60], y0_s0[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_61_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10073, mcs_out[189]}), .a ({new_AGEMA_signal_10290, y0_1[61]}), .c ({y0_s1[61], y0_s0[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_62_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10072, mcs_out[190]}), .a ({new_AGEMA_signal_10291, y0_1[62]}), .c ({y0_s1[62], y0_s0[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_63_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10617, mcs_out[191]}), .a ({new_AGEMA_signal_10779, y0_1[63]}), .c ({y0_s1[63], y0_s0[63]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_64_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10934, mcs_out[192]}), .a ({new_AGEMA_signal_10977, y0_1[64]}), .c ({y0_s1[64], y0_s0[64]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_65_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10738, mcs_out[193]}), .a ({new_AGEMA_signal_10780, y0_1[65]}), .c ({y0_s1[65], y0_s0[65]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_66_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10737, mcs_out[194]}), .a ({new_AGEMA_signal_10781, y0_1[66]}), .c ({y0_s1[66], y0_s0[66]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_67_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10736, mcs_out[195]}), .a ({new_AGEMA_signal_10782, y0_1[67]}), .c ({y0_s1[67], y0_s0[67]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_68_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10718, mcs_out[196]}), .a ({new_AGEMA_signal_10783, y0_1[68]}), .c ({y0_s1[68], y0_s0[68]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_69_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10461, mcs_out[197]}), .a ({new_AGEMA_signal_10528, y0_1[69]}), .c ({y0_s1[69], y0_s0[69]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_70_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10221, mcs_out[198]}), .a ({new_AGEMA_signal_10292, y0_1[70]}), .c ({y0_s1[70], y0_s0[70]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_71_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10717, mcs_out[199]}), .a ({new_AGEMA_signal_10784, y0_1[71]}), .c ({y0_s1[71], y0_s0[71]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_72_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11100, mcs_out[200]}), .a ({new_AGEMA_signal_11138, y0_1[72]}), .c ({y0_s1[72], y0_s0[72]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_73_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9976, mcs_out[201]}), .a ({new_AGEMA_signal_10056, y0_1[73]}), .c ({y0_s1[73], y0_s0[73]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_74_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10436, mcs_out[202]}), .a ({new_AGEMA_signal_10529, y0_1[74]}), .c ({y0_s1[74], y0_s0[74]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_75_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10916, mcs_out[203]}), .a ({new_AGEMA_signal_10979, y0_1[75]}), .c ({y0_s1[75], y0_s0[75]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_76_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10908, mcs_out[204]}), .a ({new_AGEMA_signal_10980, y0_1[76]}), .c ({y0_s1[76], y0_s0[76]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_77_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10907, mcs_out[205]}), .a ({new_AGEMA_signal_10981, y0_1[77]}), .c ({y0_s1[77], y0_s0[77]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_78_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10906, mcs_out[206]}), .a ({new_AGEMA_signal_10982, y0_1[78]}), .c ({y0_s1[78], y0_s0[78]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_79_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10905, mcs_out[207]}), .a ({new_AGEMA_signal_10983, y0_1[79]}), .c ({y0_s1[79], y0_s0[79]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_80_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10897, mcs_out[208]}), .a ({new_AGEMA_signal_10984, y0_1[80]}), .c ({y0_s1[80], y0_s0[80]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_81_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10669, mcs_out[209]}), .a ({new_AGEMA_signal_10786, y0_1[81]}), .c ({y0_s1[81], y0_s0[81]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_82_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10668, mcs_out[210]}), .a ({new_AGEMA_signal_10787, y0_1[82]}), .c ({y0_s1[82], y0_s0[82]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_83_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10667, mcs_out[211]}), .a ({new_AGEMA_signal_10788, y0_1[83]}), .c ({y0_s1[83], y0_s0[83]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_84_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10649, mcs_out[212]}), .a ({new_AGEMA_signal_10789, y0_1[84]}), .c ({y0_s1[84], y0_s0[84]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_85_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10366, mcs_out[213]}), .a ({new_AGEMA_signal_10530, y0_1[85]}), .c ({y0_s1[85], y0_s0[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_86_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10122, mcs_out[214]}), .a ({new_AGEMA_signal_10293, y0_1[86]}), .c ({y0_s1[86], y0_s0[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_87_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10648, mcs_out[215]}), .a ({new_AGEMA_signal_10790, y0_1[87]}), .c ({y0_s1[87], y0_s0[87]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_88_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11098, mcs_out[216]}), .a ({new_AGEMA_signal_11139, y0_1[88]}), .c ({y0_s1[88], y0_s0[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_89_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9883, mcs_out[217]}), .a ({new_AGEMA_signal_10057, y0_1[89]}), .c ({y0_s1[89], y0_s0[89]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_90_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10341, mcs_out[218]}), .a ({new_AGEMA_signal_10531, y0_1[90]}), .c ({y0_s1[90], y0_s0[90]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_91_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10879, mcs_out[219]}), .a ({new_AGEMA_signal_10985, y0_1[91]}), .c ({y0_s1[91], y0_s0[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_92_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10871, mcs_out[220]}), .a ({new_AGEMA_signal_10986, y0_1[92]}), .c ({y0_s1[92], y0_s0[92]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_93_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10870, mcs_out[221]}), .a ({new_AGEMA_signal_10987, y0_1[93]}), .c ({y0_s1[93], y0_s0[93]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_94_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10869, mcs_out[222]}), .a ({new_AGEMA_signal_10988, y0_1[94]}), .c ({y0_s1[94], y0_s0[94]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_95_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10868, mcs_out[223]}), .a ({new_AGEMA_signal_10989, y0_1[95]}), .c ({y0_s1[95], y0_s0[95]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_96_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10735, mcs_out[224]}), .a ({new_AGEMA_signal_10791, y0_1[96]}), .c ({y0_s1[96], y0_s0[96]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_97_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10933, mcs_out[225]}), .a ({new_AGEMA_signal_10990, y0_1[97]}), .c ({y0_s1[97], y0_s0[97]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_98_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10244, mcs_out[226]}), .a ({new_AGEMA_signal_10294, y0_1[98]}), .c ({y0_s1[98], y0_s0[98]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_99_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10932, mcs_out[227]}), .a ({new_AGEMA_signal_10991, y0_1[99]}), .c ({y0_s1[99], y0_s0[99]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_100_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10459, mcs_out[228]}), .a ({new_AGEMA_signal_10514, y0_1[100]}), .c ({y0_s1[100], y0_s0[100]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_101_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10716, mcs_out[229]}), .a ({new_AGEMA_signal_10764, y0_1[101]}), .c ({y0_s1[101], y0_s0[101]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_102_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10924, mcs_out[230]}), .a ({new_AGEMA_signal_10957, y0_1[102]}), .c ({y0_s1[102], y0_s0[102]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_103_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10923, mcs_out[231]}), .a ({new_AGEMA_signal_10958, y0_1[103]}), .c ({y0_s1[103], y0_s0[103]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_104_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10915, mcs_out[232]}), .a ({new_AGEMA_signal_10959, y0_1[104]}), .c ({y0_s1[104], y0_s0[104]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_105_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10196, mcs_out[233]}), .a ({new_AGEMA_signal_10278, y0_1[105]}), .c ({y0_s1[105], y0_s0[105]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_106_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10434, mcs_out[234]}), .a ({new_AGEMA_signal_10515, y0_1[106]}), .c ({y0_s1[106], y0_s0[106]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_107_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10698, mcs_out[235]}), .a ({new_AGEMA_signal_10765, y0_1[107]}), .c ({y0_s1[107], y0_s0[107]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_108_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9731, mcs_out[236]}), .a ({new_AGEMA_signal_9838, y0_1[108]}), .c ({y0_s1[108], y0_s0[108]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_109_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9955, mcs_out[237]}), .a ({new_AGEMA_signal_10046, y0_1[109]}), .c ({y0_s1[109], y0_s0[109]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_110_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9954, mcs_out[238]}), .a ({new_AGEMA_signal_10047, y0_1[110]}), .c ({y0_s1[110], y0_s0[110]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_111_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9728, mcs_out[239]}), .a ({new_AGEMA_signal_9839, y0_1[111]}), .c ({y0_s1[111], y0_s0[111]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_112_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10666, mcs_out[240]}), .a ({new_AGEMA_signal_10767, y0_1[112]}), .c ({y0_s1[112], y0_s0[112]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_113_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10896, mcs_out[241]}), .a ({new_AGEMA_signal_10960, y0_1[113]}), .c ({y0_s1[113], y0_s0[113]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_114_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10145, mcs_out[242]}), .a ({new_AGEMA_signal_10279, y0_1[114]}), .c ({y0_s1[114], y0_s0[114]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_115_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10895, mcs_out[243]}), .a ({new_AGEMA_signal_10961, y0_1[115]}), .c ({y0_s1[115], y0_s0[115]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_116_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10364, mcs_out[244]}), .a ({new_AGEMA_signal_10516, y0_1[116]}), .c ({y0_s1[116], y0_s0[116]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_117_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10647, mcs_out[245]}), .a ({new_AGEMA_signal_10768, y0_1[117]}), .c ({y0_s1[117], y0_s0[117]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_118_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10887, mcs_out[246]}), .a ({new_AGEMA_signal_10962, y0_1[118]}), .c ({y0_s1[118], y0_s0[118]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_119_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10886, mcs_out[247]}), .a ({new_AGEMA_signal_10963, y0_1[119]}), .c ({y0_s1[119], y0_s0[119]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_120_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10878, mcs_out[248]}), .a ({new_AGEMA_signal_10965, y0_1[120]}), .c ({y0_s1[120], y0_s0[120]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_121_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10097, mcs_out[249]}), .a ({new_AGEMA_signal_10280, y0_1[121]}), .c ({y0_s1[121], y0_s0[121]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_122_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10339, mcs_out[250]}), .a ({new_AGEMA_signal_10517, y0_1[122]}), .c ({y0_s1[122], y0_s0[122]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_123_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10629, mcs_out[251]}), .a ({new_AGEMA_signal_10769, y0_1[123]}), .c ({y0_s1[123], y0_s0[123]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_124_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9622, mcs_out[252]}), .a ({new_AGEMA_signal_9840, y0_1[124]}), .c ({y0_s1[124], y0_s0[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_125_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9862, mcs_out[253]}), .a ({new_AGEMA_signal_10048, y0_1[125]}), .c ({y0_s1[125], y0_s0[125]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_126_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9861, mcs_out[254]}), .a ({new_AGEMA_signal_10049, y0_1[126]}), .c ({y0_s1[126], y0_s0[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_inst2_MUXInst_127_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9619, mcs_out[255]}), .a ({new_AGEMA_signal_9841, y0_1[127]}), .c ({y0_s1[127], y0_s0[127]}) ) ;

endmodule
