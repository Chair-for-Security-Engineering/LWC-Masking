/* modified netlist. Source: module arx_round in file ./test/arx_round.v */
/* clock gating is added to the circuit, the latency increased 10 time(s)  */

module arx_round_HPC2_ClockGating_d3 (round_constant, round, x_round_in_s0, y_round_in_s0, clk, y_round_in_s1, y_round_in_s2, y_round_in_s3, x_round_in_s1, x_round_in_s2, x_round_in_s3, Fresh, /*rst,*/ x_round_out_s0, y_round_out_s0, x_round_out_s1, x_round_out_s2, x_round_out_s3, y_round_out_s1, y_round_out_s2, y_round_out_s3/*, Synch*/);
    input [31:0] round_constant ;
    input [1:0] round ;
    input [31:0] x_round_in_s0 ;
    input [31:0] y_round_in_s0 ;
    input clk ;
    input [31:0] y_round_in_s1 ;
    input [31:0] y_round_in_s2 ;
    input [31:0] y_round_in_s3 ;
    input [31:0] x_round_in_s1 ;
    input [31:0] x_round_in_s2 ;
    input [31:0] x_round_in_s3 ;
    //input rst ;
    input [1535:0] Fresh ;
    output [31:0] x_round_out_s0 ;
    output [31:0] y_round_out_s0 ;
    output [31:0] x_round_out_s1 ;
    output [31:0] x_round_out_s2 ;
    output [31:0] x_round_out_s3 ;
    output [31:0] y_round_out_s1 ;
    output [31:0] y_round_out_s2 ;
    output [31:0] y_round_out_s3 ;
    //output Synch ;
    wire AdderIns_s2_gc_0_a1_t ;
    wire AdderIns_s2_bc_0_a1_t ;
    wire AdderIns_s2_bc_1_a1_t ;
    wire AdderIns_s2_bc_2_a1_t ;
    wire AdderIns_s2_bc_3_a1_t ;
    wire AdderIns_s2_bc_4_a1_t ;
    wire AdderIns_s2_bc_5_a1_t ;
    wire AdderIns_s2_bc_6_a1_t ;
    wire AdderIns_s2_bc_7_a1_t ;
    wire AdderIns_s2_bc_8_a1_t ;
    wire AdderIns_s2_bc_9_a1_t ;
    wire AdderIns_s2_bc_10_a1_t ;
    wire AdderIns_s2_bc_11_a1_t ;
    wire AdderIns_s2_bc_12_a1_t ;
    wire AdderIns_s2_bc_13_a1_t ;
    wire AdderIns_s2_bc_14_a1_t ;
    wire AdderIns_s2_bc_15_a1_t ;
    wire AdderIns_s2_bc_16_a1_t ;
    wire AdderIns_s2_bc_17_a1_t ;
    wire AdderIns_s2_bc_18_a1_t ;
    wire AdderIns_s2_bc_19_a1_t ;
    wire AdderIns_s2_bc_20_a1_t ;
    wire AdderIns_s2_bc_21_a1_t ;
    wire AdderIns_s2_bc_22_a1_t ;
    wire AdderIns_s2_bc_23_a1_t ;
    wire AdderIns_s2_bc_24_a1_t ;
    wire AdderIns_s2_bc_25_a1_t ;
    wire AdderIns_s2_bc_26_a1_t ;
    wire AdderIns_s2_bc_27_a1_t ;
    wire AdderIns_s2_bc_28_a1_t ;
    wire AdderIns_s2_bc_29_a1_t ;
    wire AdderIns_s3_gc_0_a1_t ;
    wire AdderIns_s3_gc_1_a1_t ;
    wire AdderIns_s3_bc_0_a1_t ;
    wire AdderIns_s3_bc_1_a1_t ;
    wire AdderIns_s3_bc_2_a1_t ;
    wire AdderIns_s3_bc_3_a1_t ;
    wire AdderIns_s3_bc_4_a1_t ;
    wire AdderIns_s3_bc_5_a1_t ;
    wire AdderIns_s3_bc_6_a1_t ;
    wire AdderIns_s3_bc_7_a1_t ;
    wire AdderIns_s3_bc_8_a1_t ;
    wire AdderIns_s3_bc_9_a1_t ;
    wire AdderIns_s3_bc_10_a1_t ;
    wire AdderIns_s3_bc_11_a1_t ;
    wire AdderIns_s3_bc_12_a1_t ;
    wire AdderIns_s3_bc_13_a1_t ;
    wire AdderIns_s3_bc_14_a1_t ;
    wire AdderIns_s3_bc_15_a1_t ;
    wire AdderIns_s3_bc_16_a1_t ;
    wire AdderIns_s3_bc_17_a1_t ;
    wire AdderIns_s3_bc_18_a1_t ;
    wire AdderIns_s3_bc_19_a1_t ;
    wire AdderIns_s3_bc_20_a1_t ;
    wire AdderIns_s3_bc_21_a1_t ;
    wire AdderIns_s3_bc_22_a1_t ;
    wire AdderIns_s3_bc_23_a1_t ;
    wire AdderIns_s3_bc_24_a1_t ;
    wire AdderIns_s3_bc_25_a1_t ;
    wire AdderIns_s3_bc_26_a1_t ;
    wire AdderIns_s3_bc_27_a1_t ;
    wire AdderIns_s4_gc_0_a1_t ;
    wire AdderIns_s4_gc_1_a1_t ;
    wire AdderIns_s4_gc_2_a1_t ;
    wire AdderIns_s4_gc_3_a1_t ;
    wire AdderIns_s4_bc_0_a1_t ;
    wire AdderIns_s4_bc_1_a1_t ;
    wire AdderIns_s4_bc_2_a1_t ;
    wire AdderIns_s4_bc_3_a1_t ;
    wire AdderIns_s4_bc_4_a1_t ;
    wire AdderIns_s4_bc_5_a1_t ;
    wire AdderIns_s4_bc_6_a1_t ;
    wire AdderIns_s4_bc_7_a1_t ;
    wire AdderIns_s4_bc_8_a1_t ;
    wire AdderIns_s4_bc_9_a1_t ;
    wire AdderIns_s4_bc_10_a1_t ;
    wire AdderIns_s4_bc_11_a1_t ;
    wire AdderIns_s4_bc_12_a1_t ;
    wire AdderIns_s4_bc_13_a1_t ;
    wire AdderIns_s4_bc_14_a1_t ;
    wire AdderIns_s4_bc_15_a1_t ;
    wire AdderIns_s4_bc_16_a1_t ;
    wire AdderIns_s4_bc_17_a1_t ;
    wire AdderIns_s4_bc_18_a1_t ;
    wire AdderIns_s4_bc_19_a1_t ;
    wire AdderIns_s4_bc_20_a1_t ;
    wire AdderIns_s4_bc_21_a1_t ;
    wire AdderIns_s4_bc_22_a1_t ;
    wire AdderIns_s4_bc_23_a1_t ;
    wire AdderIns_s5_gc_0_a1_t ;
    wire AdderIns_s5_gc_1_a1_t ;
    wire AdderIns_s5_gc_2_a1_t ;
    wire AdderIns_s5_gc_3_a1_t ;
    wire AdderIns_s5_gc_4_a1_t ;
    wire AdderIns_s5_gc_5_a1_t ;
    wire AdderIns_s5_gc_6_a1_t ;
    wire AdderIns_s5_gc_7_a1_t ;
    wire AdderIns_s5_bc_0_a1_t ;
    wire AdderIns_s5_bc_1_a1_t ;
    wire AdderIns_s5_bc_2_a1_t ;
    wire AdderIns_s5_bc_3_a1_t ;
    wire AdderIns_s5_bc_4_a1_t ;
    wire AdderIns_s5_bc_5_a1_t ;
    wire AdderIns_s5_bc_6_a1_t ;
    wire AdderIns_s5_bc_7_a1_t ;
    wire AdderIns_s5_bc_8_a1_t ;
    wire AdderIns_s5_bc_9_a1_t ;
    wire AdderIns_s5_bc_10_a1_t ;
    wire AdderIns_s5_bc_11_a1_t ;
    wire AdderIns_s5_bc_12_a1_t ;
    wire AdderIns_s5_bc_13_a1_t ;
    wire AdderIns_s5_bc_14_a1_t ;
    wire AdderIns_s5_bc_15_a1_t ;
    wire AdderIns_s6_gc_1_a1_t ;
    wire AdderIns_s6_gc_2_a1_t ;
    wire AdderIns_s6_gc_3_a1_t ;
    wire AdderIns_s6_gc_4_a1_t ;
    wire AdderIns_s6_gc_5_a1_t ;
    wire AdderIns_s6_gc_6_a1_t ;
    wire AdderIns_s6_gc_7_a1_t ;
    wire AdderIns_s6_gc_8_a1_t ;
    wire AdderIns_s6_gc_9_a1_t ;
    wire AdderIns_s6_gc_10_a1_t ;
    wire AdderIns_s6_gc_11_a1_t ;
    wire AdderIns_s6_gc_12_a1_t ;
    wire AdderIns_s6_gc_13_a1_t ;
    wire AdderIns_s6_gc_14_a1_t ;
    wire AdderIns_s6_gc_15_a1_t ;
    wire [31:0] y_rotated01 ;
    wire [31:0] y_rotated23 ;
    wire [31:0] y_rotated ;
    wire [31:0] sum ;
    wire [31:0] sum_rotated01 ;
    wire [31:0] sum_rotated23 ;
    wire [31:0] sum_rotated ;
    wire [30:0] AdderIns_g6 ;
    wire [31:1] AdderIns_p6 ;
    wire [30:16] AdderIns_g5 ;
    wire [15:1] AdderIns_p5 ;
    wire [30:7] AdderIns_g4 ;
    wire [23:0] AdderIns_p4 ;
    wire [30:3] AdderIns_g3 ;
    wire [27:0] AdderIns_p3 ;
    wire [30:1] AdderIns_g2 ;
    wire [29:0] AdderIns_p2 ;
    wire [30:0] AdderIns_g1 ;
    wire new_AGEMA_signal_830 ;
    wire new_AGEMA_signal_831 ;
    wire new_AGEMA_signal_832 ;
    wire new_AGEMA_signal_839 ;
    wire new_AGEMA_signal_840 ;
    wire new_AGEMA_signal_841 ;
    wire new_AGEMA_signal_848 ;
    wire new_AGEMA_signal_849 ;
    wire new_AGEMA_signal_850 ;
    wire new_AGEMA_signal_857 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_859 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_868 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_886 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_902 ;
    wire new_AGEMA_signal_903 ;
    wire new_AGEMA_signal_904 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_912 ;
    wire new_AGEMA_signal_913 ;
    wire new_AGEMA_signal_920 ;
    wire new_AGEMA_signal_921 ;
    wire new_AGEMA_signal_922 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_930 ;
    wire new_AGEMA_signal_931 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_939 ;
    wire new_AGEMA_signal_940 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) U129 ( .a ({1'b0, 1'b0, 1'b0, round_constant[0]}), .b ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, new_AGEMA_signal_1211, sum[0]}), .c ({x_round_out_s3[0], x_round_out_s2[0], x_round_out_s1[0], x_round_out_s0[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_0_U1 ( .s (round[0]), .b ({y_round_in_s3[31], y_round_in_s2[31], y_round_in_s1[31], y_round_in_s0[31]}), .a ({y_round_in_s3[17], y_round_in_s2[17], y_round_in_s1[17], y_round_in_s0[17]}), .c ({new_AGEMA_signal_832, new_AGEMA_signal_831, new_AGEMA_signal_830, y_rotated01[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_1_U1 ( .s (round[0]), .b ({y_round_in_s3[0], y_round_in_s2[0], y_round_in_s1[0], y_round_in_s0[0]}), .a ({y_round_in_s3[18], y_round_in_s2[18], y_round_in_s1[18], y_round_in_s0[18]}), .c ({new_AGEMA_signal_841, new_AGEMA_signal_840, new_AGEMA_signal_839, y_rotated01[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_2_U1 ( .s (round[0]), .b ({y_round_in_s3[1], y_round_in_s2[1], y_round_in_s1[1], y_round_in_s0[1]}), .a ({y_round_in_s3[19], y_round_in_s2[19], y_round_in_s1[19], y_round_in_s0[19]}), .c ({new_AGEMA_signal_850, new_AGEMA_signal_849, new_AGEMA_signal_848, y_rotated01[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_3_U1 ( .s (round[0]), .b ({y_round_in_s3[2], y_round_in_s2[2], y_round_in_s1[2], y_round_in_s0[2]}), .a ({y_round_in_s3[20], y_round_in_s2[20], y_round_in_s1[20], y_round_in_s0[20]}), .c ({new_AGEMA_signal_859, new_AGEMA_signal_858, new_AGEMA_signal_857, y_rotated01[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_4_U1 ( .s (round[0]), .b ({y_round_in_s3[3], y_round_in_s2[3], y_round_in_s1[3], y_round_in_s0[3]}), .a ({y_round_in_s3[21], y_round_in_s2[21], y_round_in_s1[21], y_round_in_s0[21]}), .c ({new_AGEMA_signal_868, new_AGEMA_signal_867, new_AGEMA_signal_866, y_rotated01[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_5_U1 ( .s (round[0]), .b ({y_round_in_s3[4], y_round_in_s2[4], y_round_in_s1[4], y_round_in_s0[4]}), .a ({y_round_in_s3[22], y_round_in_s2[22], y_round_in_s1[22], y_round_in_s0[22]}), .c ({new_AGEMA_signal_877, new_AGEMA_signal_876, new_AGEMA_signal_875, y_rotated01[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_6_U1 ( .s (round[0]), .b ({y_round_in_s3[5], y_round_in_s2[5], y_round_in_s1[5], y_round_in_s0[5]}), .a ({y_round_in_s3[23], y_round_in_s2[23], y_round_in_s1[23], y_round_in_s0[23]}), .c ({new_AGEMA_signal_886, new_AGEMA_signal_885, new_AGEMA_signal_884, y_rotated01[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_7_U1 ( .s (round[0]), .b ({y_round_in_s3[6], y_round_in_s2[6], y_round_in_s1[6], y_round_in_s0[6]}), .a ({y_round_in_s3[24], y_round_in_s2[24], y_round_in_s1[24], y_round_in_s0[24]}), .c ({new_AGEMA_signal_895, new_AGEMA_signal_894, new_AGEMA_signal_893, y_rotated01[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_8_U1 ( .s (round[0]), .b ({y_round_in_s3[7], y_round_in_s2[7], y_round_in_s1[7], y_round_in_s0[7]}), .a ({y_round_in_s3[25], y_round_in_s2[25], y_round_in_s1[25], y_round_in_s0[25]}), .c ({new_AGEMA_signal_904, new_AGEMA_signal_903, new_AGEMA_signal_902, y_rotated01[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_9_U1 ( .s (round[0]), .b ({y_round_in_s3[8], y_round_in_s2[8], y_round_in_s1[8], y_round_in_s0[8]}), .a ({y_round_in_s3[26], y_round_in_s2[26], y_round_in_s1[26], y_round_in_s0[26]}), .c ({new_AGEMA_signal_913, new_AGEMA_signal_912, new_AGEMA_signal_911, y_rotated01[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_10_U1 ( .s (round[0]), .b ({y_round_in_s3[9], y_round_in_s2[9], y_round_in_s1[9], y_round_in_s0[9]}), .a ({y_round_in_s3[27], y_round_in_s2[27], y_round_in_s1[27], y_round_in_s0[27]}), .c ({new_AGEMA_signal_922, new_AGEMA_signal_921, new_AGEMA_signal_920, y_rotated01[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_11_U1 ( .s (round[0]), .b ({y_round_in_s3[10], y_round_in_s2[10], y_round_in_s1[10], y_round_in_s0[10]}), .a ({y_round_in_s3[28], y_round_in_s2[28], y_round_in_s1[28], y_round_in_s0[28]}), .c ({new_AGEMA_signal_931, new_AGEMA_signal_930, new_AGEMA_signal_929, y_rotated01[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_12_U1 ( .s (round[0]), .b ({y_round_in_s3[11], y_round_in_s2[11], y_round_in_s1[11], y_round_in_s0[11]}), .a ({y_round_in_s3[29], y_round_in_s2[29], y_round_in_s1[29], y_round_in_s0[29]}), .c ({new_AGEMA_signal_940, new_AGEMA_signal_939, new_AGEMA_signal_938, y_rotated01[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_13_U1 ( .s (round[0]), .b ({y_round_in_s3[12], y_round_in_s2[12], y_round_in_s1[12], y_round_in_s0[12]}), .a ({y_round_in_s3[30], y_round_in_s2[30], y_round_in_s1[30], y_round_in_s0[30]}), .c ({new_AGEMA_signal_949, new_AGEMA_signal_948, new_AGEMA_signal_947, y_rotated01[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_14_U1 ( .s (round[0]), .b ({y_round_in_s3[13], y_round_in_s2[13], y_round_in_s1[13], y_round_in_s0[13]}), .a ({y_round_in_s3[31], y_round_in_s2[31], y_round_in_s1[31], y_round_in_s0[31]}), .c ({new_AGEMA_signal_955, new_AGEMA_signal_954, new_AGEMA_signal_953, y_rotated01[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_15_U1 ( .s (round[0]), .b ({y_round_in_s3[14], y_round_in_s2[14], y_round_in_s1[14], y_round_in_s0[14]}), .a ({y_round_in_s3[0], y_round_in_s2[0], y_round_in_s1[0], y_round_in_s0[0]}), .c ({new_AGEMA_signal_961, new_AGEMA_signal_960, new_AGEMA_signal_959, y_rotated01[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_16_U1 ( .s (round[0]), .b ({y_round_in_s3[15], y_round_in_s2[15], y_round_in_s1[15], y_round_in_s0[15]}), .a ({y_round_in_s3[1], y_round_in_s2[1], y_round_in_s1[1], y_round_in_s0[1]}), .c ({new_AGEMA_signal_967, new_AGEMA_signal_966, new_AGEMA_signal_965, y_rotated01[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_17_U1 ( .s (round[0]), .b ({y_round_in_s3[16], y_round_in_s2[16], y_round_in_s1[16], y_round_in_s0[16]}), .a ({y_round_in_s3[2], y_round_in_s2[2], y_round_in_s1[2], y_round_in_s0[2]}), .c ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, y_rotated01[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_18_U1 ( .s (round[0]), .b ({y_round_in_s3[17], y_round_in_s2[17], y_round_in_s1[17], y_round_in_s0[17]}), .a ({y_round_in_s3[3], y_round_in_s2[3], y_round_in_s1[3], y_round_in_s0[3]}), .c ({new_AGEMA_signal_976, new_AGEMA_signal_975, new_AGEMA_signal_974, y_rotated01[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_19_U1 ( .s (round[0]), .b ({y_round_in_s3[18], y_round_in_s2[18], y_round_in_s1[18], y_round_in_s0[18]}), .a ({y_round_in_s3[4], y_round_in_s2[4], y_round_in_s1[4], y_round_in_s0[4]}), .c ({new_AGEMA_signal_979, new_AGEMA_signal_978, new_AGEMA_signal_977, y_rotated01[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_20_U1 ( .s (round[0]), .b ({y_round_in_s3[19], y_round_in_s2[19], y_round_in_s1[19], y_round_in_s0[19]}), .a ({y_round_in_s3[5], y_round_in_s2[5], y_round_in_s1[5], y_round_in_s0[5]}), .c ({new_AGEMA_signal_982, new_AGEMA_signal_981, new_AGEMA_signal_980, y_rotated01[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_21_U1 ( .s (round[0]), .b ({y_round_in_s3[20], y_round_in_s2[20], y_round_in_s1[20], y_round_in_s0[20]}), .a ({y_round_in_s3[6], y_round_in_s2[6], y_round_in_s1[6], y_round_in_s0[6]}), .c ({new_AGEMA_signal_985, new_AGEMA_signal_984, new_AGEMA_signal_983, y_rotated01[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_22_U1 ( .s (round[0]), .b ({y_round_in_s3[21], y_round_in_s2[21], y_round_in_s1[21], y_round_in_s0[21]}), .a ({y_round_in_s3[7], y_round_in_s2[7], y_round_in_s1[7], y_round_in_s0[7]}), .c ({new_AGEMA_signal_988, new_AGEMA_signal_987, new_AGEMA_signal_986, y_rotated01[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_23_U1 ( .s (round[0]), .b ({y_round_in_s3[22], y_round_in_s2[22], y_round_in_s1[22], y_round_in_s0[22]}), .a ({y_round_in_s3[8], y_round_in_s2[8], y_round_in_s1[8], y_round_in_s0[8]}), .c ({new_AGEMA_signal_991, new_AGEMA_signal_990, new_AGEMA_signal_989, y_rotated01[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_24_U1 ( .s (round[0]), .b ({y_round_in_s3[23], y_round_in_s2[23], y_round_in_s1[23], y_round_in_s0[23]}), .a ({y_round_in_s3[9], y_round_in_s2[9], y_round_in_s1[9], y_round_in_s0[9]}), .c ({new_AGEMA_signal_994, new_AGEMA_signal_993, new_AGEMA_signal_992, y_rotated01[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_25_U1 ( .s (round[0]), .b ({y_round_in_s3[24], y_round_in_s2[24], y_round_in_s1[24], y_round_in_s0[24]}), .a ({y_round_in_s3[10], y_round_in_s2[10], y_round_in_s1[10], y_round_in_s0[10]}), .c ({new_AGEMA_signal_997, new_AGEMA_signal_996, new_AGEMA_signal_995, y_rotated01[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_26_U1 ( .s (round[0]), .b ({y_round_in_s3[25], y_round_in_s2[25], y_round_in_s1[25], y_round_in_s0[25]}), .a ({y_round_in_s3[11], y_round_in_s2[11], y_round_in_s1[11], y_round_in_s0[11]}), .c ({new_AGEMA_signal_1000, new_AGEMA_signal_999, new_AGEMA_signal_998, y_rotated01[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_27_U1 ( .s (round[0]), .b ({y_round_in_s3[26], y_round_in_s2[26], y_round_in_s1[26], y_round_in_s0[26]}), .a ({y_round_in_s3[12], y_round_in_s2[12], y_round_in_s1[12], y_round_in_s0[12]}), .c ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, new_AGEMA_signal_1001, y_rotated01[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_28_U1 ( .s (round[0]), .b ({y_round_in_s3[27], y_round_in_s2[27], y_round_in_s1[27], y_round_in_s0[27]}), .a ({y_round_in_s3[13], y_round_in_s2[13], y_round_in_s1[13], y_round_in_s0[13]}), .c ({new_AGEMA_signal_1006, new_AGEMA_signal_1005, new_AGEMA_signal_1004, y_rotated01[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_29_U1 ( .s (round[0]), .b ({y_round_in_s3[28], y_round_in_s2[28], y_round_in_s1[28], y_round_in_s0[28]}), .a ({y_round_in_s3[14], y_round_in_s2[14], y_round_in_s1[14], y_round_in_s0[14]}), .c ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, new_AGEMA_signal_1007, y_rotated01[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_30_U1 ( .s (round[0]), .b ({y_round_in_s3[29], y_round_in_s2[29], y_round_in_s1[29], y_round_in_s0[29]}), .a ({y_round_in_s3[15], y_round_in_s2[15], y_round_in_s1[15], y_round_in_s0[15]}), .c ({new_AGEMA_signal_1012, new_AGEMA_signal_1011, new_AGEMA_signal_1010, y_rotated01[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M0_mux_inst_31_U1 ( .s (round[0]), .b ({y_round_in_s3[30], y_round_in_s2[30], y_round_in_s1[30], y_round_in_s0[30]}), .a ({y_round_in_s3[16], y_round_in_s2[16], y_round_in_s1[16], y_round_in_s0[16]}), .c ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, new_AGEMA_signal_1013, y_rotated01[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_0_U1 ( .s (round[0]), .b ({y_round_in_s3[0], y_round_in_s2[0], y_round_in_s1[0], y_round_in_s0[0]}), .a ({y_round_in_s3[24], y_round_in_s2[24], y_round_in_s1[24], y_round_in_s0[24]}), .c ({new_AGEMA_signal_1018, new_AGEMA_signal_1017, new_AGEMA_signal_1016, y_rotated23[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_1_U1 ( .s (round[0]), .b ({y_round_in_s3[1], y_round_in_s2[1], y_round_in_s1[1], y_round_in_s0[1]}), .a ({y_round_in_s3[25], y_round_in_s2[25], y_round_in_s1[25], y_round_in_s0[25]}), .c ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, y_rotated23[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_2_U1 ( .s (round[0]), .b ({y_round_in_s3[2], y_round_in_s2[2], y_round_in_s1[2], y_round_in_s0[2]}), .a ({y_round_in_s3[26], y_round_in_s2[26], y_round_in_s1[26], y_round_in_s0[26]}), .c ({new_AGEMA_signal_1024, new_AGEMA_signal_1023, new_AGEMA_signal_1022, y_rotated23[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_3_U1 ( .s (round[0]), .b ({y_round_in_s3[3], y_round_in_s2[3], y_round_in_s1[3], y_round_in_s0[3]}), .a ({y_round_in_s3[27], y_round_in_s2[27], y_round_in_s1[27], y_round_in_s0[27]}), .c ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, new_AGEMA_signal_1025, y_rotated23[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_4_U1 ( .s (round[0]), .b ({y_round_in_s3[4], y_round_in_s2[4], y_round_in_s1[4], y_round_in_s0[4]}), .a ({y_round_in_s3[28], y_round_in_s2[28], y_round_in_s1[28], y_round_in_s0[28]}), .c ({new_AGEMA_signal_1030, new_AGEMA_signal_1029, new_AGEMA_signal_1028, y_rotated23[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_5_U1 ( .s (round[0]), .b ({y_round_in_s3[5], y_round_in_s2[5], y_round_in_s1[5], y_round_in_s0[5]}), .a ({y_round_in_s3[29], y_round_in_s2[29], y_round_in_s1[29], y_round_in_s0[29]}), .c ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, y_rotated23[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_6_U1 ( .s (round[0]), .b ({y_round_in_s3[6], y_round_in_s2[6], y_round_in_s1[6], y_round_in_s0[6]}), .a ({y_round_in_s3[30], y_round_in_s2[30], y_round_in_s1[30], y_round_in_s0[30]}), .c ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, y_rotated23[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_7_U1 ( .s (round[0]), .b ({y_round_in_s3[7], y_round_in_s2[7], y_round_in_s1[7], y_round_in_s0[7]}), .a ({y_round_in_s3[31], y_round_in_s2[31], y_round_in_s1[31], y_round_in_s0[31]}), .c ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, new_AGEMA_signal_1037, y_rotated23[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_8_U1 ( .s (round[0]), .b ({y_round_in_s3[8], y_round_in_s2[8], y_round_in_s1[8], y_round_in_s0[8]}), .a ({y_round_in_s3[0], y_round_in_s2[0], y_round_in_s1[0], y_round_in_s0[0]}), .c ({new_AGEMA_signal_1042, new_AGEMA_signal_1041, new_AGEMA_signal_1040, y_rotated23[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_9_U1 ( .s (round[0]), .b ({y_round_in_s3[9], y_round_in_s2[9], y_round_in_s1[9], y_round_in_s0[9]}), .a ({y_round_in_s3[1], y_round_in_s2[1], y_round_in_s1[1], y_round_in_s0[1]}), .c ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, new_AGEMA_signal_1043, y_rotated23[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_10_U1 ( .s (round[0]), .b ({y_round_in_s3[10], y_round_in_s2[10], y_round_in_s1[10], y_round_in_s0[10]}), .a ({y_round_in_s3[2], y_round_in_s2[2], y_round_in_s1[2], y_round_in_s0[2]}), .c ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, new_AGEMA_signal_1046, y_rotated23[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_11_U1 ( .s (round[0]), .b ({y_round_in_s3[11], y_round_in_s2[11], y_round_in_s1[11], y_round_in_s0[11]}), .a ({y_round_in_s3[3], y_round_in_s2[3], y_round_in_s1[3], y_round_in_s0[3]}), .c ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, new_AGEMA_signal_1049, y_rotated23[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_12_U1 ( .s (round[0]), .b ({y_round_in_s3[12], y_round_in_s2[12], y_round_in_s1[12], y_round_in_s0[12]}), .a ({y_round_in_s3[4], y_round_in_s2[4], y_round_in_s1[4], y_round_in_s0[4]}), .c ({new_AGEMA_signal_1054, new_AGEMA_signal_1053, new_AGEMA_signal_1052, y_rotated23[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_13_U1 ( .s (round[0]), .b ({y_round_in_s3[13], y_round_in_s2[13], y_round_in_s1[13], y_round_in_s0[13]}), .a ({y_round_in_s3[5], y_round_in_s2[5], y_round_in_s1[5], y_round_in_s0[5]}), .c ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, y_rotated23[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_14_U1 ( .s (round[0]), .b ({y_round_in_s3[14], y_round_in_s2[14], y_round_in_s1[14], y_round_in_s0[14]}), .a ({y_round_in_s3[6], y_round_in_s2[6], y_round_in_s1[6], y_round_in_s0[6]}), .c ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, y_rotated23[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_15_U1 ( .s (round[0]), .b ({y_round_in_s3[15], y_round_in_s2[15], y_round_in_s1[15], y_round_in_s0[15]}), .a ({y_round_in_s3[7], y_round_in_s2[7], y_round_in_s1[7], y_round_in_s0[7]}), .c ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, new_AGEMA_signal_1061, y_rotated23[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_16_U1 ( .s (round[0]), .b ({y_round_in_s3[16], y_round_in_s2[16], y_round_in_s1[16], y_round_in_s0[16]}), .a ({y_round_in_s3[8], y_round_in_s2[8], y_round_in_s1[8], y_round_in_s0[8]}), .c ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, new_AGEMA_signal_1064, y_rotated23[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_17_U1 ( .s (round[0]), .b ({y_round_in_s3[17], y_round_in_s2[17], y_round_in_s1[17], y_round_in_s0[17]}), .a ({y_round_in_s3[9], y_round_in_s2[9], y_round_in_s1[9], y_round_in_s0[9]}), .c ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, new_AGEMA_signal_1067, y_rotated23[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_18_U1 ( .s (round[0]), .b ({y_round_in_s3[18], y_round_in_s2[18], y_round_in_s1[18], y_round_in_s0[18]}), .a ({y_round_in_s3[10], y_round_in_s2[10], y_round_in_s1[10], y_round_in_s0[10]}), .c ({new_AGEMA_signal_1072, new_AGEMA_signal_1071, new_AGEMA_signal_1070, y_rotated23[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_19_U1 ( .s (round[0]), .b ({y_round_in_s3[19], y_round_in_s2[19], y_round_in_s1[19], y_round_in_s0[19]}), .a ({y_round_in_s3[11], y_round_in_s2[11], y_round_in_s1[11], y_round_in_s0[11]}), .c ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, new_AGEMA_signal_1073, y_rotated23[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_20_U1 ( .s (round[0]), .b ({y_round_in_s3[20], y_round_in_s2[20], y_round_in_s1[20], y_round_in_s0[20]}), .a ({y_round_in_s3[12], y_round_in_s2[12], y_round_in_s1[12], y_round_in_s0[12]}), .c ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, new_AGEMA_signal_1076, y_rotated23[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_21_U1 ( .s (round[0]), .b ({y_round_in_s3[21], y_round_in_s2[21], y_round_in_s1[21], y_round_in_s0[21]}), .a ({y_round_in_s3[13], y_round_in_s2[13], y_round_in_s1[13], y_round_in_s0[13]}), .c ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, y_rotated23[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_22_U1 ( .s (round[0]), .b ({y_round_in_s3[22], y_round_in_s2[22], y_round_in_s1[22], y_round_in_s0[22]}), .a ({y_round_in_s3[14], y_round_in_s2[14], y_round_in_s1[14], y_round_in_s0[14]}), .c ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, new_AGEMA_signal_1082, y_rotated23[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_23_U1 ( .s (round[0]), .b ({y_round_in_s3[23], y_round_in_s2[23], y_round_in_s1[23], y_round_in_s0[23]}), .a ({y_round_in_s3[15], y_round_in_s2[15], y_round_in_s1[15], y_round_in_s0[15]}), .c ({new_AGEMA_signal_1087, new_AGEMA_signal_1086, new_AGEMA_signal_1085, y_rotated23[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_24_U1 ( .s (round[0]), .b ({y_round_in_s3[24], y_round_in_s2[24], y_round_in_s1[24], y_round_in_s0[24]}), .a ({y_round_in_s3[16], y_round_in_s2[16], y_round_in_s1[16], y_round_in_s0[16]}), .c ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, new_AGEMA_signal_1088, y_rotated23[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_25_U1 ( .s (round[0]), .b ({y_round_in_s3[25], y_round_in_s2[25], y_round_in_s1[25], y_round_in_s0[25]}), .a ({y_round_in_s3[17], y_round_in_s2[17], y_round_in_s1[17], y_round_in_s0[17]}), .c ({new_AGEMA_signal_1093, new_AGEMA_signal_1092, new_AGEMA_signal_1091, y_rotated23[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_26_U1 ( .s (round[0]), .b ({y_round_in_s3[26], y_round_in_s2[26], y_round_in_s1[26], y_round_in_s0[26]}), .a ({y_round_in_s3[18], y_round_in_s2[18], y_round_in_s1[18], y_round_in_s0[18]}), .c ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, new_AGEMA_signal_1094, y_rotated23[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_27_U1 ( .s (round[0]), .b ({y_round_in_s3[27], y_round_in_s2[27], y_round_in_s1[27], y_round_in_s0[27]}), .a ({y_round_in_s3[19], y_round_in_s2[19], y_round_in_s1[19], y_round_in_s0[19]}), .c ({new_AGEMA_signal_1099, new_AGEMA_signal_1098, new_AGEMA_signal_1097, y_rotated23[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_28_U1 ( .s (round[0]), .b ({y_round_in_s3[28], y_round_in_s2[28], y_round_in_s1[28], y_round_in_s0[28]}), .a ({y_round_in_s3[20], y_round_in_s2[20], y_round_in_s1[20], y_round_in_s0[20]}), .c ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, new_AGEMA_signal_1100, y_rotated23[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_29_U1 ( .s (round[0]), .b ({y_round_in_s3[29], y_round_in_s2[29], y_round_in_s1[29], y_round_in_s0[29]}), .a ({y_round_in_s3[21], y_round_in_s2[21], y_round_in_s1[21], y_round_in_s0[21]}), .c ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, y_rotated23[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_30_U1 ( .s (round[0]), .b ({y_round_in_s3[30], y_round_in_s2[30], y_round_in_s1[30], y_round_in_s0[30]}), .a ({y_round_in_s3[22], y_round_in_s2[22], y_round_in_s1[22], y_round_in_s0[22]}), .c ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, y_rotated23[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M1_mux_inst_31_U1 ( .s (round[0]), .b ({y_round_in_s3[31], y_round_in_s2[31], y_round_in_s1[31], y_round_in_s0[31]}), .a ({y_round_in_s3[23], y_round_in_s2[23], y_round_in_s1[23], y_round_in_s0[23]}), .c ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, new_AGEMA_signal_1109, y_rotated23[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_0_U1 ( .s (round[1]), .b ({new_AGEMA_signal_832, new_AGEMA_signal_831, new_AGEMA_signal_830, y_rotated01[0]}), .a ({new_AGEMA_signal_1018, new_AGEMA_signal_1017, new_AGEMA_signal_1016, y_rotated23[0]}), .c ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, new_AGEMA_signal_1112, y_rotated[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_1_U1 ( .s (round[1]), .b ({new_AGEMA_signal_841, new_AGEMA_signal_840, new_AGEMA_signal_839, y_rotated01[1]}), .a ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, new_AGEMA_signal_1019, y_rotated23[1]}), .c ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, new_AGEMA_signal_1115, y_rotated[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_2_U1 ( .s (round[1]), .b ({new_AGEMA_signal_850, new_AGEMA_signal_849, new_AGEMA_signal_848, y_rotated01[2]}), .a ({new_AGEMA_signal_1024, new_AGEMA_signal_1023, new_AGEMA_signal_1022, y_rotated23[2]}), .c ({new_AGEMA_signal_1120, new_AGEMA_signal_1119, new_AGEMA_signal_1118, y_rotated[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_3_U1 ( .s (round[1]), .b ({new_AGEMA_signal_859, new_AGEMA_signal_858, new_AGEMA_signal_857, y_rotated01[3]}), .a ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, new_AGEMA_signal_1025, y_rotated23[3]}), .c ({new_AGEMA_signal_1123, new_AGEMA_signal_1122, new_AGEMA_signal_1121, y_rotated[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_4_U1 ( .s (round[1]), .b ({new_AGEMA_signal_868, new_AGEMA_signal_867, new_AGEMA_signal_866, y_rotated01[4]}), .a ({new_AGEMA_signal_1030, new_AGEMA_signal_1029, new_AGEMA_signal_1028, y_rotated23[4]}), .c ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, new_AGEMA_signal_1124, y_rotated[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_5_U1 ( .s (round[1]), .b ({new_AGEMA_signal_877, new_AGEMA_signal_876, new_AGEMA_signal_875, y_rotated01[5]}), .a ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, y_rotated23[5]}), .c ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, new_AGEMA_signal_1127, y_rotated[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_6_U1 ( .s (round[1]), .b ({new_AGEMA_signal_886, new_AGEMA_signal_885, new_AGEMA_signal_884, y_rotated01[6]}), .a ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, y_rotated23[6]}), .c ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, new_AGEMA_signal_1130, y_rotated[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_7_U1 ( .s (round[1]), .b ({new_AGEMA_signal_895, new_AGEMA_signal_894, new_AGEMA_signal_893, y_rotated01[7]}), .a ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, new_AGEMA_signal_1037, y_rotated23[7]}), .c ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, new_AGEMA_signal_1133, y_rotated[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_8_U1 ( .s (round[1]), .b ({new_AGEMA_signal_904, new_AGEMA_signal_903, new_AGEMA_signal_902, y_rotated01[8]}), .a ({new_AGEMA_signal_1042, new_AGEMA_signal_1041, new_AGEMA_signal_1040, y_rotated23[8]}), .c ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, new_AGEMA_signal_1136, y_rotated[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_9_U1 ( .s (round[1]), .b ({new_AGEMA_signal_913, new_AGEMA_signal_912, new_AGEMA_signal_911, y_rotated01[9]}), .a ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, new_AGEMA_signal_1043, y_rotated23[9]}), .c ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, new_AGEMA_signal_1139, y_rotated[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_10_U1 ( .s (round[1]), .b ({new_AGEMA_signal_922, new_AGEMA_signal_921, new_AGEMA_signal_920, y_rotated01[10]}), .a ({new_AGEMA_signal_1048, new_AGEMA_signal_1047, new_AGEMA_signal_1046, y_rotated23[10]}), .c ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, new_AGEMA_signal_1142, y_rotated[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_11_U1 ( .s (round[1]), .b ({new_AGEMA_signal_931, new_AGEMA_signal_930, new_AGEMA_signal_929, y_rotated01[11]}), .a ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, new_AGEMA_signal_1049, y_rotated23[11]}), .c ({new_AGEMA_signal_1147, new_AGEMA_signal_1146, new_AGEMA_signal_1145, y_rotated[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_12_U1 ( .s (round[1]), .b ({new_AGEMA_signal_940, new_AGEMA_signal_939, new_AGEMA_signal_938, y_rotated01[12]}), .a ({new_AGEMA_signal_1054, new_AGEMA_signal_1053, new_AGEMA_signal_1052, y_rotated23[12]}), .c ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, new_AGEMA_signal_1148, y_rotated[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_13_U1 ( .s (round[1]), .b ({new_AGEMA_signal_949, new_AGEMA_signal_948, new_AGEMA_signal_947, y_rotated01[13]}), .a ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, y_rotated23[13]}), .c ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, y_rotated[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_14_U1 ( .s (round[1]), .b ({new_AGEMA_signal_955, new_AGEMA_signal_954, new_AGEMA_signal_953, y_rotated01[14]}), .a ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, y_rotated23[14]}), .c ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, y_rotated[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_15_U1 ( .s (round[1]), .b ({new_AGEMA_signal_961, new_AGEMA_signal_960, new_AGEMA_signal_959, y_rotated01[15]}), .a ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, new_AGEMA_signal_1061, y_rotated23[15]}), .c ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, new_AGEMA_signal_1157, y_rotated[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_16_U1 ( .s (round[1]), .b ({new_AGEMA_signal_967, new_AGEMA_signal_966, new_AGEMA_signal_965, y_rotated01[16]}), .a ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, new_AGEMA_signal_1064, y_rotated23[16]}), .c ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, new_AGEMA_signal_1160, y_rotated[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_17_U1 ( .s (round[1]), .b ({new_AGEMA_signal_973, new_AGEMA_signal_972, new_AGEMA_signal_971, y_rotated01[17]}), .a ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, new_AGEMA_signal_1067, y_rotated23[17]}), .c ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, new_AGEMA_signal_1163, y_rotated[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_18_U1 ( .s (round[1]), .b ({new_AGEMA_signal_976, new_AGEMA_signal_975, new_AGEMA_signal_974, y_rotated01[18]}), .a ({new_AGEMA_signal_1072, new_AGEMA_signal_1071, new_AGEMA_signal_1070, y_rotated23[18]}), .c ({new_AGEMA_signal_1168, new_AGEMA_signal_1167, new_AGEMA_signal_1166, y_rotated[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_19_U1 ( .s (round[1]), .b ({new_AGEMA_signal_979, new_AGEMA_signal_978, new_AGEMA_signal_977, y_rotated01[19]}), .a ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, new_AGEMA_signal_1073, y_rotated23[19]}), .c ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, new_AGEMA_signal_1169, y_rotated[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_20_U1 ( .s (round[1]), .b ({new_AGEMA_signal_982, new_AGEMA_signal_981, new_AGEMA_signal_980, y_rotated01[20]}), .a ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, new_AGEMA_signal_1076, y_rotated23[20]}), .c ({new_AGEMA_signal_1174, new_AGEMA_signal_1173, new_AGEMA_signal_1172, y_rotated[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_21_U1 ( .s (round[1]), .b ({new_AGEMA_signal_985, new_AGEMA_signal_984, new_AGEMA_signal_983, y_rotated01[21]}), .a ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, y_rotated23[21]}), .c ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, new_AGEMA_signal_1175, y_rotated[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_22_U1 ( .s (round[1]), .b ({new_AGEMA_signal_988, new_AGEMA_signal_987, new_AGEMA_signal_986, y_rotated01[22]}), .a ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, new_AGEMA_signal_1082, y_rotated23[22]}), .c ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, y_rotated[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_23_U1 ( .s (round[1]), .b ({new_AGEMA_signal_991, new_AGEMA_signal_990, new_AGEMA_signal_989, y_rotated01[23]}), .a ({new_AGEMA_signal_1087, new_AGEMA_signal_1086, new_AGEMA_signal_1085, y_rotated23[23]}), .c ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, new_AGEMA_signal_1181, y_rotated[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_24_U1 ( .s (round[1]), .b ({new_AGEMA_signal_994, new_AGEMA_signal_993, new_AGEMA_signal_992, y_rotated01[24]}), .a ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, new_AGEMA_signal_1088, y_rotated23[24]}), .c ({new_AGEMA_signal_1186, new_AGEMA_signal_1185, new_AGEMA_signal_1184, y_rotated[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_25_U1 ( .s (round[1]), .b ({new_AGEMA_signal_997, new_AGEMA_signal_996, new_AGEMA_signal_995, y_rotated01[25]}), .a ({new_AGEMA_signal_1093, new_AGEMA_signal_1092, new_AGEMA_signal_1091, y_rotated23[25]}), .c ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, new_AGEMA_signal_1187, y_rotated[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_26_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1000, new_AGEMA_signal_999, new_AGEMA_signal_998, y_rotated01[26]}), .a ({new_AGEMA_signal_1096, new_AGEMA_signal_1095, new_AGEMA_signal_1094, y_rotated23[26]}), .c ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, new_AGEMA_signal_1190, y_rotated[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_27_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, new_AGEMA_signal_1001, y_rotated01[27]}), .a ({new_AGEMA_signal_1099, new_AGEMA_signal_1098, new_AGEMA_signal_1097, y_rotated23[27]}), .c ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, new_AGEMA_signal_1193, y_rotated[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_28_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1006, new_AGEMA_signal_1005, new_AGEMA_signal_1004, y_rotated01[28]}), .a ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, new_AGEMA_signal_1100, y_rotated23[28]}), .c ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, new_AGEMA_signal_1196, y_rotated[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_29_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, new_AGEMA_signal_1007, y_rotated01[29]}), .a ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, y_rotated23[29]}), .c ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, new_AGEMA_signal_1199, y_rotated[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_30_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1012, new_AGEMA_signal_1011, new_AGEMA_signal_1010, y_rotated01[30]}), .a ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, y_rotated23[30]}), .c ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, y_rotated[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M3_mux_inst_31_U1 ( .s (round[1]), .b ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, new_AGEMA_signal_1013, y_rotated01[31]}), .a ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, new_AGEMA_signal_1109, y_rotated23[31]}), .c ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, new_AGEMA_signal_1205, y_rotated[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_0_U1 ( .a ({x_round_in_s3[0], x_round_in_s2[0], x_round_in_s1[0], x_round_in_s0[0]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, new_AGEMA_signal_1112, y_rotated[0]}), .c ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, new_AGEMA_signal_1211, sum[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_1_U1 ( .a ({x_round_in_s3[1], x_round_in_s2[1], x_round_in_s1[1], x_round_in_s0[1]}), .b ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, new_AGEMA_signal_1115, y_rotated[1]}), .c ({new_AGEMA_signal_1222, new_AGEMA_signal_1221, new_AGEMA_signal_1220, AdderIns_p6[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_2_U1 ( .a ({x_round_in_s3[2], x_round_in_s2[2], x_round_in_s1[2], x_round_in_s0[2]}), .b ({new_AGEMA_signal_1120, new_AGEMA_signal_1119, new_AGEMA_signal_1118, y_rotated[2]}), .c ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, new_AGEMA_signal_1229, AdderIns_p6[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_3_U1 ( .a ({x_round_in_s3[3], x_round_in_s2[3], x_round_in_s1[3], x_round_in_s0[3]}), .b ({new_AGEMA_signal_1123, new_AGEMA_signal_1122, new_AGEMA_signal_1121, y_rotated[3]}), .c ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, new_AGEMA_signal_1238, AdderIns_p6[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_4_U1 ( .a ({x_round_in_s3[4], x_round_in_s2[4], x_round_in_s1[4], x_round_in_s0[4]}), .b ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, new_AGEMA_signal_1124, y_rotated[4]}), .c ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, new_AGEMA_signal_1247, AdderIns_p6[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_5_U1 ( .a ({x_round_in_s3[5], x_round_in_s2[5], x_round_in_s1[5], x_round_in_s0[5]}), .b ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, new_AGEMA_signal_1127, y_rotated[5]}), .c ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, new_AGEMA_signal_1256, AdderIns_p6[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_6_U1 ( .a ({x_round_in_s3[6], x_round_in_s2[6], x_round_in_s1[6], x_round_in_s0[6]}), .b ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, new_AGEMA_signal_1130, y_rotated[6]}), .c ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, new_AGEMA_signal_1265, AdderIns_p6[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_7_U1 ( .a ({x_round_in_s3[7], x_round_in_s2[7], x_round_in_s1[7], x_round_in_s0[7]}), .b ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, new_AGEMA_signal_1133, y_rotated[7]}), .c ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, AdderIns_p6[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_8_U1 ( .a ({x_round_in_s3[8], x_round_in_s2[8], x_round_in_s1[8], x_round_in_s0[8]}), .b ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, new_AGEMA_signal_1136, y_rotated[8]}), .c ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, AdderIns_p6[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_9_U1 ( .a ({x_round_in_s3[9], x_round_in_s2[9], x_round_in_s1[9], x_round_in_s0[9]}), .b ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, new_AGEMA_signal_1139, y_rotated[9]}), .c ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, new_AGEMA_signal_1292, AdderIns_p6[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_10_U1 ( .a ({x_round_in_s3[10], x_round_in_s2[10], x_round_in_s1[10], x_round_in_s0[10]}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, new_AGEMA_signal_1142, y_rotated[10]}), .c ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, new_AGEMA_signal_1301, AdderIns_p6[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_11_U1 ( .a ({x_round_in_s3[11], x_round_in_s2[11], x_round_in_s1[11], x_round_in_s0[11]}), .b ({new_AGEMA_signal_1147, new_AGEMA_signal_1146, new_AGEMA_signal_1145, y_rotated[11]}), .c ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, new_AGEMA_signal_1310, AdderIns_p6[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_12_U1 ( .a ({x_round_in_s3[12], x_round_in_s2[12], x_round_in_s1[12], x_round_in_s0[12]}), .b ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, new_AGEMA_signal_1148, y_rotated[12]}), .c ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, new_AGEMA_signal_1319, AdderIns_p6[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_13_U1 ( .a ({x_round_in_s3[13], x_round_in_s2[13], x_round_in_s1[13], x_round_in_s0[13]}), .b ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, y_rotated[13]}), .c ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, new_AGEMA_signal_1328, AdderIns_p6[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_14_U1 ( .a ({x_round_in_s3[14], x_round_in_s2[14], x_round_in_s1[14], x_round_in_s0[14]}), .b ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, y_rotated[14]}), .c ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, new_AGEMA_signal_1337, AdderIns_p6[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_15_U1 ( .a ({x_round_in_s3[15], x_round_in_s2[15], x_round_in_s1[15], x_round_in_s0[15]}), .b ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, new_AGEMA_signal_1157, y_rotated[15]}), .c ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, AdderIns_p6[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_16_U1 ( .a ({x_round_in_s3[16], x_round_in_s2[16], x_round_in_s1[16], x_round_in_s0[16]}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, new_AGEMA_signal_1160, y_rotated[16]}), .c ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, AdderIns_p6[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_17_U1 ( .a ({x_round_in_s3[17], x_round_in_s2[17], x_round_in_s1[17], x_round_in_s0[17]}), .b ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, new_AGEMA_signal_1163, y_rotated[17]}), .c ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, new_AGEMA_signal_1364, AdderIns_p6[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_18_U1 ( .a ({x_round_in_s3[18], x_round_in_s2[18], x_round_in_s1[18], x_round_in_s0[18]}), .b ({new_AGEMA_signal_1168, new_AGEMA_signal_1167, new_AGEMA_signal_1166, y_rotated[18]}), .c ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, new_AGEMA_signal_1373, AdderIns_p6[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_19_U1 ( .a ({x_round_in_s3[19], x_round_in_s2[19], x_round_in_s1[19], x_round_in_s0[19]}), .b ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, new_AGEMA_signal_1169, y_rotated[19]}), .c ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, new_AGEMA_signal_1382, AdderIns_p6[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_20_U1 ( .a ({x_round_in_s3[20], x_round_in_s2[20], x_round_in_s1[20], x_round_in_s0[20]}), .b ({new_AGEMA_signal_1174, new_AGEMA_signal_1173, new_AGEMA_signal_1172, y_rotated[20]}), .c ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, AdderIns_p6[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_21_U1 ( .a ({x_round_in_s3[21], x_round_in_s2[21], x_round_in_s1[21], x_round_in_s0[21]}), .b ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, new_AGEMA_signal_1175, y_rotated[21]}), .c ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, new_AGEMA_signal_1400, AdderIns_p6[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_22_U1 ( .a ({x_round_in_s3[22], x_round_in_s2[22], x_round_in_s1[22], x_round_in_s0[22]}), .b ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, y_rotated[22]}), .c ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, new_AGEMA_signal_1409, AdderIns_p6[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_23_U1 ( .a ({x_round_in_s3[23], x_round_in_s2[23], x_round_in_s1[23], x_round_in_s0[23]}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, new_AGEMA_signal_1181, y_rotated[23]}), .c ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, AdderIns_p6[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_24_U1 ( .a ({x_round_in_s3[24], x_round_in_s2[24], x_round_in_s1[24], x_round_in_s0[24]}), .b ({new_AGEMA_signal_1186, new_AGEMA_signal_1185, new_AGEMA_signal_1184, y_rotated[24]}), .c ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, AdderIns_p6[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_25_U1 ( .a ({x_round_in_s3[25], x_round_in_s2[25], x_round_in_s1[25], x_round_in_s0[25]}), .b ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, new_AGEMA_signal_1187, y_rotated[25]}), .c ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, new_AGEMA_signal_1436, AdderIns_p6[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_26_U1 ( .a ({x_round_in_s3[26], x_round_in_s2[26], x_round_in_s1[26], x_round_in_s0[26]}), .b ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, new_AGEMA_signal_1190, y_rotated[26]}), .c ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, new_AGEMA_signal_1445, AdderIns_p6[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_27_U1 ( .a ({x_round_in_s3[27], x_round_in_s2[27], x_round_in_s1[27], x_round_in_s0[27]}), .b ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, new_AGEMA_signal_1193, y_rotated[27]}), .c ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, AdderIns_p6[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_28_U1 ( .a ({x_round_in_s3[28], x_round_in_s2[28], x_round_in_s1[28], x_round_in_s0[28]}), .b ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, new_AGEMA_signal_1196, y_rotated[28]}), .c ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, new_AGEMA_signal_1463, AdderIns_p6[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_29_U1 ( .a ({x_round_in_s3[29], x_round_in_s2[29], x_round_in_s1[29], x_round_in_s0[29]}), .b ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, new_AGEMA_signal_1199, y_rotated[29]}), .c ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, new_AGEMA_signal_1472, AdderIns_p6[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_30_U1 ( .a ({x_round_in_s3[30], x_round_in_s2[30], x_round_in_s1[30], x_round_in_s0[30]}), .b ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, y_rotated[30]}), .c ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, new_AGEMA_signal_1481, AdderIns_p6[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_31_U1 ( .a ({x_round_in_s3[31], x_round_in_s2[31], x_round_in_s1[31], x_round_in_s0[31]}), .b ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, new_AGEMA_signal_1205, y_rotated[31]}), .c ({new_AGEMA_signal_1492, new_AGEMA_signal_1491, new_AGEMA_signal_1490, AdderIns_p6[31]}) ) ;
    //ClockGatingController #(10) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) U140 ( .a ({1'b0, 1'b0, 1'b0, round_constant[1]}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, new_AGEMA_signal_2027, sum[1]}), .c ({x_round_out_s3[1], x_round_out_s2[1], x_round_out_s1[1], x_round_out_s0[1]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_0_a1_U1 ( .a ({x_round_in_s3[0], x_round_in_s2[0], x_round_in_s1[0], x_round_in_s0[0]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, new_AGEMA_signal_1112, y_rotated[0]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, new_AGEMA_signal_1214, AdderIns_g1[0]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_1_a1_U1 ( .a ({x_round_in_s3[1], x_round_in_s2[1], x_round_in_s1[1], x_round_in_s0[1]}), .b ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, new_AGEMA_signal_1115, y_rotated[1]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, AdderIns_g1[1]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_2_a1_U1 ( .a ({x_round_in_s3[2], x_round_in_s2[2], x_round_in_s1[2], x_round_in_s0[2]}), .b ({new_AGEMA_signal_1120, new_AGEMA_signal_1119, new_AGEMA_signal_1118, y_rotated[2]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, new_AGEMA_signal_1232, AdderIns_g1[2]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_3_a1_U1 ( .a ({x_round_in_s3[3], x_round_in_s2[3], x_round_in_s1[3], x_round_in_s0[3]}), .b ({new_AGEMA_signal_1123, new_AGEMA_signal_1122, new_AGEMA_signal_1121, y_rotated[3]}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, new_AGEMA_signal_1241, AdderIns_g1[3]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_4_a1_U1 ( .a ({x_round_in_s3[4], x_round_in_s2[4], x_round_in_s1[4], x_round_in_s0[4]}), .b ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, new_AGEMA_signal_1124, y_rotated[4]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, new_AGEMA_signal_1250, AdderIns_g1[4]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_5_a1_U1 ( .a ({x_round_in_s3[5], x_round_in_s2[5], x_round_in_s1[5], x_round_in_s0[5]}), .b ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, new_AGEMA_signal_1127, y_rotated[5]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, new_AGEMA_signal_1259, AdderIns_g1[5]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_6_a1_U1 ( .a ({x_round_in_s3[6], x_round_in_s2[6], x_round_in_s1[6], x_round_in_s0[6]}), .b ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, new_AGEMA_signal_1130, y_rotated[6]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, new_AGEMA_signal_1268, AdderIns_g1[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_7_a1_U1 ( .a ({x_round_in_s3[7], x_round_in_s2[7], x_round_in_s1[7], x_round_in_s0[7]}), .b ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, new_AGEMA_signal_1133, y_rotated[7]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, new_AGEMA_signal_1277, AdderIns_g1[7]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_8_a1_U1 ( .a ({x_round_in_s3[8], x_round_in_s2[8], x_round_in_s1[8], x_round_in_s0[8]}), .b ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, new_AGEMA_signal_1136, y_rotated[8]}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, AdderIns_g1[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_9_a1_U1 ( .a ({x_round_in_s3[9], x_round_in_s2[9], x_round_in_s1[9], x_round_in_s0[9]}), .b ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, new_AGEMA_signal_1139, y_rotated[9]}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, new_AGEMA_signal_1295, AdderIns_g1[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_10_a1_U1 ( .a ({x_round_in_s3[10], x_round_in_s2[10], x_round_in_s1[10], x_round_in_s0[10]}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, new_AGEMA_signal_1142, y_rotated[10]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, new_AGEMA_signal_1304, AdderIns_g1[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_11_a1_U1 ( .a ({x_round_in_s3[11], x_round_in_s2[11], x_round_in_s1[11], x_round_in_s0[11]}), .b ({new_AGEMA_signal_1147, new_AGEMA_signal_1146, new_AGEMA_signal_1145, y_rotated[11]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, new_AGEMA_signal_1313, AdderIns_g1[11]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_12_a1_U1 ( .a ({x_round_in_s3[12], x_round_in_s2[12], x_round_in_s1[12], x_round_in_s0[12]}), .b ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, new_AGEMA_signal_1148, y_rotated[12]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, AdderIns_g1[12]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_13_a1_U1 ( .a ({x_round_in_s3[13], x_round_in_s2[13], x_round_in_s1[13], x_round_in_s0[13]}), .b ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, y_rotated[13]}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, AdderIns_g1[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_14_a1_U1 ( .a ({x_round_in_s3[14], x_round_in_s2[14], x_round_in_s1[14], x_round_in_s0[14]}), .b ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, y_rotated[14]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, new_AGEMA_signal_1340, AdderIns_g1[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_15_a1_U1 ( .a ({x_round_in_s3[15], x_round_in_s2[15], x_round_in_s1[15], x_round_in_s0[15]}), .b ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, new_AGEMA_signal_1157, y_rotated[15]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, new_AGEMA_signal_1349, AdderIns_g1[15]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_16_a1_U1 ( .a ({x_round_in_s3[16], x_round_in_s2[16], x_round_in_s1[16], x_round_in_s0[16]}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, new_AGEMA_signal_1160, y_rotated[16]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, new_AGEMA_signal_1358, AdderIns_g1[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_17_a1_U1 ( .a ({x_round_in_s3[17], x_round_in_s2[17], x_round_in_s1[17], x_round_in_s0[17]}), .b ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, new_AGEMA_signal_1163, y_rotated[17]}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, AdderIns_g1[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_18_a1_U1 ( .a ({x_round_in_s3[18], x_round_in_s2[18], x_round_in_s1[18], x_round_in_s0[18]}), .b ({new_AGEMA_signal_1168, new_AGEMA_signal_1167, new_AGEMA_signal_1166, y_rotated[18]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, new_AGEMA_signal_1376, AdderIns_g1[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_19_a1_U1 ( .a ({x_round_in_s3[19], x_round_in_s2[19], x_round_in_s1[19], x_round_in_s0[19]}), .b ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, new_AGEMA_signal_1169, y_rotated[19]}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, new_AGEMA_signal_1385, AdderIns_g1[19]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_20_a1_U1 ( .a ({x_round_in_s3[20], x_round_in_s2[20], x_round_in_s1[20], x_round_in_s0[20]}), .b ({new_AGEMA_signal_1174, new_AGEMA_signal_1173, new_AGEMA_signal_1172, y_rotated[20]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, AdderIns_g1[20]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_21_a1_U1 ( .a ({x_round_in_s3[21], x_round_in_s2[21], x_round_in_s1[21], x_round_in_s0[21]}), .b ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, new_AGEMA_signal_1175, y_rotated[21]}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, new_AGEMA_signal_1403, AdderIns_g1[21]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_22_a1_U1 ( .a ({x_round_in_s3[22], x_round_in_s2[22], x_round_in_s1[22], x_round_in_s0[22]}), .b ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, y_rotated[22]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, new_AGEMA_signal_1412, AdderIns_g1[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_23_a1_U1 ( .a ({x_round_in_s3[23], x_round_in_s2[23], x_round_in_s1[23], x_round_in_s0[23]}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, new_AGEMA_signal_1181, y_rotated[23]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, new_AGEMA_signal_1421, AdderIns_g1[23]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_24_a1_U1 ( .a ({x_round_in_s3[24], x_round_in_s2[24], x_round_in_s1[24], x_round_in_s0[24]}), .b ({new_AGEMA_signal_1186, new_AGEMA_signal_1185, new_AGEMA_signal_1184, y_rotated[24]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, new_AGEMA_signal_1430, AdderIns_g1[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_25_a1_U1 ( .a ({x_round_in_s3[25], x_round_in_s2[25], x_round_in_s1[25], x_round_in_s0[25]}), .b ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, new_AGEMA_signal_1187, y_rotated[25]}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, AdderIns_g1[25]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_26_a1_U1 ( .a ({x_round_in_s3[26], x_round_in_s2[26], x_round_in_s1[26], x_round_in_s0[26]}), .b ({new_AGEMA_signal_1192, new_AGEMA_signal_1191, new_AGEMA_signal_1190, y_rotated[26]}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, new_AGEMA_signal_1448, AdderIns_g1[26]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_27_a1_U1 ( .a ({x_round_in_s3[27], x_round_in_s2[27], x_round_in_s1[27], x_round_in_s0[27]}), .b ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, new_AGEMA_signal_1193, y_rotated[27]}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, new_AGEMA_signal_1457, AdderIns_g1[27]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_28_a1_U1 ( .a ({x_round_in_s3[28], x_round_in_s2[28], x_round_in_s1[28], x_round_in_s0[28]}), .b ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, new_AGEMA_signal_1196, y_rotated[28]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, new_AGEMA_signal_1466, AdderIns_g1[28]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_29_a1_U1 ( .a ({x_round_in_s3[29], x_round_in_s2[29], x_round_in_s1[29], x_round_in_s0[29]}), .b ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, new_AGEMA_signal_1199, y_rotated[29]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, new_AGEMA_signal_1475, AdderIns_g1[29]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s1_pg_30_a1_U1 ( .a ({x_round_in_s3[30], x_round_in_s2[30], x_round_in_s1[30], x_round_in_s0[30]}), .b ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, y_rotated[30]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, new_AGEMA_signal_1484, AdderIns_g1[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_gc_0_a1_U1 ( .a ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, new_AGEMA_signal_1214, AdderIns_g1[0]}), .b ({new_AGEMA_signal_1498, new_AGEMA_signal_1497, new_AGEMA_signal_1496, AdderIns_s2_gc_0_a1_t}), .c ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, AdderIns_g6[0]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, new_AGEMA_signal_1211, sum[0]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1498, new_AGEMA_signal_1497, new_AGEMA_signal_1496, AdderIns_s2_gc_0_a1_t}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_0_a2_U1 ( .a ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, new_AGEMA_signal_1211, sum[0]}), .b ({new_AGEMA_signal_1222, new_AGEMA_signal_1221, new_AGEMA_signal_1220, AdderIns_p6[1]}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, new_AGEMA_signal_1502, AdderIns_p2[0]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1222, new_AGEMA_signal_1221, new_AGEMA_signal_1220, AdderIns_p6[1]}), .b ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, new_AGEMA_signal_1229, AdderIns_p6[2]}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, new_AGEMA_signal_1508, AdderIns_p2[1]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, new_AGEMA_signal_1229, AdderIns_p6[2]}), .b ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, new_AGEMA_signal_1238, AdderIns_p6[3]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, new_AGEMA_signal_1514, AdderIns_p2[2]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, new_AGEMA_signal_1238, AdderIns_p6[3]}), .b ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, new_AGEMA_signal_1247, AdderIns_p6[4]}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, new_AGEMA_signal_1520, AdderIns_p2[3]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, new_AGEMA_signal_1247, AdderIns_p6[4]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, new_AGEMA_signal_1256, AdderIns_p6[5]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, new_AGEMA_signal_1526, AdderIns_p2[4]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, new_AGEMA_signal_1256, AdderIns_p6[5]}), .b ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, new_AGEMA_signal_1265, AdderIns_p6[6]}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1534, new_AGEMA_signal_1533, new_AGEMA_signal_1532, AdderIns_p2[5]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, new_AGEMA_signal_1265, AdderIns_p6[6]}), .b ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, AdderIns_p6[7]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, new_AGEMA_signal_1538, AdderIns_p2[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, AdderIns_p6[7]}), .b ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, AdderIns_p6[8]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, new_AGEMA_signal_1544, AdderIns_p2[7]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, AdderIns_p6[8]}), .b ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, new_AGEMA_signal_1292, AdderIns_p6[9]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, new_AGEMA_signal_1550, AdderIns_p2[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, new_AGEMA_signal_1292, AdderIns_p6[9]}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, new_AGEMA_signal_1301, AdderIns_p6[10]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, new_AGEMA_signal_1556, AdderIns_p2[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, new_AGEMA_signal_1301, AdderIns_p6[10]}), .b ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, new_AGEMA_signal_1310, AdderIns_p6[11]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, new_AGEMA_signal_1562, AdderIns_p2[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, new_AGEMA_signal_1310, AdderIns_p6[11]}), .b ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, new_AGEMA_signal_1319, AdderIns_p6[12]}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, new_AGEMA_signal_1568, AdderIns_p2[11]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, new_AGEMA_signal_1319, AdderIns_p6[12]}), .b ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, new_AGEMA_signal_1328, AdderIns_p6[13]}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1574, AdderIns_p2[12]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, new_AGEMA_signal_1328, AdderIns_p6[13]}), .b ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, new_AGEMA_signal_1337, AdderIns_p6[14]}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, new_AGEMA_signal_1580, AdderIns_p2[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, new_AGEMA_signal_1337, AdderIns_p6[14]}), .b ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, AdderIns_p6[15]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1586, AdderIns_p2[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_15_a2_U1 ( .a ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, AdderIns_p6[15]}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, AdderIns_p6[16]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, new_AGEMA_signal_1592, AdderIns_p2[15]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_16_a2_U1 ( .a ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, AdderIns_p6[16]}), .b ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, new_AGEMA_signal_1364, AdderIns_p6[17]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, new_AGEMA_signal_1598, AdderIns_p2[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_17_a2_U1 ( .a ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, new_AGEMA_signal_1364, AdderIns_p6[17]}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, new_AGEMA_signal_1373, AdderIns_p6[18]}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, new_AGEMA_signal_1604, AdderIns_p2[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_18_a2_U1 ( .a ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, new_AGEMA_signal_1373, AdderIns_p6[18]}), .b ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, new_AGEMA_signal_1382, AdderIns_p6[19]}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1610, AdderIns_p2[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_19_a2_U1 ( .a ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, new_AGEMA_signal_1382, AdderIns_p6[19]}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, AdderIns_p6[20]}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, new_AGEMA_signal_1616, AdderIns_p2[19]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_20_a2_U1 ( .a ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, AdderIns_p6[20]}), .b ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, new_AGEMA_signal_1400, AdderIns_p6[21]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, new_AGEMA_signal_1622, AdderIns_p2[20]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_21_a2_U1 ( .a ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, new_AGEMA_signal_1400, AdderIns_p6[21]}), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, new_AGEMA_signal_1409, AdderIns_p6[22]}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, new_AGEMA_signal_1628, AdderIns_p2[21]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_22_a2_U1 ( .a ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, new_AGEMA_signal_1409, AdderIns_p6[22]}), .b ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, AdderIns_p6[23]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, new_AGEMA_signal_1634, AdderIns_p2[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_23_a2_U1 ( .a ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, AdderIns_p6[23]}), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, AdderIns_p6[24]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, new_AGEMA_signal_1640, AdderIns_p2[23]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_24_a2_U1 ( .a ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, AdderIns_p6[24]}), .b ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, new_AGEMA_signal_1436, AdderIns_p6[25]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1646, AdderIns_p2[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_25_a2_U1 ( .a ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, new_AGEMA_signal_1436, AdderIns_p6[25]}), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, new_AGEMA_signal_1445, AdderIns_p6[26]}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1654, new_AGEMA_signal_1653, new_AGEMA_signal_1652, AdderIns_p2[25]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_26_a2_U1 ( .a ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, new_AGEMA_signal_1445, AdderIns_p6[26]}), .b ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, AdderIns_p6[27]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, new_AGEMA_signal_1658, AdderIns_p2[26]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_27_a2_U1 ( .a ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, AdderIns_p6[27]}), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, new_AGEMA_signal_1463, AdderIns_p6[28]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, new_AGEMA_signal_1664, AdderIns_p2[27]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_28_a2_U1 ( .a ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, new_AGEMA_signal_1463, AdderIns_p6[28]}), .b ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, new_AGEMA_signal_1472, AdderIns_p6[29]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, new_AGEMA_signal_1670, AdderIns_p2[28]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_29_a2_U1 ( .a ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, new_AGEMA_signal_1472, AdderIns_p6[29]}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, new_AGEMA_signal_1481, AdderIns_p6[30]}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, new_AGEMA_signal_1676, AdderIns_p2[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U11 ( .a ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1222, new_AGEMA_signal_1221, new_AGEMA_signal_1220, AdderIns_p6[1]}), .c ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, new_AGEMA_signal_2027, sum[1]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) U151 ( .a ({1'b0, 1'b0, 1'b0, round_constant[2]}), .b ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, sum[2]}), .c ({x_round_out_s3[2], x_round_out_s2[2], x_round_out_s1[2], x_round_out_s0[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U154 ( .a ({1'b0, 1'b0, 1'b0, round_constant[3]}), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, sum[3]}), .c ({x_round_out_s3[3], x_round_out_s2[3], x_round_out_s1[3], x_round_out_s0[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_0_a1_U1 ( .a ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, AdderIns_g1[1]}), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, new_AGEMA_signal_1499, AdderIns_s2_bc_0_a1_t}), .c ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, new_AGEMA_signal_1682, AdderIns_g2[1]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, new_AGEMA_signal_1214, AdderIns_g1[0]}), .b ({new_AGEMA_signal_1222, new_AGEMA_signal_1221, new_AGEMA_signal_1220, AdderIns_p6[1]}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, new_AGEMA_signal_1499, AdderIns_s2_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_1_a1_U1 ( .a ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, new_AGEMA_signal_1232, AdderIns_g1[2]}), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, new_AGEMA_signal_1505, AdderIns_s2_bc_1_a1_t}), .c ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, new_AGEMA_signal_1685, AdderIns_g2[2]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, AdderIns_g1[1]}), .b ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, new_AGEMA_signal_1229, AdderIns_p6[2]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, new_AGEMA_signal_1505, AdderIns_s2_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_2_a1_U1 ( .a ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, new_AGEMA_signal_1241, AdderIns_g1[3]}), .b ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, new_AGEMA_signal_1511, AdderIns_s2_bc_2_a1_t}), .c ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, new_AGEMA_signal_1688, AdderIns_g2[3]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, new_AGEMA_signal_1232, AdderIns_g1[2]}), .b ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, new_AGEMA_signal_1238, AdderIns_p6[3]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, new_AGEMA_signal_1511, AdderIns_s2_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_3_a1_U1 ( .a ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, new_AGEMA_signal_1250, AdderIns_g1[4]}), .b ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, new_AGEMA_signal_1517, AdderIns_s2_bc_3_a1_t}), .c ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, new_AGEMA_signal_1691, AdderIns_g2[4]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, new_AGEMA_signal_1241, AdderIns_g1[3]}), .b ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, new_AGEMA_signal_1247, AdderIns_p6[4]}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, new_AGEMA_signal_1517, AdderIns_s2_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_4_a1_U1 ( .a ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, new_AGEMA_signal_1259, AdderIns_g1[5]}), .b ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1523, AdderIns_s2_bc_4_a1_t}), .c ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, new_AGEMA_signal_1694, AdderIns_g2[5]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, new_AGEMA_signal_1250, AdderIns_g1[4]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, new_AGEMA_signal_1256, AdderIns_p6[5]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1523, AdderIns_s2_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_5_a1_U1 ( .a ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, new_AGEMA_signal_1268, AdderIns_g1[6]}), .b ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, new_AGEMA_signal_1529, AdderIns_s2_bc_5_a1_t}), .c ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, new_AGEMA_signal_1697, AdderIns_g2[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, new_AGEMA_signal_1259, AdderIns_g1[5]}), .b ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, new_AGEMA_signal_1265, AdderIns_p6[6]}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, new_AGEMA_signal_1529, AdderIns_s2_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_6_a1_U1 ( .a ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, new_AGEMA_signal_1277, AdderIns_g1[7]}), .b ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, new_AGEMA_signal_1535, AdderIns_s2_bc_6_a1_t}), .c ({new_AGEMA_signal_1702, new_AGEMA_signal_1701, new_AGEMA_signal_1700, AdderIns_g2[7]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, new_AGEMA_signal_1268, AdderIns_g1[6]}), .b ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, AdderIns_p6[7]}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, new_AGEMA_signal_1535, AdderIns_s2_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_7_a1_U1 ( .a ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, AdderIns_g1[8]}), .b ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, new_AGEMA_signal_1541, AdderIns_s2_bc_7_a1_t}), .c ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1703, AdderIns_g2[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, new_AGEMA_signal_1277, AdderIns_g1[7]}), .b ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, AdderIns_p6[8]}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, new_AGEMA_signal_1541, AdderIns_s2_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_8_a1_U1 ( .a ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, new_AGEMA_signal_1295, AdderIns_g1[9]}), .b ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, new_AGEMA_signal_1547, AdderIns_s2_bc_8_a1_t}), .c ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, new_AGEMA_signal_1706, AdderIns_g2[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, AdderIns_g1[8]}), .b ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, new_AGEMA_signal_1292, AdderIns_p6[9]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, new_AGEMA_signal_1547, AdderIns_s2_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_9_a1_U1 ( .a ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, new_AGEMA_signal_1304, AdderIns_g1[10]}), .b ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, new_AGEMA_signal_1553, AdderIns_s2_bc_9_a1_t}), .c ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, new_AGEMA_signal_1709, AdderIns_g2[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, new_AGEMA_signal_1295, AdderIns_g1[9]}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, new_AGEMA_signal_1301, AdderIns_p6[10]}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, new_AGEMA_signal_1553, AdderIns_s2_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_10_a1_U1 ( .a ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, new_AGEMA_signal_1313, AdderIns_g1[11]}), .b ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, new_AGEMA_signal_1559, AdderIns_s2_bc_10_a1_t}), .c ({new_AGEMA_signal_1714, new_AGEMA_signal_1713, new_AGEMA_signal_1712, AdderIns_g2[11]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, new_AGEMA_signal_1304, AdderIns_g1[10]}), .b ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, new_AGEMA_signal_1310, AdderIns_p6[11]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, new_AGEMA_signal_1559, AdderIns_s2_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_11_a1_U1 ( .a ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, AdderIns_g1[12]}), .b ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, new_AGEMA_signal_1565, AdderIns_s2_bc_11_a1_t}), .c ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, AdderIns_g2[12]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, new_AGEMA_signal_1313, AdderIns_g1[11]}), .b ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, new_AGEMA_signal_1319, AdderIns_p6[12]}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, new_AGEMA_signal_1565, AdderIns_s2_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_12_a1_U1 ( .a ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, AdderIns_g1[13]}), .b ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, new_AGEMA_signal_1571, AdderIns_s2_bc_12_a1_t}), .c ({new_AGEMA_signal_1720, new_AGEMA_signal_1719, new_AGEMA_signal_1718, AdderIns_g2[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, AdderIns_g1[12]}), .b ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, new_AGEMA_signal_1328, AdderIns_p6[13]}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, new_AGEMA_signal_1571, AdderIns_s2_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_13_a1_U1 ( .a ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, new_AGEMA_signal_1340, AdderIns_g1[14]}), .b ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, new_AGEMA_signal_1577, AdderIns_s2_bc_13_a1_t}), .c ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, new_AGEMA_signal_1721, AdderIns_g2[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, AdderIns_g1[13]}), .b ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, new_AGEMA_signal_1337, AdderIns_p6[14]}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, new_AGEMA_signal_1577, AdderIns_s2_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_14_a1_U1 ( .a ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, new_AGEMA_signal_1349, AdderIns_g1[15]}), .b ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, new_AGEMA_signal_1583, AdderIns_s2_bc_14_a1_t}), .c ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, new_AGEMA_signal_1724, AdderIns_g2[15]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, new_AGEMA_signal_1340, AdderIns_g1[14]}), .b ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, AdderIns_p6[15]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, new_AGEMA_signal_1583, AdderIns_s2_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_15_a1_U1 ( .a ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, new_AGEMA_signal_1358, AdderIns_g1[16]}), .b ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, new_AGEMA_signal_1589, AdderIns_s2_bc_15_a1_t}), .c ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, new_AGEMA_signal_1727, AdderIns_g2[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, new_AGEMA_signal_1349, AdderIns_g1[15]}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, AdderIns_p6[16]}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, new_AGEMA_signal_1589, AdderIns_s2_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_16_a1_U1 ( .a ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, AdderIns_g1[17]}), .b ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, new_AGEMA_signal_1595, AdderIns_s2_bc_16_a1_t}), .c ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, new_AGEMA_signal_1730, AdderIns_g2[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_16_a1_a1_U1 ( .a ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, new_AGEMA_signal_1358, AdderIns_g1[16]}), .b ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, new_AGEMA_signal_1364, AdderIns_p6[17]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, new_AGEMA_signal_1595, AdderIns_s2_bc_16_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_17_a1_U1 ( .a ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, new_AGEMA_signal_1376, AdderIns_g1[18]}), .b ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, new_AGEMA_signal_1601, AdderIns_s2_bc_17_a1_t}), .c ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, new_AGEMA_signal_1733, AdderIns_g2[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_17_a1_a1_U1 ( .a ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, AdderIns_g1[17]}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, new_AGEMA_signal_1373, AdderIns_p6[18]}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, new_AGEMA_signal_1601, AdderIns_s2_bc_17_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_18_a1_U1 ( .a ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, new_AGEMA_signal_1385, AdderIns_g1[19]}), .b ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, new_AGEMA_signal_1607, AdderIns_s2_bc_18_a1_t}), .c ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, new_AGEMA_signal_1736, AdderIns_g2[19]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_18_a1_a1_U1 ( .a ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, new_AGEMA_signal_1376, AdderIns_g1[18]}), .b ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, new_AGEMA_signal_1382, AdderIns_p6[19]}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, new_AGEMA_signal_1607, AdderIns_s2_bc_18_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_19_a1_U1 ( .a ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, AdderIns_g1[20]}), .b ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, new_AGEMA_signal_1613, AdderIns_s2_bc_19_a1_t}), .c ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, new_AGEMA_signal_1739, AdderIns_g2[20]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_19_a1_a1_U1 ( .a ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, new_AGEMA_signal_1385, AdderIns_g1[19]}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, AdderIns_p6[20]}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, new_AGEMA_signal_1613, AdderIns_s2_bc_19_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_20_a1_U1 ( .a ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, new_AGEMA_signal_1403, AdderIns_g1[21]}), .b ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, new_AGEMA_signal_1619, AdderIns_s2_bc_20_a1_t}), .c ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, new_AGEMA_signal_1742, AdderIns_g2[21]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_20_a1_a1_U1 ( .a ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, AdderIns_g1[20]}), .b ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, new_AGEMA_signal_1400, AdderIns_p6[21]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, new_AGEMA_signal_1619, AdderIns_s2_bc_20_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_21_a1_U1 ( .a ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, new_AGEMA_signal_1412, AdderIns_g1[22]}), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, new_AGEMA_signal_1625, AdderIns_s2_bc_21_a1_t}), .c ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, new_AGEMA_signal_1745, AdderIns_g2[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_21_a1_a1_U1 ( .a ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, new_AGEMA_signal_1403, AdderIns_g1[21]}), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, new_AGEMA_signal_1409, AdderIns_p6[22]}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, new_AGEMA_signal_1625, AdderIns_s2_bc_21_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_22_a1_U1 ( .a ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, new_AGEMA_signal_1421, AdderIns_g1[23]}), .b ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, new_AGEMA_signal_1631, AdderIns_s2_bc_22_a1_t}), .c ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, new_AGEMA_signal_1748, AdderIns_g2[23]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_22_a1_a1_U1 ( .a ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, new_AGEMA_signal_1412, AdderIns_g1[22]}), .b ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, AdderIns_p6[23]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, new_AGEMA_signal_1631, AdderIns_s2_bc_22_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_23_a1_U1 ( .a ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, new_AGEMA_signal_1430, AdderIns_g1[24]}), .b ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, new_AGEMA_signal_1637, AdderIns_s2_bc_23_a1_t}), .c ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, AdderIns_g2[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_23_a1_a1_U1 ( .a ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, new_AGEMA_signal_1421, AdderIns_g1[23]}), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, AdderIns_p6[24]}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, new_AGEMA_signal_1637, AdderIns_s2_bc_23_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_24_a1_U1 ( .a ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, AdderIns_g1[25]}), .b ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, new_AGEMA_signal_1643, AdderIns_s2_bc_24_a1_t}), .c ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, new_AGEMA_signal_1754, AdderIns_g2[25]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_24_a1_a1_U1 ( .a ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, new_AGEMA_signal_1430, AdderIns_g1[24]}), .b ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, new_AGEMA_signal_1436, AdderIns_p6[25]}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, new_AGEMA_signal_1643, AdderIns_s2_bc_24_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_25_a1_U1 ( .a ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, new_AGEMA_signal_1448, AdderIns_g1[26]}), .b ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, new_AGEMA_signal_1649, AdderIns_s2_bc_25_a1_t}), .c ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, new_AGEMA_signal_1757, AdderIns_g2[26]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_25_a1_a1_U1 ( .a ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, AdderIns_g1[25]}), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, new_AGEMA_signal_1445, AdderIns_p6[26]}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, new_AGEMA_signal_1649, AdderIns_s2_bc_25_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_26_a1_U1 ( .a ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, new_AGEMA_signal_1457, AdderIns_g1[27]}), .b ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, new_AGEMA_signal_1655, AdderIns_s2_bc_26_a1_t}), .c ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, new_AGEMA_signal_1760, AdderIns_g2[27]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_26_a1_a1_U1 ( .a ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, new_AGEMA_signal_1448, AdderIns_g1[26]}), .b ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, AdderIns_p6[27]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, new_AGEMA_signal_1655, AdderIns_s2_bc_26_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_27_a1_U1 ( .a ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, new_AGEMA_signal_1466, AdderIns_g1[28]}), .b ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, new_AGEMA_signal_1661, AdderIns_s2_bc_27_a1_t}), .c ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, new_AGEMA_signal_1763, AdderIns_g2[28]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_27_a1_a1_U1 ( .a ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, new_AGEMA_signal_1457, AdderIns_g1[27]}), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, new_AGEMA_signal_1463, AdderIns_p6[28]}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, new_AGEMA_signal_1661, AdderIns_s2_bc_27_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_28_a1_U1 ( .a ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, new_AGEMA_signal_1475, AdderIns_g1[29]}), .b ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, new_AGEMA_signal_1667, AdderIns_s2_bc_28_a1_t}), .c ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, new_AGEMA_signal_1766, AdderIns_g2[29]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_28_a1_a1_U1 ( .a ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, new_AGEMA_signal_1466, AdderIns_g1[28]}), .b ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, new_AGEMA_signal_1472, AdderIns_p6[29]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, new_AGEMA_signal_1667, AdderIns_s2_bc_28_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_29_a1_U1 ( .a ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, new_AGEMA_signal_1484, AdderIns_g1[30]}), .b ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, new_AGEMA_signal_1673, AdderIns_s2_bc_29_a1_t}), .c ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, new_AGEMA_signal_1769, AdderIns_g2[30]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s2_bc_29_a1_a1_U1 ( .a ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, new_AGEMA_signal_1475, AdderIns_g1[29]}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, new_AGEMA_signal_1481, AdderIns_p6[30]}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, new_AGEMA_signal_1673, AdderIns_s2_bc_29_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_gc_0_a1_U1 ( .a ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, new_AGEMA_signal_1682, AdderIns_g2[1]}), .b ({new_AGEMA_signal_1774, new_AGEMA_signal_1773, new_AGEMA_signal_1772, AdderIns_s3_gc_0_a1_t}), .c ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, new_AGEMA_signal_1859, AdderIns_g6[1]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, new_AGEMA_signal_1502, AdderIns_p2[0]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1774, new_AGEMA_signal_1773, new_AGEMA_signal_1772, AdderIns_s3_gc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_gc_1_a1_U1 ( .a ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, new_AGEMA_signal_1685, AdderIns_g2[2]}), .b ({new_AGEMA_signal_1864, new_AGEMA_signal_1863, new_AGEMA_signal_1862, AdderIns_s3_gc_1_a1_t}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, AdderIns_g6[2]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, new_AGEMA_signal_1508, AdderIns_p2[1]}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1864, new_AGEMA_signal_1863, new_AGEMA_signal_1862, AdderIns_s3_gc_1_a1_t}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_0_a2_U1 ( .a ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, new_AGEMA_signal_1502, AdderIns_p2[0]}), .b ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, new_AGEMA_signal_1514, AdderIns_p2[2]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, new_AGEMA_signal_1775, AdderIns_p3[0]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, new_AGEMA_signal_1508, AdderIns_p2[1]}), .b ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, new_AGEMA_signal_1520, AdderIns_p2[3]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, new_AGEMA_signal_1778, AdderIns_p3[1]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, new_AGEMA_signal_1514, AdderIns_p2[2]}), .b ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, new_AGEMA_signal_1526, AdderIns_p2[4]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, new_AGEMA_signal_1781, AdderIns_p3[2]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, new_AGEMA_signal_1520, AdderIns_p2[3]}), .b ({new_AGEMA_signal_1534, new_AGEMA_signal_1533, new_AGEMA_signal_1532, AdderIns_p2[5]}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, new_AGEMA_signal_1784, AdderIns_p3[3]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, new_AGEMA_signal_1526, AdderIns_p2[4]}), .b ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, new_AGEMA_signal_1538, AdderIns_p2[6]}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, new_AGEMA_signal_1787, AdderIns_p3[4]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1534, new_AGEMA_signal_1533, new_AGEMA_signal_1532, AdderIns_p2[5]}), .b ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, new_AGEMA_signal_1544, AdderIns_p2[7]}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_1792, new_AGEMA_signal_1791, new_AGEMA_signal_1790, AdderIns_p3[5]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, new_AGEMA_signal_1538, AdderIns_p2[6]}), .b ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, new_AGEMA_signal_1550, AdderIns_p2[8]}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, new_AGEMA_signal_1793, AdderIns_p3[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, new_AGEMA_signal_1544, AdderIns_p2[7]}), .b ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, new_AGEMA_signal_1556, AdderIns_p2[9]}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, new_AGEMA_signal_1796, AdderIns_p3[7]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, new_AGEMA_signal_1550, AdderIns_p2[8]}), .b ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, new_AGEMA_signal_1562, AdderIns_p2[10]}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, new_AGEMA_signal_1799, AdderIns_p3[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, new_AGEMA_signal_1556, AdderIns_p2[9]}), .b ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, new_AGEMA_signal_1568, AdderIns_p2[11]}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, new_AGEMA_signal_1802, AdderIns_p3[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, new_AGEMA_signal_1562, AdderIns_p2[10]}), .b ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1574, AdderIns_p2[12]}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, new_AGEMA_signal_1805, AdderIns_p3[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, new_AGEMA_signal_1568, AdderIns_p2[11]}), .b ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, new_AGEMA_signal_1580, AdderIns_p2[13]}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, new_AGEMA_signal_1808, AdderIns_p3[11]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1574, AdderIns_p2[12]}), .b ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1586, AdderIns_p2[14]}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, new_AGEMA_signal_1811, AdderIns_p3[12]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, new_AGEMA_signal_1580, AdderIns_p2[13]}), .b ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, new_AGEMA_signal_1592, AdderIns_p2[15]}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, new_AGEMA_signal_1814, AdderIns_p3[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1586, AdderIns_p2[14]}), .b ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, new_AGEMA_signal_1598, AdderIns_p2[16]}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, new_AGEMA_signal_1817, AdderIns_p3[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_15_a2_U1 ( .a ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, new_AGEMA_signal_1592, AdderIns_p2[15]}), .b ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, new_AGEMA_signal_1604, AdderIns_p2[17]}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_1822, new_AGEMA_signal_1821, new_AGEMA_signal_1820, AdderIns_p3[15]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_16_a2_U1 ( .a ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, new_AGEMA_signal_1598, AdderIns_p2[16]}), .b ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1610, AdderIns_p2[18]}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, new_AGEMA_signal_1823, AdderIns_p3[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_17_a2_U1 ( .a ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, new_AGEMA_signal_1604, AdderIns_p2[17]}), .b ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, new_AGEMA_signal_1616, AdderIns_p2[19]}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, AdderIns_p3[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_18_a2_U1 ( .a ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1610, AdderIns_p2[18]}), .b ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, new_AGEMA_signal_1622, AdderIns_p2[20]}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, new_AGEMA_signal_1829, AdderIns_p3[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_19_a2_U1 ( .a ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, new_AGEMA_signal_1616, AdderIns_p2[19]}), .b ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, new_AGEMA_signal_1628, AdderIns_p2[21]}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, new_AGEMA_signal_1832, AdderIns_p3[19]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_20_a2_U1 ( .a ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, new_AGEMA_signal_1622, AdderIns_p2[20]}), .b ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, new_AGEMA_signal_1634, AdderIns_p2[22]}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, new_AGEMA_signal_1835, AdderIns_p3[20]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_21_a2_U1 ( .a ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, new_AGEMA_signal_1628, AdderIns_p2[21]}), .b ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, new_AGEMA_signal_1640, AdderIns_p2[23]}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, new_AGEMA_signal_1838, AdderIns_p3[21]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_22_a2_U1 ( .a ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, new_AGEMA_signal_1634, AdderIns_p2[22]}), .b ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1646, AdderIns_p2[24]}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, new_AGEMA_signal_1841, AdderIns_p3[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_23_a2_U1 ( .a ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, new_AGEMA_signal_1640, AdderIns_p2[23]}), .b ({new_AGEMA_signal_1654, new_AGEMA_signal_1653, new_AGEMA_signal_1652, AdderIns_p2[25]}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, new_AGEMA_signal_1844, AdderIns_p3[23]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_24_a2_U1 ( .a ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1646, AdderIns_p2[24]}), .b ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, new_AGEMA_signal_1658, AdderIns_p2[26]}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1847, AdderIns_p3[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_25_a2_U1 ( .a ({new_AGEMA_signal_1654, new_AGEMA_signal_1653, new_AGEMA_signal_1652, AdderIns_p2[25]}), .b ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, new_AGEMA_signal_1664, AdderIns_p2[27]}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_1852, new_AGEMA_signal_1851, new_AGEMA_signal_1850, AdderIns_p3[25]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_26_a2_U1 ( .a ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, new_AGEMA_signal_1658, AdderIns_p2[26]}), .b ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, new_AGEMA_signal_1670, AdderIns_p2[28]}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, new_AGEMA_signal_1853, AdderIns_p3[26]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_27_a2_U1 ( .a ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, new_AGEMA_signal_1664, AdderIns_p2[27]}), .b ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, new_AGEMA_signal_1676, AdderIns_p2[29]}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, new_AGEMA_signal_1856, AdderIns_p3[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U25 ( .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, AdderIns_g6[2]}), .b ({new_AGEMA_signal_1240, new_AGEMA_signal_1239, new_AGEMA_signal_1238, AdderIns_p6[3]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, sum[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U22 ( .a ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, new_AGEMA_signal_1859, AdderIns_g6[1]}), .b ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, new_AGEMA_signal_1229, AdderIns_p6[2]}), .c ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, sum[2]}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) U155 ( .a ({1'b0, 1'b0, 1'b0, round_constant[4]}), .b ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, new_AGEMA_signal_2384, sum[4]}), .c ({x_round_out_s3[4], x_round_out_s2[4], x_round_out_s1[4], x_round_out_s0[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U156 ( .a ({1'b0, 1'b0, 1'b0, round_constant[5]}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, sum[5]}), .c ({x_round_out_s3[5], x_round_out_s2[5], x_round_out_s1[5], x_round_out_s0[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U157 ( .a ({1'b0, 1'b0, 1'b0, round_constant[6]}), .b ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, new_AGEMA_signal_2378, sum[6]}), .c ({x_round_out_s3[6], x_round_out_s2[6], x_round_out_s1[6], x_round_out_s0[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U158 ( .a ({1'b0, 1'b0, 1'b0, round_constant[7]}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, sum[7]}), .c ({x_round_out_s3[7], x_round_out_s2[7], x_round_out_s1[7], x_round_out_s0[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_0_a1_U1 ( .a ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, new_AGEMA_signal_1688, AdderIns_g2[3]}), .b ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, new_AGEMA_signal_1865, AdderIns_s3_bc_0_a1_t}), .c ({new_AGEMA_signal_2038, new_AGEMA_signal_2037, new_AGEMA_signal_2036, AdderIns_g3[3]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, new_AGEMA_signal_1682, AdderIns_g2[1]}), .b ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, new_AGEMA_signal_1514, AdderIns_p2[2]}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, new_AGEMA_signal_1865, AdderIns_s3_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_1_a1_U1 ( .a ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, new_AGEMA_signal_1691, AdderIns_g2[4]}), .b ({new_AGEMA_signal_1870, new_AGEMA_signal_1869, new_AGEMA_signal_1868, AdderIns_s3_bc_1_a1_t}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, AdderIns_g3[4]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, new_AGEMA_signal_1685, AdderIns_g2[2]}), .b ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, new_AGEMA_signal_1520, AdderIns_p2[3]}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_1870, new_AGEMA_signal_1869, new_AGEMA_signal_1868, AdderIns_s3_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_2_a1_U1 ( .a ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, new_AGEMA_signal_1694, AdderIns_g2[5]}), .b ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, new_AGEMA_signal_1871, AdderIns_s3_bc_2_a1_t}), .c ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, AdderIns_g3[5]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, new_AGEMA_signal_1688, AdderIns_g2[3]}), .b ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, new_AGEMA_signal_1526, AdderIns_p2[4]}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, new_AGEMA_signal_1871, AdderIns_s3_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_3_a1_U1 ( .a ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, new_AGEMA_signal_1697, AdderIns_g2[6]}), .b ({new_AGEMA_signal_1876, new_AGEMA_signal_1875, new_AGEMA_signal_1874, AdderIns_s3_bc_3_a1_t}), .c ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, new_AGEMA_signal_2045, AdderIns_g3[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, new_AGEMA_signal_1691, AdderIns_g2[4]}), .b ({new_AGEMA_signal_1534, new_AGEMA_signal_1533, new_AGEMA_signal_1532, AdderIns_p2[5]}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_1876, new_AGEMA_signal_1875, new_AGEMA_signal_1874, AdderIns_s3_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_4_a1_U1 ( .a ({new_AGEMA_signal_1702, new_AGEMA_signal_1701, new_AGEMA_signal_1700, AdderIns_g2[7]}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, new_AGEMA_signal_1877, AdderIns_s3_bc_4_a1_t}), .c ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, AdderIns_g3[7]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, new_AGEMA_signal_1694, AdderIns_g2[5]}), .b ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, new_AGEMA_signal_1538, AdderIns_p2[6]}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, new_AGEMA_signal_1877, AdderIns_s3_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_5_a1_U1 ( .a ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1703, AdderIns_g2[8]}), .b ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, new_AGEMA_signal_1880, AdderIns_s3_bc_5_a1_t}), .c ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, new_AGEMA_signal_2051, AdderIns_g3[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, new_AGEMA_signal_1697, AdderIns_g2[6]}), .b ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, new_AGEMA_signal_1544, AdderIns_p2[7]}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, new_AGEMA_signal_1880, AdderIns_s3_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_6_a1_U1 ( .a ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, new_AGEMA_signal_1706, AdderIns_g2[9]}), .b ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, new_AGEMA_signal_1883, AdderIns_s3_bc_6_a1_t}), .c ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, AdderIns_g3[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_1702, new_AGEMA_signal_1701, new_AGEMA_signal_1700, AdderIns_g2[7]}), .b ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, new_AGEMA_signal_1550, AdderIns_p2[8]}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, new_AGEMA_signal_1883, AdderIns_s3_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_7_a1_U1 ( .a ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, new_AGEMA_signal_1709, AdderIns_g2[10]}), .b ({new_AGEMA_signal_1888, new_AGEMA_signal_1887, new_AGEMA_signal_1886, AdderIns_s3_bc_7_a1_t}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, new_AGEMA_signal_2057, AdderIns_g3[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1703, AdderIns_g2[8]}), .b ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, new_AGEMA_signal_1556, AdderIns_p2[9]}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_1888, new_AGEMA_signal_1887, new_AGEMA_signal_1886, AdderIns_s3_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_8_a1_U1 ( .a ({new_AGEMA_signal_1714, new_AGEMA_signal_1713, new_AGEMA_signal_1712, AdderIns_g2[11]}), .b ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, new_AGEMA_signal_1889, AdderIns_s3_bc_8_a1_t}), .c ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, new_AGEMA_signal_2060, AdderIns_g3[11]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, new_AGEMA_signal_1706, AdderIns_g2[9]}), .b ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, new_AGEMA_signal_1562, AdderIns_p2[10]}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, new_AGEMA_signal_1889, AdderIns_s3_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_9_a1_U1 ( .a ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, AdderIns_g2[12]}), .b ({new_AGEMA_signal_1894, new_AGEMA_signal_1893, new_AGEMA_signal_1892, AdderIns_s3_bc_9_a1_t}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, AdderIns_g3[12]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, new_AGEMA_signal_1709, AdderIns_g2[10]}), .b ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, new_AGEMA_signal_1568, AdderIns_p2[11]}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_1894, new_AGEMA_signal_1893, new_AGEMA_signal_1892, AdderIns_s3_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_10_a1_U1 ( .a ({new_AGEMA_signal_1720, new_AGEMA_signal_1719, new_AGEMA_signal_1718, AdderIns_g2[13]}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, new_AGEMA_signal_1895, AdderIns_s3_bc_10_a1_t}), .c ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, AdderIns_g3[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_1714, new_AGEMA_signal_1713, new_AGEMA_signal_1712, AdderIns_g2[11]}), .b ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1574, AdderIns_p2[12]}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, new_AGEMA_signal_1895, AdderIns_s3_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_11_a1_U1 ( .a ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, new_AGEMA_signal_1721, AdderIns_g2[14]}), .b ({new_AGEMA_signal_1900, new_AGEMA_signal_1899, new_AGEMA_signal_1898, AdderIns_s3_bc_11_a1_t}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, AdderIns_g3[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, AdderIns_g2[12]}), .b ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, new_AGEMA_signal_1580, AdderIns_p2[13]}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_1900, new_AGEMA_signal_1899, new_AGEMA_signal_1898, AdderIns_s3_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_12_a1_U1 ( .a ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, new_AGEMA_signal_1724, AdderIns_g2[15]}), .b ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, new_AGEMA_signal_1901, AdderIns_s3_bc_12_a1_t}), .c ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, AdderIns_g3[15]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_1720, new_AGEMA_signal_1719, new_AGEMA_signal_1718, AdderIns_g2[13]}), .b ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1586, AdderIns_p2[14]}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, new_AGEMA_signal_1901, AdderIns_s3_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_13_a1_U1 ( .a ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, new_AGEMA_signal_1727, AdderIns_g2[16]}), .b ({new_AGEMA_signal_1906, new_AGEMA_signal_1905, new_AGEMA_signal_1904, AdderIns_s3_bc_13_a1_t}), .c ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, new_AGEMA_signal_2075, AdderIns_g3[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, new_AGEMA_signal_1721, AdderIns_g2[14]}), .b ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, new_AGEMA_signal_1592, AdderIns_p2[15]}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_1906, new_AGEMA_signal_1905, new_AGEMA_signal_1904, AdderIns_s3_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_14_a1_U1 ( .a ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, new_AGEMA_signal_1730, AdderIns_g2[17]}), .b ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, new_AGEMA_signal_1907, AdderIns_s3_bc_14_a1_t}), .c ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, AdderIns_g3[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, new_AGEMA_signal_1724, AdderIns_g2[15]}), .b ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, new_AGEMA_signal_1598, AdderIns_p2[16]}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, new_AGEMA_signal_1907, AdderIns_s3_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_15_a1_U1 ( .a ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, new_AGEMA_signal_1733, AdderIns_g2[18]}), .b ({new_AGEMA_signal_1912, new_AGEMA_signal_1911, new_AGEMA_signal_1910, AdderIns_s3_bc_15_a1_t}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, new_AGEMA_signal_2081, AdderIns_g3[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, new_AGEMA_signal_1727, AdderIns_g2[16]}), .b ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, new_AGEMA_signal_1604, AdderIns_p2[17]}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_1912, new_AGEMA_signal_1911, new_AGEMA_signal_1910, AdderIns_s3_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_16_a1_U1 ( .a ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, new_AGEMA_signal_1736, AdderIns_g2[19]}), .b ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, new_AGEMA_signal_1913, AdderIns_s3_bc_16_a1_t}), .c ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, AdderIns_g3[19]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_16_a1_a1_U1 ( .a ({new_AGEMA_signal_1732, new_AGEMA_signal_1731, new_AGEMA_signal_1730, AdderIns_g2[17]}), .b ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1610, AdderIns_p2[18]}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, new_AGEMA_signal_1913, AdderIns_s3_bc_16_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_17_a1_U1 ( .a ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, new_AGEMA_signal_1739, AdderIns_g2[20]}), .b ({new_AGEMA_signal_1918, new_AGEMA_signal_1917, new_AGEMA_signal_1916, AdderIns_s3_bc_17_a1_t}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, AdderIns_g3[20]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_17_a1_a1_U1 ( .a ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, new_AGEMA_signal_1733, AdderIns_g2[18]}), .b ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, new_AGEMA_signal_1616, AdderIns_p2[19]}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_1918, new_AGEMA_signal_1917, new_AGEMA_signal_1916, AdderIns_s3_bc_17_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_18_a1_U1 ( .a ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, new_AGEMA_signal_1742, AdderIns_g2[21]}), .b ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, new_AGEMA_signal_1919, AdderIns_s3_bc_18_a1_t}), .c ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, AdderIns_g3[21]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_18_a1_a1_U1 ( .a ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, new_AGEMA_signal_1736, AdderIns_g2[19]}), .b ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, new_AGEMA_signal_1622, AdderIns_p2[20]}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, new_AGEMA_signal_1919, AdderIns_s3_bc_18_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_19_a1_U1 ( .a ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, new_AGEMA_signal_1745, AdderIns_g2[22]}), .b ({new_AGEMA_signal_1924, new_AGEMA_signal_1923, new_AGEMA_signal_1922, AdderIns_s3_bc_19_a1_t}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, AdderIns_g3[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_19_a1_a1_U1 ( .a ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, new_AGEMA_signal_1739, AdderIns_g2[20]}), .b ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, new_AGEMA_signal_1628, AdderIns_p2[21]}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_1924, new_AGEMA_signal_1923, new_AGEMA_signal_1922, AdderIns_s3_bc_19_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_20_a1_U1 ( .a ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, new_AGEMA_signal_1748, AdderIns_g2[23]}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, new_AGEMA_signal_1925, AdderIns_s3_bc_20_a1_t}), .c ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, new_AGEMA_signal_2096, AdderIns_g3[23]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_20_a1_a1_U1 ( .a ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, new_AGEMA_signal_1742, AdderIns_g2[21]}), .b ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, new_AGEMA_signal_1634, AdderIns_p2[22]}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, new_AGEMA_signal_1925, AdderIns_s3_bc_20_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_21_a1_U1 ( .a ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, AdderIns_g2[24]}), .b ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, new_AGEMA_signal_1928, AdderIns_s3_bc_21_a1_t}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, AdderIns_g3[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_21_a1_a1_U1 ( .a ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, new_AGEMA_signal_1745, AdderIns_g2[22]}), .b ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, new_AGEMA_signal_1640, AdderIns_p2[23]}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, new_AGEMA_signal_1928, AdderIns_s3_bc_21_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_22_a1_U1 ( .a ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, new_AGEMA_signal_1754, AdderIns_g2[25]}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, new_AGEMA_signal_1931, AdderIns_s3_bc_22_a1_t}), .c ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, AdderIns_g3[25]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_22_a1_a1_U1 ( .a ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, new_AGEMA_signal_1748, AdderIns_g2[23]}), .b ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1646, AdderIns_p2[24]}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, new_AGEMA_signal_1931, AdderIns_s3_bc_22_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_23_a1_U1 ( .a ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, new_AGEMA_signal_1757, AdderIns_g2[26]}), .b ({new_AGEMA_signal_1936, new_AGEMA_signal_1935, new_AGEMA_signal_1934, AdderIns_s3_bc_23_a1_t}), .c ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, new_AGEMA_signal_2105, AdderIns_g3[26]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_23_a1_a1_U1 ( .a ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, AdderIns_g2[24]}), .b ({new_AGEMA_signal_1654, new_AGEMA_signal_1653, new_AGEMA_signal_1652, AdderIns_p2[25]}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_1936, new_AGEMA_signal_1935, new_AGEMA_signal_1934, AdderIns_s3_bc_23_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_24_a1_U1 ( .a ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, new_AGEMA_signal_1760, AdderIns_g2[27]}), .b ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, new_AGEMA_signal_1937, AdderIns_s3_bc_24_a1_t}), .c ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, AdderIns_g3[27]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_24_a1_a1_U1 ( .a ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, new_AGEMA_signal_1754, AdderIns_g2[25]}), .b ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, new_AGEMA_signal_1658, AdderIns_p2[26]}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, new_AGEMA_signal_1937, AdderIns_s3_bc_24_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_25_a1_U1 ( .a ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, new_AGEMA_signal_1763, AdderIns_g2[28]}), .b ({new_AGEMA_signal_1942, new_AGEMA_signal_1941, new_AGEMA_signal_1940, AdderIns_s3_bc_25_a1_t}), .c ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, new_AGEMA_signal_2111, AdderIns_g3[28]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_25_a1_a1_U1 ( .a ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, new_AGEMA_signal_1757, AdderIns_g2[26]}), .b ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, new_AGEMA_signal_1664, AdderIns_p2[27]}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_1942, new_AGEMA_signal_1941, new_AGEMA_signal_1940, AdderIns_s3_bc_25_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_26_a1_U1 ( .a ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, new_AGEMA_signal_1766, AdderIns_g2[29]}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, new_AGEMA_signal_1943, AdderIns_s3_bc_26_a1_t}), .c ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, new_AGEMA_signal_2114, AdderIns_g3[29]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_26_a1_a1_U1 ( .a ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, new_AGEMA_signal_1760, AdderIns_g2[27]}), .b ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, new_AGEMA_signal_1670, AdderIns_p2[28]}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, new_AGEMA_signal_1943, AdderIns_s3_bc_26_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_27_a1_U1 ( .a ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, new_AGEMA_signal_1769, AdderIns_g2[30]}), .b ({new_AGEMA_signal_1948, new_AGEMA_signal_1947, new_AGEMA_signal_1946, AdderIns_s3_bc_27_a1_t}), .c ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, new_AGEMA_signal_2117, AdderIns_g3[30]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s3_bc_27_a1_a1_U1 ( .a ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, new_AGEMA_signal_1763, AdderIns_g2[28]}), .b ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, new_AGEMA_signal_1676, AdderIns_p2[29]}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_1948, new_AGEMA_signal_1947, new_AGEMA_signal_1946, AdderIns_s3_bc_27_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_gc_0_a1_U1 ( .a ({new_AGEMA_signal_2038, new_AGEMA_signal_2037, new_AGEMA_signal_2036, AdderIns_g3[3]}), .b ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, new_AGEMA_signal_1949, AdderIns_s4_gc_0_a1_t}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, AdderIns_g6[3]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, new_AGEMA_signal_1775, AdderIns_p3[0]}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, new_AGEMA_signal_1949, AdderIns_s4_gc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_gc_1_a1_U1 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, AdderIns_g3[4]}), .b ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, new_AGEMA_signal_1952, AdderIns_s4_gc_1_a1_t}), .c ({new_AGEMA_signal_2188, new_AGEMA_signal_2187, new_AGEMA_signal_2186, AdderIns_g6[4]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, new_AGEMA_signal_1778, AdderIns_p3[1]}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, new_AGEMA_signal_1952, AdderIns_s4_gc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_gc_2_a1_U1 ( .a ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, AdderIns_g3[5]}), .b ({new_AGEMA_signal_2122, new_AGEMA_signal_2121, new_AGEMA_signal_2120, AdderIns_s4_gc_2_a1_t}), .c ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, AdderIns_g6[5]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_gc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, new_AGEMA_signal_1859, AdderIns_g6[1]}), .b ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, new_AGEMA_signal_1781, AdderIns_p3[2]}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_2122, new_AGEMA_signal_2121, new_AGEMA_signal_2120, AdderIns_s4_gc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_gc_3_a1_U1 ( .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, new_AGEMA_signal_2045, AdderIns_g3[6]}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, new_AGEMA_signal_2192, AdderIns_s4_gc_3_a1_t}), .c ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, new_AGEMA_signal_2285, AdderIns_g6[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_gc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, AdderIns_g6[2]}), .b ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, new_AGEMA_signal_1784, AdderIns_p3[3]}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, new_AGEMA_signal_2192, AdderIns_s4_gc_3_a1_t}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_0_a2_U1 ( .a ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, new_AGEMA_signal_1775, AdderIns_p3[0]}), .b ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, new_AGEMA_signal_1787, AdderIns_p3[4]}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, new_AGEMA_signal_1955, AdderIns_p4[0]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, new_AGEMA_signal_1778, AdderIns_p3[1]}), .b ({new_AGEMA_signal_1792, new_AGEMA_signal_1791, new_AGEMA_signal_1790, AdderIns_p3[5]}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_1960, new_AGEMA_signal_1959, new_AGEMA_signal_1958, AdderIns_p4[1]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, new_AGEMA_signal_1781, AdderIns_p3[2]}), .b ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, new_AGEMA_signal_1793, AdderIns_p3[6]}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, new_AGEMA_signal_1961, AdderIns_p4[2]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, new_AGEMA_signal_1784, AdderIns_p3[3]}), .b ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, new_AGEMA_signal_1796, AdderIns_p3[7]}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_1966, new_AGEMA_signal_1965, new_AGEMA_signal_1964, AdderIns_p4[3]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, new_AGEMA_signal_1787, AdderIns_p3[4]}), .b ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, new_AGEMA_signal_1799, AdderIns_p3[8]}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, new_AGEMA_signal_1967, AdderIns_p4[4]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1792, new_AGEMA_signal_1791, new_AGEMA_signal_1790, AdderIns_p3[5]}), .b ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, new_AGEMA_signal_1802, AdderIns_p3[9]}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_1972, new_AGEMA_signal_1971, new_AGEMA_signal_1970, AdderIns_p4[5]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, new_AGEMA_signal_1793, AdderIns_p3[6]}), .b ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, new_AGEMA_signal_1805, AdderIns_p3[10]}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, new_AGEMA_signal_1973, AdderIns_p4[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, new_AGEMA_signal_1796, AdderIns_p3[7]}), .b ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, new_AGEMA_signal_1808, AdderIns_p3[11]}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, new_AGEMA_signal_1976, AdderIns_p4[7]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, new_AGEMA_signal_1799, AdderIns_p3[8]}), .b ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, new_AGEMA_signal_1811, AdderIns_p3[12]}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, new_AGEMA_signal_1979, AdderIns_p4[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, new_AGEMA_signal_1802, AdderIns_p3[9]}), .b ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, new_AGEMA_signal_1814, AdderIns_p3[13]}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1982, AdderIns_p4[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, new_AGEMA_signal_1805, AdderIns_p3[10]}), .b ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, new_AGEMA_signal_1817, AdderIns_p3[14]}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, AdderIns_p4[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, new_AGEMA_signal_1808, AdderIns_p3[11]}), .b ({new_AGEMA_signal_1822, new_AGEMA_signal_1821, new_AGEMA_signal_1820, AdderIns_p3[15]}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, new_AGEMA_signal_1988, AdderIns_p4[11]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, new_AGEMA_signal_1811, AdderIns_p3[12]}), .b ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, new_AGEMA_signal_1823, AdderIns_p3[16]}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1991, AdderIns_p4[12]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, new_AGEMA_signal_1814, AdderIns_p3[13]}), .b ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, AdderIns_p3[17]}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, AdderIns_p4[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, new_AGEMA_signal_1817, AdderIns_p3[14]}), .b ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, new_AGEMA_signal_1829, AdderIns_p3[18]}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, new_AGEMA_signal_1997, AdderIns_p4[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_15_a2_U1 ( .a ({new_AGEMA_signal_1822, new_AGEMA_signal_1821, new_AGEMA_signal_1820, AdderIns_p3[15]}), .b ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, new_AGEMA_signal_1832, AdderIns_p3[19]}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_2002, new_AGEMA_signal_2001, new_AGEMA_signal_2000, AdderIns_p4[15]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_16_a2_U1 ( .a ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, new_AGEMA_signal_1823, AdderIns_p3[16]}), .b ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, new_AGEMA_signal_1835, AdderIns_p3[20]}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, AdderIns_p4[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_17_a2_U1 ( .a ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, AdderIns_p3[17]}), .b ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, new_AGEMA_signal_1838, AdderIns_p3[21]}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, AdderIns_p4[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_18_a2_U1 ( .a ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, new_AGEMA_signal_1829, AdderIns_p3[18]}), .b ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, new_AGEMA_signal_1841, AdderIns_p3[22]}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, new_AGEMA_signal_2009, AdderIns_p4[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_19_a2_U1 ( .a ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, new_AGEMA_signal_1832, AdderIns_p3[19]}), .b ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, new_AGEMA_signal_1844, AdderIns_p3[23]}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, AdderIns_p4[19]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_20_a2_U1 ( .a ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, new_AGEMA_signal_1835, AdderIns_p3[20]}), .b ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1847, AdderIns_p3[24]}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2015, AdderIns_p4[20]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_21_a2_U1 ( .a ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, new_AGEMA_signal_1838, AdderIns_p3[21]}), .b ({new_AGEMA_signal_1852, new_AGEMA_signal_1851, new_AGEMA_signal_1850, AdderIns_p3[25]}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_2020, new_AGEMA_signal_2019, new_AGEMA_signal_2018, AdderIns_p4[21]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_22_a2_U1 ( .a ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, new_AGEMA_signal_1841, AdderIns_p3[22]}), .b ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, new_AGEMA_signal_1853, AdderIns_p3[26]}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, AdderIns_p4[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_23_a2_U1 ( .a ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, new_AGEMA_signal_1844, AdderIns_p3[23]}), .b ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, new_AGEMA_signal_1856, AdderIns_p3[27]}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2024, AdderIns_p4[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U29 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, new_AGEMA_signal_2285, AdderIns_g6[6]}), .b ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, AdderIns_p6[7]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, sum[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U28 ( .a ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, AdderIns_g6[5]}), .b ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, new_AGEMA_signal_1265, AdderIns_p6[6]}), .c ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, new_AGEMA_signal_2378, sum[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U27 ( .a ({new_AGEMA_signal_2188, new_AGEMA_signal_2187, new_AGEMA_signal_2186, AdderIns_g6[4]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, new_AGEMA_signal_1256, AdderIns_p6[5]}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, sum[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U26 ( .a ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, AdderIns_g6[3]}), .b ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, new_AGEMA_signal_1247, AdderIns_p6[4]}), .c ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, new_AGEMA_signal_2384, sum[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_15_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, sum[7]}), .a ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, new_AGEMA_signal_1211, sum[0]}), .c ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, new_AGEMA_signal_2570, sum_rotated01[15]}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) U130 ( .a ({1'b0, 1'b0, 1'b0, round_constant[10]}), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, sum[10]}), .c ({x_round_out_s3[10], x_round_out_s2[10], x_round_out_s1[10], x_round_out_s0[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U131 ( .a ({1'b0, 1'b0, 1'b0, round_constant[11]}), .b ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, new_AGEMA_signal_2564, sum[11]}), .c ({x_round_out_s3[11], x_round_out_s2[11], x_round_out_s1[11], x_round_out_s0[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U132 ( .a ({1'b0, 1'b0, 1'b0, round_constant[12]}), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, new_AGEMA_signal_2561, sum[12]}), .c ({x_round_out_s3[12], x_round_out_s2[12], x_round_out_s1[12], x_round_out_s0[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U133 ( .a ({1'b0, 1'b0, 1'b0, round_constant[13]}), .b ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, sum[13]}), .c ({x_round_out_s3[13], x_round_out_s2[13], x_round_out_s1[13], x_round_out_s0[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U134 ( .a ({1'b0, 1'b0, 1'b0, round_constant[14]}), .b ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, new_AGEMA_signal_2555, sum[14]}), .c ({x_round_out_s3[14], x_round_out_s2[14], x_round_out_s1[14], x_round_out_s0[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U135 ( .a ({1'b0, 1'b0, 1'b0, round_constant[15]}), .b ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, new_AGEMA_signal_2642, sum[15]}), .c ({x_round_out_s3[15], x_round_out_s2[15], x_round_out_s1[15], x_round_out_s0[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U159 ( .a ({1'b0, 1'b0, 1'b0, round_constant[8]}), .b ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, new_AGEMA_signal_2552, sum[8]}), .c ({x_round_out_s3[8], x_round_out_s2[8], x_round_out_s1[8], x_round_out_s0[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U160 ( .a ({1'b0, 1'b0, 1'b0, round_constant[9]}), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, new_AGEMA_signal_2549, sum[9]}), .c ({x_round_out_s3[9], x_round_out_s2[9], x_round_out_s1[9], x_round_out_s0[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U168 ( .a ({new_AGEMA_signal_2920, new_AGEMA_signal_2919, new_AGEMA_signal_2918, sum_rotated[16]}), .b ({y_round_in_s3[16], y_round_in_s2[16], y_round_in_s1[16], y_round_in_s0[16]}), .c ({y_round_out_s3[16], y_round_out_s2[16], y_round_out_s1[16], y_round_out_s0[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_0_a1_U1 ( .a ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, AdderIns_g3[7]}), .b ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, new_AGEMA_signal_2195, AdderIns_s4_bc_0_a1_t}), .c ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, new_AGEMA_signal_2288, AdderIns_g4[7]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_2038, new_AGEMA_signal_2037, new_AGEMA_signal_2036, AdderIns_g3[3]}), .b ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, new_AGEMA_signal_1787, AdderIns_p3[4]}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, new_AGEMA_signal_2195, AdderIns_s4_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_1_a1_U1 ( .a ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, new_AGEMA_signal_2051, AdderIns_g3[8]}), .b ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, new_AGEMA_signal_2198, AdderIns_s4_bc_1_a1_t}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, new_AGEMA_signal_2291, AdderIns_g4[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, AdderIns_g3[4]}), .b ({new_AGEMA_signal_1792, new_AGEMA_signal_1791, new_AGEMA_signal_1790, AdderIns_p3[5]}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, new_AGEMA_signal_2198, AdderIns_s4_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_2_a1_U1 ( .a ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, AdderIns_g3[9]}), .b ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, new_AGEMA_signal_2201, AdderIns_s4_bc_2_a1_t}), .c ({new_AGEMA_signal_2296, new_AGEMA_signal_2295, new_AGEMA_signal_2294, AdderIns_g4[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, AdderIns_g3[5]}), .b ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, new_AGEMA_signal_1793, AdderIns_p3[6]}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, new_AGEMA_signal_2201, AdderIns_s4_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_3_a1_U1 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, new_AGEMA_signal_2057, AdderIns_g3[10]}), .b ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, new_AGEMA_signal_2204, AdderIns_s4_bc_3_a1_t}), .c ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, new_AGEMA_signal_2297, AdderIns_g4[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, new_AGEMA_signal_2045, AdderIns_g3[6]}), .b ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, new_AGEMA_signal_1796, AdderIns_p3[7]}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, new_AGEMA_signal_2204, AdderIns_s4_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_4_a1_U1 ( .a ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, new_AGEMA_signal_2060, AdderIns_g3[11]}), .b ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, new_AGEMA_signal_2207, AdderIns_s4_bc_4_a1_t}), .c ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, new_AGEMA_signal_2300, AdderIns_g4[11]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, AdderIns_g3[7]}), .b ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, new_AGEMA_signal_1799, AdderIns_p3[8]}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, new_AGEMA_signal_2207, AdderIns_s4_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_5_a1_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, AdderIns_g3[12]}), .b ({new_AGEMA_signal_2212, new_AGEMA_signal_2211, new_AGEMA_signal_2210, AdderIns_s4_bc_5_a1_t}), .c ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, new_AGEMA_signal_2303, AdderIns_g4[12]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, new_AGEMA_signal_2051, AdderIns_g3[8]}), .b ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, new_AGEMA_signal_1802, AdderIns_p3[9]}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_2212, new_AGEMA_signal_2211, new_AGEMA_signal_2210, AdderIns_s4_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_6_a1_U1 ( .a ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, AdderIns_g3[13]}), .b ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, new_AGEMA_signal_2213, AdderIns_s4_bc_6_a1_t}), .c ({new_AGEMA_signal_2308, new_AGEMA_signal_2307, new_AGEMA_signal_2306, AdderIns_g4[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, AdderIns_g3[9]}), .b ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, new_AGEMA_signal_1805, AdderIns_p3[10]}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, new_AGEMA_signal_2213, AdderIns_s4_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_7_a1_U1 ( .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, AdderIns_g3[14]}), .b ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, new_AGEMA_signal_2216, AdderIns_s4_bc_7_a1_t}), .c ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, new_AGEMA_signal_2309, AdderIns_g4[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, new_AGEMA_signal_2057, AdderIns_g3[10]}), .b ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, new_AGEMA_signal_1808, AdderIns_p3[11]}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, new_AGEMA_signal_2216, AdderIns_s4_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_8_a1_U1 ( .a ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, AdderIns_g3[15]}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, new_AGEMA_signal_2219, AdderIns_s4_bc_8_a1_t}), .c ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, new_AGEMA_signal_2312, AdderIns_g4[15]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, new_AGEMA_signal_2060, AdderIns_g3[11]}), .b ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, new_AGEMA_signal_1811, AdderIns_p3[12]}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, new_AGEMA_signal_2219, AdderIns_s4_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_9_a1_U1 ( .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, new_AGEMA_signal_2075, AdderIns_g3[16]}), .b ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, AdderIns_s4_bc_9_a1_t}), .c ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, new_AGEMA_signal_2315, AdderIns_g4[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, AdderIns_g3[12]}), .b ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, new_AGEMA_signal_1814, AdderIns_p3[13]}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, AdderIns_s4_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_10_a1_U1 ( .a ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, AdderIns_g3[17]}), .b ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, new_AGEMA_signal_2225, AdderIns_s4_bc_10_a1_t}), .c ({new_AGEMA_signal_2320, new_AGEMA_signal_2319, new_AGEMA_signal_2318, AdderIns_g4[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, AdderIns_g3[13]}), .b ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, new_AGEMA_signal_1817, AdderIns_p3[14]}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, new_AGEMA_signal_2225, AdderIns_s4_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_11_a1_U1 ( .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, new_AGEMA_signal_2081, AdderIns_g3[18]}), .b ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, new_AGEMA_signal_2228, AdderIns_s4_bc_11_a1_t}), .c ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, new_AGEMA_signal_2321, AdderIns_g4[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, AdderIns_g3[14]}), .b ({new_AGEMA_signal_1822, new_AGEMA_signal_1821, new_AGEMA_signal_1820, AdderIns_p3[15]}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, new_AGEMA_signal_2228, AdderIns_s4_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_12_a1_U1 ( .a ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, AdderIns_g3[19]}), .b ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, new_AGEMA_signal_2231, AdderIns_s4_bc_12_a1_t}), .c ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, new_AGEMA_signal_2324, AdderIns_g4[19]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, AdderIns_g3[15]}), .b ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, new_AGEMA_signal_1823, AdderIns_p3[16]}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, new_AGEMA_signal_2231, AdderIns_s4_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_13_a1_U1 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, AdderIns_g3[20]}), .b ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, AdderIns_s4_bc_13_a1_t}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, AdderIns_g4[20]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, new_AGEMA_signal_2075, AdderIns_g3[16]}), .b ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1826, AdderIns_p3[17]}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, AdderIns_s4_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_14_a1_U1 ( .a ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, AdderIns_g3[21]}), .b ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, new_AGEMA_signal_2237, AdderIns_s4_bc_14_a1_t}), .c ({new_AGEMA_signal_2332, new_AGEMA_signal_2331, new_AGEMA_signal_2330, AdderIns_g4[21]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, AdderIns_g3[17]}), .b ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, new_AGEMA_signal_1829, AdderIns_p3[18]}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, new_AGEMA_signal_2237, AdderIns_s4_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_15_a1_U1 ( .a ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, AdderIns_g3[22]}), .b ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, new_AGEMA_signal_2240, AdderIns_s4_bc_15_a1_t}), .c ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, new_AGEMA_signal_2333, AdderIns_g4[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, new_AGEMA_signal_2081, AdderIns_g3[18]}), .b ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, new_AGEMA_signal_1832, AdderIns_p3[19]}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, new_AGEMA_signal_2240, AdderIns_s4_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_16_a1_U1 ( .a ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, new_AGEMA_signal_2096, AdderIns_g3[23]}), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, AdderIns_s4_bc_16_a1_t}), .c ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, new_AGEMA_signal_2336, AdderIns_g4[23]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_16_a1_a1_U1 ( .a ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, AdderIns_g3[19]}), .b ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, new_AGEMA_signal_1835, AdderIns_p3[20]}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, AdderIns_s4_bc_16_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_17_a1_U1 ( .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, AdderIns_g3[24]}), .b ({new_AGEMA_signal_2248, new_AGEMA_signal_2247, new_AGEMA_signal_2246, AdderIns_s4_bc_17_a1_t}), .c ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, new_AGEMA_signal_2339, AdderIns_g4[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_17_a1_a1_U1 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, AdderIns_g3[20]}), .b ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, new_AGEMA_signal_1838, AdderIns_p3[21]}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_2248, new_AGEMA_signal_2247, new_AGEMA_signal_2246, AdderIns_s4_bc_17_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_18_a1_U1 ( .a ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, AdderIns_g3[25]}), .b ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, new_AGEMA_signal_2249, AdderIns_s4_bc_18_a1_t}), .c ({new_AGEMA_signal_2344, new_AGEMA_signal_2343, new_AGEMA_signal_2342, AdderIns_g4[25]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_18_a1_a1_U1 ( .a ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, AdderIns_g3[21]}), .b ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, new_AGEMA_signal_1841, AdderIns_p3[22]}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, new_AGEMA_signal_2249, AdderIns_s4_bc_18_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_19_a1_U1 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, new_AGEMA_signal_2105, AdderIns_g3[26]}), .b ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, new_AGEMA_signal_2252, AdderIns_s4_bc_19_a1_t}), .c ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, new_AGEMA_signal_2345, AdderIns_g4[26]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_19_a1_a1_U1 ( .a ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, AdderIns_g3[22]}), .b ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, new_AGEMA_signal_1844, AdderIns_p3[23]}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, new_AGEMA_signal_2252, AdderIns_s4_bc_19_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_20_a1_U1 ( .a ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, AdderIns_g3[27]}), .b ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, new_AGEMA_signal_2255, AdderIns_s4_bc_20_a1_t}), .c ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, new_AGEMA_signal_2348, AdderIns_g4[27]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_20_a1_a1_U1 ( .a ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, new_AGEMA_signal_2096, AdderIns_g3[23]}), .b ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1847, AdderIns_p3[24]}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, new_AGEMA_signal_2255, AdderIns_s4_bc_20_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_21_a1_U1 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, new_AGEMA_signal_2111, AdderIns_g3[28]}), .b ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, AdderIns_s4_bc_21_a1_t}), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, new_AGEMA_signal_2351, AdderIns_g4[28]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_21_a1_a1_U1 ( .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, AdderIns_g3[24]}), .b ({new_AGEMA_signal_1852, new_AGEMA_signal_1851, new_AGEMA_signal_1850, AdderIns_p3[25]}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, AdderIns_s4_bc_21_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_22_a1_U1 ( .a ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, new_AGEMA_signal_2114, AdderIns_g3[29]}), .b ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, new_AGEMA_signal_2261, AdderIns_s4_bc_22_a1_t}), .c ({new_AGEMA_signal_2356, new_AGEMA_signal_2355, new_AGEMA_signal_2354, AdderIns_g4[29]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_22_a1_a1_U1 ( .a ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, AdderIns_g3[25]}), .b ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, new_AGEMA_signal_1853, AdderIns_p3[26]}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, new_AGEMA_signal_2261, AdderIns_s4_bc_22_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_23_a1_U1 ( .a ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, new_AGEMA_signal_2117, AdderIns_g3[30]}), .b ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, new_AGEMA_signal_2264, AdderIns_s4_bc_23_a1_t}), .c ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, new_AGEMA_signal_2357, AdderIns_g4[30]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s4_bc_23_a1_a1_U1 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, new_AGEMA_signal_2105, AdderIns_g3[26]}), .b ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, new_AGEMA_signal_1856, AdderIns_p3[27]}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, new_AGEMA_signal_2264, AdderIns_s4_bc_23_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_0_a1_U1 ( .a ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, new_AGEMA_signal_2288, AdderIns_g4[7]}), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, new_AGEMA_signal_2123, AdderIns_s5_gc_0_a1_t}), .c ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, new_AGEMA_signal_2396, AdderIns_g6[7]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_0_a1_a1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, new_AGEMA_signal_1955, AdderIns_p4[0]}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, new_AGEMA_signal_2123, AdderIns_s5_gc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_1_a1_U1 ( .a ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, new_AGEMA_signal_2291, AdderIns_g4[8]}), .b ({new_AGEMA_signal_2128, new_AGEMA_signal_2127, new_AGEMA_signal_2126, AdderIns_s5_gc_1_a1_t}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, AdderIns_g6[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, AdderIns_g6[0]}), .b ({new_AGEMA_signal_1960, new_AGEMA_signal_1959, new_AGEMA_signal_1958, AdderIns_p4[1]}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_2128, new_AGEMA_signal_2127, new_AGEMA_signal_2126, AdderIns_s5_gc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_2_a1_U1 ( .a ({new_AGEMA_signal_2296, new_AGEMA_signal_2295, new_AGEMA_signal_2294, AdderIns_g4[9]}), .b ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, new_AGEMA_signal_2129, AdderIns_s5_gc_2_a1_t}), .c ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, new_AGEMA_signal_2402, AdderIns_g6[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, new_AGEMA_signal_1859, AdderIns_g6[1]}), .b ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, new_AGEMA_signal_1961, AdderIns_p4[2]}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, new_AGEMA_signal_2129, AdderIns_s5_gc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_3_a1_U1 ( .a ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, new_AGEMA_signal_2297, AdderIns_g4[10]}), .b ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, new_AGEMA_signal_2267, AdderIns_s5_gc_3_a1_t}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, new_AGEMA_signal_2405, AdderIns_g6[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, AdderIns_g6[2]}), .b ({new_AGEMA_signal_1966, new_AGEMA_signal_1965, new_AGEMA_signal_1964, AdderIns_p4[3]}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, new_AGEMA_signal_2267, AdderIns_s5_gc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_4_a1_U1 ( .a ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, new_AGEMA_signal_2300, AdderIns_g4[11]}), .b ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, new_AGEMA_signal_2360, AdderIns_s5_gc_4_a1_t}), .c ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, new_AGEMA_signal_2408, AdderIns_g6[11]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, AdderIns_g6[3]}), .b ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, new_AGEMA_signal_1967, AdderIns_p4[4]}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, new_AGEMA_signal_2360, AdderIns_s5_gc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_5_a1_U1 ( .a ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, new_AGEMA_signal_2303, AdderIns_g4[12]}), .b ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, new_AGEMA_signal_2363, AdderIns_s5_gc_5_a1_t}), .c ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, new_AGEMA_signal_2411, AdderIns_g6[12]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_2188, new_AGEMA_signal_2187, new_AGEMA_signal_2186, AdderIns_g6[4]}), .b ({new_AGEMA_signal_1972, new_AGEMA_signal_1971, new_AGEMA_signal_1970, AdderIns_p4[5]}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, new_AGEMA_signal_2363, AdderIns_s5_gc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_6_a1_U1 ( .a ({new_AGEMA_signal_2308, new_AGEMA_signal_2307, new_AGEMA_signal_2306, AdderIns_g4[13]}), .b ({new_AGEMA_signal_2368, new_AGEMA_signal_2367, new_AGEMA_signal_2366, AdderIns_s5_gc_6_a1_t}), .c ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, new_AGEMA_signal_2414, AdderIns_g6[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, AdderIns_g6[5]}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, new_AGEMA_signal_1973, AdderIns_p4[6]}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_2368, new_AGEMA_signal_2367, new_AGEMA_signal_2366, AdderIns_s5_gc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_7_a1_U1 ( .a ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, new_AGEMA_signal_2309, AdderIns_g4[14]}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, new_AGEMA_signal_2417, AdderIns_s5_gc_7_a1_t}), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, new_AGEMA_signal_2477, AdderIns_g6[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_gc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, new_AGEMA_signal_2285, AdderIns_g6[6]}), .b ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, new_AGEMA_signal_1976, AdderIns_p4[7]}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, new_AGEMA_signal_2417, AdderIns_s5_gc_7_a1_t}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_1_a2_U1 ( .a ({new_AGEMA_signal_1960, new_AGEMA_signal_1959, new_AGEMA_signal_1958, AdderIns_p4[1]}), .b ({new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1982, AdderIns_p4[9]}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, new_AGEMA_signal_2132, AdderIns_p5[1]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_2_a2_U1 ( .a ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, new_AGEMA_signal_1961, AdderIns_p4[2]}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, AdderIns_p4[10]}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, new_AGEMA_signal_2135, AdderIns_p5[2]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_3_a2_U1 ( .a ({new_AGEMA_signal_1966, new_AGEMA_signal_1965, new_AGEMA_signal_1964, AdderIns_p4[3]}), .b ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, new_AGEMA_signal_1988, AdderIns_p4[11]}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, new_AGEMA_signal_2138, AdderIns_p5[3]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_4_a2_U1 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, new_AGEMA_signal_1967, AdderIns_p4[4]}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1991, AdderIns_p4[12]}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, new_AGEMA_signal_2141, AdderIns_p5[4]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_5_a2_U1 ( .a ({new_AGEMA_signal_1972, new_AGEMA_signal_1971, new_AGEMA_signal_1970, AdderIns_p4[5]}), .b ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, AdderIns_p4[13]}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, AdderIns_p5[5]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_6_a2_U1 ( .a ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, new_AGEMA_signal_1973, AdderIns_p4[6]}), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, new_AGEMA_signal_1997, AdderIns_p4[14]}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, new_AGEMA_signal_2147, AdderIns_p5[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_7_a2_U1 ( .a ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, new_AGEMA_signal_1976, AdderIns_p4[7]}), .b ({new_AGEMA_signal_2002, new_AGEMA_signal_2001, new_AGEMA_signal_2000, AdderIns_p4[15]}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_2152, new_AGEMA_signal_2151, new_AGEMA_signal_2150, AdderIns_p5[7]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_8_a2_U1 ( .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, new_AGEMA_signal_1979, AdderIns_p4[8]}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, AdderIns_p4[16]}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, AdderIns_p5[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_9_a2_U1 ( .a ({new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1982, AdderIns_p4[9]}), .b ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, AdderIns_p4[17]}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, new_AGEMA_signal_2156, AdderIns_p5[9]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_10_a2_U1 ( .a ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, AdderIns_p4[10]}), .b ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, new_AGEMA_signal_2009, AdderIns_p4[18]}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, new_AGEMA_signal_2159, AdderIns_p5[10]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_11_a2_U1 ( .a ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, new_AGEMA_signal_1988, AdderIns_p4[11]}), .b ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, AdderIns_p4[19]}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, AdderIns_p5[11]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_12_a2_U1 ( .a ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1991, AdderIns_p4[12]}), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2015, AdderIns_p4[20]}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, new_AGEMA_signal_2165, AdderIns_p5[12]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_13_a2_U1 ( .a ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, AdderIns_p4[13]}), .b ({new_AGEMA_signal_2020, new_AGEMA_signal_2019, new_AGEMA_signal_2018, AdderIns_p4[21]}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, new_AGEMA_signal_2168, AdderIns_p5[13]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_14_a2_U1 ( .a ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, new_AGEMA_signal_1997, AdderIns_p4[14]}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, AdderIns_p4[22]}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, new_AGEMA_signal_2171, AdderIns_p5[14]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_15_a2_U1 ( .a ({new_AGEMA_signal_2002, new_AGEMA_signal_2001, new_AGEMA_signal_2000, AdderIns_p4[15]}), .b ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2024, AdderIns_p4[23]}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, AdderIns_p5[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U31 ( .a ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, AdderIns_g6[8]}), .b ({new_AGEMA_signal_1294, new_AGEMA_signal_1293, new_AGEMA_signal_1292, AdderIns_p6[9]}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, new_AGEMA_signal_2549, sum[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U30 ( .a ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, new_AGEMA_signal_2396, AdderIns_g6[7]}), .b ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, new_AGEMA_signal_1283, AdderIns_p6[8]}), .c ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, new_AGEMA_signal_2552, sum[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U6 ( .a ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, new_AGEMA_signal_2477, AdderIns_g6[14]}), .b ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, AdderIns_p6[15]}), .c ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, new_AGEMA_signal_2642, sum[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U5 ( .a ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, new_AGEMA_signal_2414, AdderIns_g6[13]}), .b ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, new_AGEMA_signal_1337, AdderIns_p6[14]}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, new_AGEMA_signal_2555, sum[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U4 ( .a ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, new_AGEMA_signal_2411, AdderIns_g6[12]}), .b ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, new_AGEMA_signal_1328, AdderIns_p6[13]}), .c ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, sum[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U3 ( .a ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, new_AGEMA_signal_2408, AdderIns_g6[11]}), .b ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, new_AGEMA_signal_1319, AdderIns_p6[12]}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, new_AGEMA_signal_2561, sum[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U2 ( .a ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, new_AGEMA_signal_2405, AdderIns_g6[10]}), .b ({new_AGEMA_signal_1312, new_AGEMA_signal_1311, new_AGEMA_signal_1310, AdderIns_p6[11]}), .c ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, new_AGEMA_signal_2564, sum[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U1 ( .a ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, new_AGEMA_signal_2402, AdderIns_g6[9]}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, new_AGEMA_signal_1301, AdderIns_p6[10]}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, sum[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_16_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, new_AGEMA_signal_2552, sum[8]}), .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, new_AGEMA_signal_2027, sum[1]}), .c ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, new_AGEMA_signal_2645, sum_rotated01[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_17_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, new_AGEMA_signal_2549, sum[9]}), .a ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, sum[2]}), .c ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, new_AGEMA_signal_2648, sum_rotated01[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_18_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, sum[10]}), .a ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, sum[3]}), .c ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, new_AGEMA_signal_2651, sum_rotated01[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_19_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, new_AGEMA_signal_2564, sum[11]}), .a ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, new_AGEMA_signal_2384, sum[4]}), .c ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, new_AGEMA_signal_2654, sum_rotated01[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_20_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, new_AGEMA_signal_2561, sum[12]}), .a ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, sum[5]}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, new_AGEMA_signal_2657, sum_rotated01[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_21_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, sum[13]}), .a ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, new_AGEMA_signal_2378, sum[6]}), .c ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, new_AGEMA_signal_2660, sum_rotated01[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_22_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, new_AGEMA_signal_2555, sum[14]}), .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, sum[7]}), .c ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, new_AGEMA_signal_2663, sum_rotated01[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_23_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, new_AGEMA_signal_2642, sum[15]}), .a ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, new_AGEMA_signal_2552, sum[8]}), .c ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, new_AGEMA_signal_2717, sum_rotated01[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_16_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, new_AGEMA_signal_2642, sum[15]}), .a ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, new_AGEMA_signal_1211, sum[0]}), .c ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, new_AGEMA_signal_2723, sum_rotated23[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_16_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, new_AGEMA_signal_2645, sum_rotated01[16]}), .a ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, new_AGEMA_signal_2723, sum_rotated23[16]}), .c ({new_AGEMA_signal_2920, new_AGEMA_signal_2919, new_AGEMA_signal_2918, sum_rotated[16]}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) U136 ( .a ({1'b0, 1'b0, 1'b0, round_constant[16]}), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, sum[16]}), .c ({x_round_out_s3[16], x_round_out_s2[16], x_round_out_s1[16], x_round_out_s0[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U137 ( .a ({1'b0, 1'b0, 1'b0, round_constant[17]}), .b ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, sum[17]}), .c ({x_round_out_s3[17], x_round_out_s2[17], x_round_out_s1[17], x_round_out_s0[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U138 ( .a ({1'b0, 1'b0, 1'b0, round_constant[18]}), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, sum[18]}), .c ({x_round_out_s3[18], x_round_out_s2[18], x_round_out_s1[18], x_round_out_s0[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U139 ( .a ({1'b0, 1'b0, 1'b0, round_constant[19]}), .b ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, sum[19]}), .c ({x_round_out_s3[19], x_round_out_s2[19], x_round_out_s1[19], x_round_out_s0[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U141 ( .a ({1'b0, 1'b0, 1'b0, round_constant[20]}), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, new_AGEMA_signal_2705, sum[20]}), .c ({x_round_out_s3[20], x_round_out_s2[20], x_round_out_s1[20], x_round_out_s0[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U142 ( .a ({1'b0, 1'b0, 1'b0, round_constant[21]}), .b ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, sum[21]}), .c ({x_round_out_s3[21], x_round_out_s2[21], x_round_out_s1[21], x_round_out_s0[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U143 ( .a ({1'b0, 1'b0, 1'b0, round_constant[22]}), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, sum[22]}), .c ({x_round_out_s3[22], x_round_out_s2[22], x_round_out_s1[22], x_round_out_s0[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U144 ( .a ({1'b0, 1'b0, 1'b0, round_constant[23]}), .b ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, new_AGEMA_signal_2696, sum[23]}), .c ({x_round_out_s3[23], x_round_out_s2[23], x_round_out_s1[23], x_round_out_s0[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U145 ( .a ({1'b0, 1'b0, 1'b0, round_constant[24]}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, sum[24]}), .c ({x_round_out_s3[24], x_round_out_s2[24], x_round_out_s1[24], x_round_out_s0[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U146 ( .a ({1'b0, 1'b0, 1'b0, round_constant[25]}), .b ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, sum[25]}), .c ({x_round_out_s3[25], x_round_out_s2[25], x_round_out_s1[25], x_round_out_s0[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U147 ( .a ({1'b0, 1'b0, 1'b0, round_constant[26]}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2687, sum[26]}), .c ({x_round_out_s3[26], x_round_out_s2[26], x_round_out_s1[26], x_round_out_s0[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U148 ( .a ({1'b0, 1'b0, 1'b0, round_constant[27]}), .b ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, sum[27]}), .c ({x_round_out_s3[27], x_round_out_s2[27], x_round_out_s1[27], x_round_out_s0[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U149 ( .a ({1'b0, 1'b0, 1'b0, round_constant[28]}), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, new_AGEMA_signal_2681, sum[28]}), .c ({x_round_out_s3[28], x_round_out_s2[28], x_round_out_s1[28], x_round_out_s0[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U150 ( .a ({1'b0, 1'b0, 1'b0, round_constant[29]}), .b ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, new_AGEMA_signal_2678, sum[29]}), .c ({x_round_out_s3[29], x_round_out_s2[29], x_round_out_s1[29], x_round_out_s0[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U152 ( .a ({1'b0, 1'b0, 1'b0, round_constant[30]}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, sum[30]}), .c ({x_round_out_s3[30], x_round_out_s2[30], x_round_out_s1[30], x_round_out_s0[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U153 ( .a ({1'b0, 1'b0, 1'b0, round_constant[31]}), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2771, sum[31]}), .c ({x_round_out_s3[31], x_round_out_s2[31], x_round_out_s1[31], x_round_out_s0[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U161 ( .a ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, new_AGEMA_signal_3101, sum_rotated[0]}), .b ({y_round_in_s3[0], y_round_in_s2[0], y_round_in_s1[0], y_round_in_s0[0]}), .c ({y_round_out_s3[0], y_round_out_s2[0], y_round_out_s1[0], y_round_out_s0[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U162 ( .a ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, new_AGEMA_signal_2969, sum_rotated[10]}), .b ({y_round_in_s3[10], y_round_in_s2[10], y_round_in_s1[10], y_round_in_s0[10]}), .c ({y_round_out_s3[10], y_round_out_s2[10], y_round_out_s1[10], y_round_out_s0[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U163 ( .a ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, new_AGEMA_signal_2972, sum_rotated[11]}), .b ({y_round_in_s3[11], y_round_in_s2[11], y_round_in_s1[11], y_round_in_s0[11]}), .c ({y_round_out_s3[11], y_round_out_s2[11], y_round_out_s1[11], y_round_out_s0[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U164 ( .a ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, new_AGEMA_signal_2975, sum_rotated[12]}), .b ({y_round_in_s3[12], y_round_in_s2[12], y_round_in_s1[12], y_round_in_s0[12]}), .c ({y_round_out_s3[12], y_round_out_s2[12], y_round_out_s1[12], y_round_out_s0[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U165 ( .a ({new_AGEMA_signal_2980, new_AGEMA_signal_2979, new_AGEMA_signal_2978, sum_rotated[13]}), .b ({y_round_in_s3[13], y_round_in_s2[13], y_round_in_s1[13], y_round_in_s0[13]}), .c ({y_round_out_s3[13], y_round_out_s2[13], y_round_out_s1[13], y_round_out_s0[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U166 ( .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3107, sum_rotated[14]}), .b ({y_round_in_s3[14], y_round_in_s2[14], y_round_in_s1[14], y_round_in_s0[14]}), .c ({y_round_out_s3[14], y_round_out_s2[14], y_round_out_s1[14], y_round_out_s0[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U167 ( .a ({new_AGEMA_signal_3112, new_AGEMA_signal_3111, new_AGEMA_signal_3110, sum_rotated[15]}), .b ({y_round_in_s3[15], y_round_in_s2[15], y_round_in_s1[15], y_round_in_s0[15]}), .c ({y_round_out_s3[15], y_round_out_s2[15], y_round_out_s1[15], y_round_out_s0[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U169 ( .a ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, new_AGEMA_signal_2921, sum_rotated[17]}), .b ({y_round_in_s3[17], y_round_in_s2[17], y_round_in_s1[17], y_round_in_s0[17]}), .c ({y_round_out_s3[17], y_round_out_s2[17], y_round_out_s1[17], y_round_out_s0[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U170 ( .a ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, new_AGEMA_signal_2981, sum_rotated[18]}), .b ({y_round_in_s3[18], y_round_in_s2[18], y_round_in_s1[18], y_round_in_s0[18]}), .c ({y_round_out_s3[18], y_round_out_s2[18], y_round_out_s1[18], y_round_out_s0[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U171 ( .a ({new_AGEMA_signal_2986, new_AGEMA_signal_2985, new_AGEMA_signal_2984, sum_rotated[19]}), .b ({y_round_in_s3[19], y_round_in_s2[19], y_round_in_s1[19], y_round_in_s0[19]}), .c ({y_round_out_s3[19], y_round_out_s2[19], y_round_out_s1[19], y_round_out_s0[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U172 ( .a ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, new_AGEMA_signal_2945, sum_rotated[1]}), .b ({y_round_in_s3[1], y_round_in_s2[1], y_round_in_s1[1], y_round_in_s0[1]}), .c ({y_round_out_s3[1], y_round_out_s2[1], y_round_out_s1[1], y_round_out_s0[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U173 ( .a ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, new_AGEMA_signal_2987, sum_rotated[20]}), .b ({y_round_in_s3[20], y_round_in_s2[20], y_round_in_s1[20], y_round_in_s0[20]}), .c ({y_round_out_s3[20], y_round_out_s2[20], y_round_out_s1[20], y_round_out_s0[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U174 ( .a ({new_AGEMA_signal_2992, new_AGEMA_signal_2991, new_AGEMA_signal_2990, sum_rotated[21]}), .b ({y_round_in_s3[21], y_round_in_s2[21], y_round_in_s1[21], y_round_in_s0[21]}), .c ({y_round_out_s3[21], y_round_out_s2[21], y_round_out_s1[21], y_round_out_s0[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U175 ( .a ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, new_AGEMA_signal_2993, sum_rotated[22]}), .b ({y_round_in_s3[22], y_round_in_s2[22], y_round_in_s1[22], y_round_in_s0[22]}), .c ({y_round_out_s3[22], y_round_out_s2[22], y_round_out_s1[22], y_round_out_s0[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U176 ( .a ({new_AGEMA_signal_2998, new_AGEMA_signal_2997, new_AGEMA_signal_2996, sum_rotated[23]}), .b ({y_round_in_s3[23], y_round_in_s2[23], y_round_in_s1[23], y_round_in_s0[23]}), .c ({y_round_out_s3[23], y_round_out_s2[23], y_round_out_s1[23], y_round_out_s0[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U177 ( .a ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, new_AGEMA_signal_2999, sum_rotated[24]}), .b ({y_round_in_s3[24], y_round_in_s2[24], y_round_in_s1[24], y_round_in_s0[24]}), .c ({y_round_out_s3[24], y_round_out_s2[24], y_round_out_s1[24], y_round_out_s0[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U178 ( .a ({new_AGEMA_signal_3004, new_AGEMA_signal_3003, new_AGEMA_signal_3002, sum_rotated[25]}), .b ({y_round_in_s3[25], y_round_in_s2[25], y_round_in_s1[25], y_round_in_s0[25]}), .c ({y_round_out_s3[25], y_round_out_s2[25], y_round_out_s1[25], y_round_out_s0[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U179 ( .a ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, new_AGEMA_signal_3005, sum_rotated[26]}), .b ({y_round_in_s3[26], y_round_in_s2[26], y_round_in_s1[26], y_round_in_s0[26]}), .c ({y_round_out_s3[26], y_round_out_s2[26], y_round_out_s1[26], y_round_out_s0[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U180 ( .a ({new_AGEMA_signal_3010, new_AGEMA_signal_3009, new_AGEMA_signal_3008, sum_rotated[27]}), .b ({y_round_in_s3[27], y_round_in_s2[27], y_round_in_s1[27], y_round_in_s0[27]}), .c ({y_round_out_s3[27], y_round_out_s2[27], y_round_out_s1[27], y_round_out_s0[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U181 ( .a ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, new_AGEMA_signal_3011, sum_rotated[28]}), .b ({y_round_in_s3[28], y_round_in_s2[28], y_round_in_s1[28], y_round_in_s0[28]}), .c ({y_round_out_s3[28], y_round_out_s2[28], y_round_out_s1[28], y_round_out_s0[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U182 ( .a ({new_AGEMA_signal_3016, new_AGEMA_signal_3015, new_AGEMA_signal_3014, sum_rotated[29]}), .b ({y_round_in_s3[29], y_round_in_s2[29], y_round_in_s1[29], y_round_in_s0[29]}), .c ({y_round_out_s3[29], y_round_out_s2[29], y_round_out_s1[29], y_round_out_s0[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U183 ( .a ({new_AGEMA_signal_2950, new_AGEMA_signal_2949, new_AGEMA_signal_2948, sum_rotated[2]}), .b ({y_round_in_s3[2], y_round_in_s2[2], y_round_in_s1[2], y_round_in_s0[2]}), .c ({y_round_out_s3[2], y_round_out_s2[2], y_round_out_s1[2], y_round_out_s0[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U184 ( .a ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, new_AGEMA_signal_3017, sum_rotated[30]}), .b ({y_round_in_s3[30], y_round_in_s2[30], y_round_in_s1[30], y_round_in_s0[30]}), .c ({y_round_out_s3[30], y_round_out_s2[30], y_round_out_s1[30], y_round_out_s0[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U185 ( .a ({new_AGEMA_signal_3022, new_AGEMA_signal_3021, new_AGEMA_signal_3020, sum_rotated[31]}), .b ({y_round_in_s3[31], y_round_in_s2[31], y_round_in_s1[31], y_round_in_s0[31]}), .c ({y_round_out_s3[31], y_round_out_s2[31], y_round_out_s1[31], y_round_out_s0[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U186 ( .a ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, new_AGEMA_signal_2951, sum_rotated[3]}), .b ({y_round_in_s3[3], y_round_in_s2[3], y_round_in_s1[3], y_round_in_s0[3]}), .c ({y_round_out_s3[3], y_round_out_s2[3], y_round_out_s1[3], y_round_out_s0[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U187 ( .a ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, new_AGEMA_signal_2954, sum_rotated[4]}), .b ({y_round_in_s3[4], y_round_in_s2[4], y_round_in_s1[4], y_round_in_s0[4]}), .c ({y_round_out_s3[4], y_round_out_s2[4], y_round_out_s1[4], y_round_out_s0[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U188 ( .a ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, new_AGEMA_signal_2957, sum_rotated[5]}), .b ({y_round_in_s3[5], y_round_in_s2[5], y_round_in_s1[5], y_round_in_s0[5]}), .c ({y_round_out_s3[5], y_round_out_s2[5], y_round_out_s1[5], y_round_out_s0[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U189 ( .a ({new_AGEMA_signal_2962, new_AGEMA_signal_2961, new_AGEMA_signal_2960, sum_rotated[6]}), .b ({y_round_in_s3[6], y_round_in_s2[6], y_round_in_s1[6], y_round_in_s0[6]}), .c ({y_round_out_s3[6], y_round_out_s2[6], y_round_out_s1[6], y_round_out_s0[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U190 ( .a ({new_AGEMA_signal_3106, new_AGEMA_signal_3105, new_AGEMA_signal_3104, sum_rotated[7]}), .b ({y_round_in_s3[7], y_round_in_s2[7], y_round_in_s1[7], y_round_in_s0[7]}), .c ({y_round_out_s3[7], y_round_out_s2[7], y_round_out_s1[7], y_round_out_s0[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U191 ( .a ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, new_AGEMA_signal_2963, sum_rotated[8]}), .b ({y_round_in_s3[8], y_round_in_s2[8], y_round_in_s1[8], y_round_in_s0[8]}), .c ({y_round_out_s3[8], y_round_out_s2[8], y_round_out_s1[8], y_round_out_s0[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U192 ( .a ({new_AGEMA_signal_2968, new_AGEMA_signal_2967, new_AGEMA_signal_2966, sum_rotated[9]}), .b ({y_round_in_s3[9], y_round_in_s2[9], y_round_in_s1[9], y_round_in_s0[9]}), .c ({y_round_out_s3[9], y_round_out_s2[9], y_round_out_s1[9], y_round_out_s0[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_0_a1_U1 ( .a ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, new_AGEMA_signal_2312, AdderIns_g4[15]}), .b ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, new_AGEMA_signal_2420, AdderIns_s5_bc_0_a1_t}), .c ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, new_AGEMA_signal_2480, AdderIns_g6[15]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_0_a1_a1_U1 ( .a ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, new_AGEMA_signal_2288, AdderIns_g4[7]}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, new_AGEMA_signal_1979, AdderIns_p4[8]}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, new_AGEMA_signal_2420, AdderIns_s5_bc_0_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_1_a1_U1 ( .a ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, new_AGEMA_signal_2315, AdderIns_g4[16]}), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, new_AGEMA_signal_2423, AdderIns_s5_bc_1_a1_t}), .c ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, new_AGEMA_signal_2483, AdderIns_g5[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, new_AGEMA_signal_2291, AdderIns_g4[8]}), .b ({new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1982, AdderIns_p4[9]}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, new_AGEMA_signal_2423, AdderIns_s5_bc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_2_a1_U1 ( .a ({new_AGEMA_signal_2320, new_AGEMA_signal_2319, new_AGEMA_signal_2318, AdderIns_g4[17]}), .b ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, AdderIns_s5_bc_2_a1_t}), .c ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, new_AGEMA_signal_2486, AdderIns_g5[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_2296, new_AGEMA_signal_2295, new_AGEMA_signal_2294, AdderIns_g4[9]}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, AdderIns_p4[10]}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, AdderIns_s5_bc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_3_a1_U1 ( .a ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, new_AGEMA_signal_2321, AdderIns_g4[18]}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, new_AGEMA_signal_2429, AdderIns_s5_bc_3_a1_t}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, new_AGEMA_signal_2489, AdderIns_g5[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, new_AGEMA_signal_2297, AdderIns_g4[10]}), .b ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, new_AGEMA_signal_1988, AdderIns_p4[11]}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, new_AGEMA_signal_2429, AdderIns_s5_bc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_4_a1_U1 ( .a ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, new_AGEMA_signal_2324, AdderIns_g4[19]}), .b ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, new_AGEMA_signal_2432, AdderIns_s5_bc_4_a1_t}), .c ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, new_AGEMA_signal_2492, AdderIns_g5[19]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, new_AGEMA_signal_2300, AdderIns_g4[11]}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1991, AdderIns_p4[12]}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, new_AGEMA_signal_2432, AdderIns_s5_bc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_5_a1_U1 ( .a ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, AdderIns_g4[20]}), .b ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, new_AGEMA_signal_2435, AdderIns_s5_bc_5_a1_t}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, new_AGEMA_signal_2495, AdderIns_g5[20]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, new_AGEMA_signal_2303, AdderIns_g4[12]}), .b ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, AdderIns_p4[13]}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, new_AGEMA_signal_2435, AdderIns_s5_bc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_6_a1_U1 ( .a ({new_AGEMA_signal_2332, new_AGEMA_signal_2331, new_AGEMA_signal_2330, AdderIns_g4[21]}), .b ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, new_AGEMA_signal_2438, AdderIns_s5_bc_6_a1_t}), .c ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, new_AGEMA_signal_2498, AdderIns_g5[21]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_2308, new_AGEMA_signal_2307, new_AGEMA_signal_2306, AdderIns_g4[13]}), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, new_AGEMA_signal_1997, AdderIns_p4[14]}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, new_AGEMA_signal_2438, AdderIns_s5_bc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_7_a1_U1 ( .a ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, new_AGEMA_signal_2333, AdderIns_g4[22]}), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, new_AGEMA_signal_2441, AdderIns_s5_bc_7_a1_t}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, new_AGEMA_signal_2501, AdderIns_g5[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, new_AGEMA_signal_2309, AdderIns_g4[14]}), .b ({new_AGEMA_signal_2002, new_AGEMA_signal_2001, new_AGEMA_signal_2000, AdderIns_p4[15]}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, new_AGEMA_signal_2441, AdderIns_s5_bc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_8_a1_U1 ( .a ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, new_AGEMA_signal_2336, AdderIns_g4[23]}), .b ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, new_AGEMA_signal_2444, AdderIns_s5_bc_8_a1_t}), .c ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, new_AGEMA_signal_2504, AdderIns_g5[23]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, new_AGEMA_signal_2312, AdderIns_g4[15]}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, AdderIns_p4[16]}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, new_AGEMA_signal_2444, AdderIns_s5_bc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_9_a1_U1 ( .a ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, new_AGEMA_signal_2339, AdderIns_g4[24]}), .b ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, new_AGEMA_signal_2447, AdderIns_s5_bc_9_a1_t}), .c ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, new_AGEMA_signal_2507, AdderIns_g5[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, new_AGEMA_signal_2315, AdderIns_g4[16]}), .b ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, AdderIns_p4[17]}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, new_AGEMA_signal_2447, AdderIns_s5_bc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_10_a1_U1 ( .a ({new_AGEMA_signal_2344, new_AGEMA_signal_2343, new_AGEMA_signal_2342, AdderIns_g4[25]}), .b ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, new_AGEMA_signal_2450, AdderIns_s5_bc_10_a1_t}), .c ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, new_AGEMA_signal_2510, AdderIns_g5[25]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_2320, new_AGEMA_signal_2319, new_AGEMA_signal_2318, AdderIns_g4[17]}), .b ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, new_AGEMA_signal_2009, AdderIns_p4[18]}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, new_AGEMA_signal_2450, AdderIns_s5_bc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_11_a1_U1 ( .a ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, new_AGEMA_signal_2345, AdderIns_g4[26]}), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, new_AGEMA_signal_2453, AdderIns_s5_bc_11_a1_t}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, new_AGEMA_signal_2513, AdderIns_g5[26]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, new_AGEMA_signal_2321, AdderIns_g4[18]}), .b ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, AdderIns_p4[19]}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, new_AGEMA_signal_2453, AdderIns_s5_bc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_12_a1_U1 ( .a ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, new_AGEMA_signal_2348, AdderIns_g4[27]}), .b ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, new_AGEMA_signal_2456, AdderIns_s5_bc_12_a1_t}), .c ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, new_AGEMA_signal_2516, AdderIns_g5[27]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, new_AGEMA_signal_2324, AdderIns_g4[19]}), .b ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2015, AdderIns_p4[20]}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, new_AGEMA_signal_2456, AdderIns_s5_bc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_13_a1_U1 ( .a ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, new_AGEMA_signal_2351, AdderIns_g4[28]}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, new_AGEMA_signal_2459, AdderIns_s5_bc_13_a1_t}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, new_AGEMA_signal_2519, AdderIns_g5[28]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, AdderIns_g4[20]}), .b ({new_AGEMA_signal_2020, new_AGEMA_signal_2019, new_AGEMA_signal_2018, AdderIns_p4[21]}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, new_AGEMA_signal_2459, AdderIns_s5_bc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_14_a1_U1 ( .a ({new_AGEMA_signal_2356, new_AGEMA_signal_2355, new_AGEMA_signal_2354, AdderIns_g4[29]}), .b ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, new_AGEMA_signal_2462, AdderIns_s5_bc_14_a1_t}), .c ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, new_AGEMA_signal_2522, AdderIns_g5[29]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_2332, new_AGEMA_signal_2331, new_AGEMA_signal_2330, AdderIns_g4[21]}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, AdderIns_p4[22]}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, new_AGEMA_signal_2462, AdderIns_s5_bc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_15_a1_U1 ( .a ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, new_AGEMA_signal_2357, AdderIns_g4[30]}), .b ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, new_AGEMA_signal_2465, AdderIns_s5_bc_15_a1_t}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, new_AGEMA_signal_2525, AdderIns_g5[30]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s5_bc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, new_AGEMA_signal_2333, AdderIns_g4[22]}), .b ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2024, AdderIns_p4[23]}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, new_AGEMA_signal_2465, AdderIns_s5_bc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_1_a1_U1 ( .a ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, new_AGEMA_signal_2483, AdderIns_g5[16]}), .b ({new_AGEMA_signal_2272, new_AGEMA_signal_2271, new_AGEMA_signal_2270, AdderIns_s6_gc_1_a1_t}), .c ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, new_AGEMA_signal_2594, AdderIns_g6[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_1_a1_a1_U1 ( .a ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, AdderIns_g6[0]}), .b ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, new_AGEMA_signal_2132, AdderIns_p5[1]}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_2272, new_AGEMA_signal_2271, new_AGEMA_signal_2270, AdderIns_s6_gc_1_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_2_a1_U1 ( .a ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, new_AGEMA_signal_2486, AdderIns_g5[17]}), .b ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, new_AGEMA_signal_2273, AdderIns_s6_gc_2_a1_t}), .c ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, new_AGEMA_signal_2597, AdderIns_g6[17]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_2_a1_a1_U1 ( .a ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, new_AGEMA_signal_1859, AdderIns_g6[1]}), .b ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, new_AGEMA_signal_2135, AdderIns_p5[2]}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, new_AGEMA_signal_2273, AdderIns_s6_gc_2_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_3_a1_U1 ( .a ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, new_AGEMA_signal_2489, AdderIns_g5[18]}), .b ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, new_AGEMA_signal_2276, AdderIns_s6_gc_3_a1_t}), .c ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, new_AGEMA_signal_2600, AdderIns_g6[18]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_3_a1_a1_U1 ( .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, AdderIns_g6[2]}), .b ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, new_AGEMA_signal_2138, AdderIns_p5[3]}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, new_AGEMA_signal_2276, AdderIns_s6_gc_3_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_4_a1_U1 ( .a ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, new_AGEMA_signal_2492, AdderIns_g5[19]}), .b ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, new_AGEMA_signal_2369, AdderIns_s6_gc_4_a1_t}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, new_AGEMA_signal_2603, AdderIns_g6[19]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_4_a1_a1_U1 ( .a ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, AdderIns_g6[3]}), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, new_AGEMA_signal_2141, AdderIns_p5[4]}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, new_AGEMA_signal_2369, AdderIns_s6_gc_4_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_5_a1_U1 ( .a ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, new_AGEMA_signal_2495, AdderIns_g5[20]}), .b ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, new_AGEMA_signal_2372, AdderIns_s6_gc_5_a1_t}), .c ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, new_AGEMA_signal_2606, AdderIns_g6[20]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_5_a1_a1_U1 ( .a ({new_AGEMA_signal_2188, new_AGEMA_signal_2187, new_AGEMA_signal_2186, AdderIns_g6[4]}), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, AdderIns_p5[5]}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, new_AGEMA_signal_2372, AdderIns_s6_gc_5_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_6_a1_U1 ( .a ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, new_AGEMA_signal_2498, AdderIns_g5[21]}), .b ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, new_AGEMA_signal_2375, AdderIns_s6_gc_6_a1_t}), .c ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, new_AGEMA_signal_2609, AdderIns_g6[21]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_6_a1_a1_U1 ( .a ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, AdderIns_g6[5]}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, new_AGEMA_signal_2147, AdderIns_p5[6]}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, new_AGEMA_signal_2375, AdderIns_s6_gc_6_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_7_a1_U1 ( .a ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, new_AGEMA_signal_2501, AdderIns_g5[22]}), .b ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, new_AGEMA_signal_2468, AdderIns_s6_gc_7_a1_t}), .c ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, new_AGEMA_signal_2612, AdderIns_g6[22]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_7_a1_a1_U1 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, new_AGEMA_signal_2285, AdderIns_g6[6]}), .b ({new_AGEMA_signal_2152, new_AGEMA_signal_2151, new_AGEMA_signal_2150, AdderIns_p5[7]}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, new_AGEMA_signal_2468, AdderIns_s6_gc_7_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_8_a1_U1 ( .a ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, new_AGEMA_signal_2504, AdderIns_g5[23]}), .b ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, new_AGEMA_signal_2528, AdderIns_s6_gc_8_a1_t}), .c ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, new_AGEMA_signal_2615, AdderIns_g6[23]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_8_a1_a1_U1 ( .a ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, new_AGEMA_signal_2396, AdderIns_g6[7]}), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, AdderIns_p5[8]}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, new_AGEMA_signal_2528, AdderIns_s6_gc_8_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_9_a1_U1 ( .a ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, new_AGEMA_signal_2507, AdderIns_g5[24]}), .b ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, new_AGEMA_signal_2531, AdderIns_s6_gc_9_a1_t}), .c ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, new_AGEMA_signal_2618, AdderIns_g6[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_9_a1_a1_U1 ( .a ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, AdderIns_g6[8]}), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, new_AGEMA_signal_2156, AdderIns_p5[9]}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, new_AGEMA_signal_2531, AdderIns_s6_gc_9_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_10_a1_U1 ( .a ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, new_AGEMA_signal_2510, AdderIns_g5[25]}), .b ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, new_AGEMA_signal_2534, AdderIns_s6_gc_10_a1_t}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, new_AGEMA_signal_2621, AdderIns_g6[25]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_10_a1_a1_U1 ( .a ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, new_AGEMA_signal_2402, AdderIns_g6[9]}), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, new_AGEMA_signal_2159, AdderIns_p5[10]}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, new_AGEMA_signal_2534, AdderIns_s6_gc_10_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_11_a1_U1 ( .a ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, new_AGEMA_signal_2513, AdderIns_g5[26]}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, new_AGEMA_signal_2537, AdderIns_s6_gc_11_a1_t}), .c ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, new_AGEMA_signal_2624, AdderIns_g6[26]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_11_a1_a1_U1 ( .a ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, new_AGEMA_signal_2405, AdderIns_g6[10]}), .b ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, AdderIns_p5[11]}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, new_AGEMA_signal_2537, AdderIns_s6_gc_11_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_12_a1_U1 ( .a ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, new_AGEMA_signal_2516, AdderIns_g5[27]}), .b ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, new_AGEMA_signal_2540, AdderIns_s6_gc_12_a1_t}), .c ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, new_AGEMA_signal_2627, AdderIns_g6[27]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_12_a1_a1_U1 ( .a ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, new_AGEMA_signal_2408, AdderIns_g6[11]}), .b ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, new_AGEMA_signal_2165, AdderIns_p5[12]}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, new_AGEMA_signal_2540, AdderIns_s6_gc_12_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_13_a1_U1 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, new_AGEMA_signal_2519, AdderIns_g5[28]}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, new_AGEMA_signal_2543, AdderIns_s6_gc_13_a1_t}), .c ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, new_AGEMA_signal_2630, AdderIns_g6[28]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_13_a1_a1_U1 ( .a ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, new_AGEMA_signal_2411, AdderIns_g6[12]}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, new_AGEMA_signal_2168, AdderIns_p5[13]}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, new_AGEMA_signal_2543, AdderIns_s6_gc_13_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_14_a1_U1 ( .a ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, new_AGEMA_signal_2522, AdderIns_g5[29]}), .b ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, new_AGEMA_signal_2546, AdderIns_s6_gc_14_a1_t}), .c ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, new_AGEMA_signal_2633, AdderIns_g6[29]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_14_a1_a1_U1 ( .a ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, new_AGEMA_signal_2414, AdderIns_g6[13]}), .b ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, new_AGEMA_signal_2171, AdderIns_p5[14]}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, new_AGEMA_signal_2546, AdderIns_s6_gc_14_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_15_a1_U1 ( .a ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, new_AGEMA_signal_2525, AdderIns_g5[30]}), .b ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, new_AGEMA_signal_2636, AdderIns_s6_gc_15_a1_t}), .c ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, new_AGEMA_signal_2672, AdderIns_g6[30]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s6_gc_15_a1_a1_U1 ( .a ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, new_AGEMA_signal_2477, AdderIns_g6[14]}), .b ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, AdderIns_p5[15]}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, new_AGEMA_signal_2636, AdderIns_s6_gc_15_a1_t}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U24 ( .a ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, new_AGEMA_signal_2672, AdderIns_g6[30]}), .b ({new_AGEMA_signal_1492, new_AGEMA_signal_1491, new_AGEMA_signal_1490, AdderIns_p6[31]}), .c ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2771, sum[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U23 ( .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, new_AGEMA_signal_2633, AdderIns_g6[29]}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, new_AGEMA_signal_1481, AdderIns_p6[30]}), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, sum[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U21 ( .a ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, new_AGEMA_signal_2630, AdderIns_g6[28]}), .b ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, new_AGEMA_signal_1472, AdderIns_p6[29]}), .c ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, new_AGEMA_signal_2678, sum[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U20 ( .a ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, new_AGEMA_signal_2627, AdderIns_g6[27]}), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, new_AGEMA_signal_1463, AdderIns_p6[28]}), .c ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, new_AGEMA_signal_2681, sum[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U19 ( .a ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, new_AGEMA_signal_2624, AdderIns_g6[26]}), .b ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, AdderIns_p6[27]}), .c ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, sum[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U18 ( .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, new_AGEMA_signal_2621, AdderIns_g6[25]}), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, new_AGEMA_signal_1445, AdderIns_p6[26]}), .c ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2687, sum[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U17 ( .a ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, new_AGEMA_signal_2618, AdderIns_g6[24]}), .b ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, new_AGEMA_signal_1436, AdderIns_p6[25]}), .c ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, sum[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U16 ( .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, new_AGEMA_signal_2615, AdderIns_g6[23]}), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, AdderIns_p6[24]}), .c ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, sum[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U15 ( .a ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, new_AGEMA_signal_2612, AdderIns_g6[22]}), .b ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, AdderIns_p6[23]}), .c ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, new_AGEMA_signal_2696, sum[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U14 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, new_AGEMA_signal_2609, AdderIns_g6[21]}), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, new_AGEMA_signal_1409, AdderIns_p6[22]}), .c ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, sum[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U13 ( .a ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, new_AGEMA_signal_2606, AdderIns_g6[20]}), .b ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, new_AGEMA_signal_1400, AdderIns_p6[21]}), .c ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, sum[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U12 ( .a ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, new_AGEMA_signal_2603, AdderIns_g6[19]}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, AdderIns_p6[20]}), .c ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, new_AGEMA_signal_2705, sum[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U10 ( .a ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, new_AGEMA_signal_2600, AdderIns_g6[18]}), .b ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, new_AGEMA_signal_1382, AdderIns_p6[19]}), .c ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, sum[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U9 ( .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, new_AGEMA_signal_2597, AdderIns_g6[17]}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, new_AGEMA_signal_1373, AdderIns_p6[18]}), .c ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, sum[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U8 ( .a ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, new_AGEMA_signal_2594, AdderIns_g6[16]}), .b ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, new_AGEMA_signal_1364, AdderIns_p6[17]}), .c ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, sum[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AdderIns_s7_U7 ( .a ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, new_AGEMA_signal_2480, AdderIns_g6[15]}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, new_AGEMA_signal_1355, AdderIns_p6[16]}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, sum[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_0_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, sum[24]}), .a ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, sum[17]}), .c ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, new_AGEMA_signal_2774, sum_rotated01[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_1_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, sum[25]}), .a ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, sum[18]}), .c ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, new_AGEMA_signal_2777, sum_rotated01[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_2_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2687, sum[26]}), .a ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, sum[19]}), .c ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, new_AGEMA_signal_2780, sum_rotated01[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_3_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, sum[27]}), .a ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, new_AGEMA_signal_2705, sum[20]}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, new_AGEMA_signal_2783, sum_rotated01[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_4_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, new_AGEMA_signal_2681, sum[28]}), .a ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, sum[21]}), .c ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, new_AGEMA_signal_2786, sum_rotated01[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_5_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, new_AGEMA_signal_2678, sum[29]}), .a ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, sum[22]}), .c ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, new_AGEMA_signal_2789, sum_rotated01[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_6_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, sum[30]}), .a ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, new_AGEMA_signal_2696, sum[23]}), .c ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, new_AGEMA_signal_2792, sum_rotated01[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_7_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2771, sum[31]}), .a ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, sum[24]}), .c ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, new_AGEMA_signal_2933, sum_rotated01[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_8_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, new_AGEMA_signal_1211, sum[0]}), .a ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, sum[25]}), .c ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, new_AGEMA_signal_2795, sum_rotated01[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_9_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, new_AGEMA_signal_2027, sum[1]}), .a ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2687, sum[26]}), .c ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, new_AGEMA_signal_2798, sum_rotated01[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_10_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, sum[2]}), .a ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, sum[27]}), .c ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, new_AGEMA_signal_2801, sum_rotated01[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_11_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, sum[3]}), .a ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, new_AGEMA_signal_2681, sum[28]}), .c ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, new_AGEMA_signal_2804, sum_rotated01[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_12_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, new_AGEMA_signal_2384, sum[4]}), .a ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, new_AGEMA_signal_2678, sum[29]}), .c ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, new_AGEMA_signal_2807, sum_rotated01[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_13_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, sum[5]}), .a ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, sum[30]}), .c ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810, sum_rotated01[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_14_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, new_AGEMA_signal_2378, sum[6]}), .a ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2771, sum[31]}), .c ({new_AGEMA_signal_2938, new_AGEMA_signal_2937, new_AGEMA_signal_2936, sum_rotated01[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_24_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, sum[16]}), .a ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, new_AGEMA_signal_2549, sum[9]}), .c ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, sum_rotated01[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_25_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, sum[17]}), .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, sum[10]}), .c ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, new_AGEMA_signal_2813, sum_rotated01[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_26_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, sum[18]}), .a ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, new_AGEMA_signal_2564, sum[11]}), .c ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, new_AGEMA_signal_2816, sum_rotated01[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_27_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, sum[19]}), .a ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, new_AGEMA_signal_2561, sum[12]}), .c ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, new_AGEMA_signal_2819, sum_rotated01[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_28_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, new_AGEMA_signal_2705, sum[20]}), .a ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, sum[13]}), .c ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, new_AGEMA_signal_2822, sum_rotated01[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_29_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, sum[21]}), .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, new_AGEMA_signal_2555, sum[14]}), .c ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, new_AGEMA_signal_2825, sum_rotated01[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_30_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, sum[22]}), .a ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, new_AGEMA_signal_2642, sum[15]}), .c ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, new_AGEMA_signal_2828, sum_rotated01[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M4_mux_inst_31_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, new_AGEMA_signal_2696, sum[23]}), .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, sum[16]}), .c ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, new_AGEMA_signal_2831, sum_rotated01[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_0_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2771, sum[31]}), .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, sum[16]}), .c ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, new_AGEMA_signal_2939, sum_rotated23[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_1_U1 ( .s (round[0]), .b ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, new_AGEMA_signal_1211, sum[0]}), .a ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, sum[17]}), .c ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, new_AGEMA_signal_2834, sum_rotated23[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_2_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, new_AGEMA_signal_2027, sum[1]}), .a ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, sum[18]}), .c ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, new_AGEMA_signal_2837, sum_rotated23[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_3_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, sum[2]}), .a ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, sum[19]}), .c ({new_AGEMA_signal_2842, new_AGEMA_signal_2841, new_AGEMA_signal_2840, sum_rotated23[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_4_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, sum[3]}), .a ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, new_AGEMA_signal_2705, sum[20]}), .c ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, new_AGEMA_signal_2843, sum_rotated23[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_5_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, new_AGEMA_signal_2384, sum[4]}), .a ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, sum[21]}), .c ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, sum_rotated23[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_6_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, sum[5]}), .a ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, sum[22]}), .c ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, new_AGEMA_signal_2849, sum_rotated23[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_7_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, new_AGEMA_signal_2378, sum[6]}), .a ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, new_AGEMA_signal_2696, sum[23]}), .c ({new_AGEMA_signal_2854, new_AGEMA_signal_2853, new_AGEMA_signal_2852, sum_rotated23[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_8_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, sum[7]}), .a ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, sum[24]}), .c ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, new_AGEMA_signal_2855, sum_rotated23[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_9_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, new_AGEMA_signal_2552, sum[8]}), .a ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, sum[25]}), .c ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, new_AGEMA_signal_2858, sum_rotated23[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_10_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, new_AGEMA_signal_2549, sum[9]}), .a ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2687, sum[26]}), .c ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, new_AGEMA_signal_2861, sum_rotated23[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_11_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, sum[10]}), .a ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, sum[27]}), .c ({new_AGEMA_signal_2866, new_AGEMA_signal_2865, new_AGEMA_signal_2864, sum_rotated23[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_12_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, new_AGEMA_signal_2564, sum[11]}), .a ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, new_AGEMA_signal_2681, sum[28]}), .c ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, new_AGEMA_signal_2867, sum_rotated23[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_13_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, new_AGEMA_signal_2561, sum[12]}), .a ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, new_AGEMA_signal_2678, sum[29]}), .c ({new_AGEMA_signal_2872, new_AGEMA_signal_2871, new_AGEMA_signal_2870, sum_rotated23[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_14_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, sum[13]}), .a ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, sum[30]}), .c ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, new_AGEMA_signal_2873, sum_rotated23[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_15_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, new_AGEMA_signal_2555, sum[14]}), .a ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2771, sum[31]}), .c ({new_AGEMA_signal_2944, new_AGEMA_signal_2943, new_AGEMA_signal_2942, sum_rotated23[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_17_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, sum[16]}), .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, new_AGEMA_signal_2027, sum[1]}), .c ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, sum_rotated23[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_18_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, sum[17]}), .a ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, sum[2]}), .c ({new_AGEMA_signal_2878, new_AGEMA_signal_2877, new_AGEMA_signal_2876, sum_rotated23[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_19_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, sum[18]}), .a ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, sum[3]}), .c ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, new_AGEMA_signal_2879, sum_rotated23[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_20_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, sum[19]}), .a ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, new_AGEMA_signal_2384, sum[4]}), .c ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, new_AGEMA_signal_2882, sum_rotated23[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_21_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, new_AGEMA_signal_2705, sum[20]}), .a ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, sum[5]}), .c ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, new_AGEMA_signal_2885, sum_rotated23[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_22_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, sum[21]}), .a ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, new_AGEMA_signal_2378, sum[6]}), .c ({new_AGEMA_signal_2890, new_AGEMA_signal_2889, new_AGEMA_signal_2888, sum_rotated23[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_23_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, sum[22]}), .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, sum[7]}), .c ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, new_AGEMA_signal_2891, sum_rotated23[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_24_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, new_AGEMA_signal_2696, sum[23]}), .a ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, new_AGEMA_signal_2552, sum[8]}), .c ({new_AGEMA_signal_2896, new_AGEMA_signal_2895, new_AGEMA_signal_2894, sum_rotated23[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_25_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, sum[24]}), .a ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, new_AGEMA_signal_2549, sum[9]}), .c ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, new_AGEMA_signal_2897, sum_rotated23[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_26_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, sum[25]}), .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, sum[10]}), .c ({new_AGEMA_signal_2902, new_AGEMA_signal_2901, new_AGEMA_signal_2900, sum_rotated23[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_27_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2687, sum[26]}), .a ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, new_AGEMA_signal_2564, sum[11]}), .c ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, new_AGEMA_signal_2903, sum_rotated23[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_28_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, sum[27]}), .a ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, new_AGEMA_signal_2561, sum[12]}), .c ({new_AGEMA_signal_2908, new_AGEMA_signal_2907, new_AGEMA_signal_2906, sum_rotated23[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_29_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, new_AGEMA_signal_2681, sum[28]}), .a ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, sum[13]}), .c ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, new_AGEMA_signal_2909, sum_rotated23[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_30_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, new_AGEMA_signal_2678, sum[29]}), .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, new_AGEMA_signal_2555, sum[14]}), .c ({new_AGEMA_signal_2914, new_AGEMA_signal_2913, new_AGEMA_signal_2912, sum_rotated23[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M5_mux_inst_31_U1 ( .s (round[0]), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, sum[30]}), .a ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, new_AGEMA_signal_2642, sum[15]}), .c ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, new_AGEMA_signal_2915, sum_rotated23[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_0_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, new_AGEMA_signal_2774, sum_rotated01[0]}), .a ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, new_AGEMA_signal_2939, sum_rotated23[0]}), .c ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, new_AGEMA_signal_3101, sum_rotated[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_1_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, new_AGEMA_signal_2777, sum_rotated01[1]}), .a ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, new_AGEMA_signal_2834, sum_rotated23[1]}), .c ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, new_AGEMA_signal_2945, sum_rotated[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_2_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, new_AGEMA_signal_2780, sum_rotated01[2]}), .a ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, new_AGEMA_signal_2837, sum_rotated23[2]}), .c ({new_AGEMA_signal_2950, new_AGEMA_signal_2949, new_AGEMA_signal_2948, sum_rotated[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_3_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, new_AGEMA_signal_2783, sum_rotated01[3]}), .a ({new_AGEMA_signal_2842, new_AGEMA_signal_2841, new_AGEMA_signal_2840, sum_rotated23[3]}), .c ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, new_AGEMA_signal_2951, sum_rotated[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_4_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, new_AGEMA_signal_2786, sum_rotated01[4]}), .a ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, new_AGEMA_signal_2843, sum_rotated23[4]}), .c ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, new_AGEMA_signal_2954, sum_rotated[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_5_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, new_AGEMA_signal_2789, sum_rotated01[5]}), .a ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, sum_rotated23[5]}), .c ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, new_AGEMA_signal_2957, sum_rotated[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_6_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, new_AGEMA_signal_2792, sum_rotated01[6]}), .a ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, new_AGEMA_signal_2849, sum_rotated23[6]}), .c ({new_AGEMA_signal_2962, new_AGEMA_signal_2961, new_AGEMA_signal_2960, sum_rotated[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_7_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, new_AGEMA_signal_2933, sum_rotated01[7]}), .a ({new_AGEMA_signal_2854, new_AGEMA_signal_2853, new_AGEMA_signal_2852, sum_rotated23[7]}), .c ({new_AGEMA_signal_3106, new_AGEMA_signal_3105, new_AGEMA_signal_3104, sum_rotated[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_8_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, new_AGEMA_signal_2795, sum_rotated01[8]}), .a ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, new_AGEMA_signal_2855, sum_rotated23[8]}), .c ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, new_AGEMA_signal_2963, sum_rotated[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_9_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, new_AGEMA_signal_2798, sum_rotated01[9]}), .a ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, new_AGEMA_signal_2858, sum_rotated23[9]}), .c ({new_AGEMA_signal_2968, new_AGEMA_signal_2967, new_AGEMA_signal_2966, sum_rotated[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_10_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, new_AGEMA_signal_2801, sum_rotated01[10]}), .a ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, new_AGEMA_signal_2861, sum_rotated23[10]}), .c ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, new_AGEMA_signal_2969, sum_rotated[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_11_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, new_AGEMA_signal_2804, sum_rotated01[11]}), .a ({new_AGEMA_signal_2866, new_AGEMA_signal_2865, new_AGEMA_signal_2864, sum_rotated23[11]}), .c ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, new_AGEMA_signal_2972, sum_rotated[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_12_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, new_AGEMA_signal_2807, sum_rotated01[12]}), .a ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, new_AGEMA_signal_2867, sum_rotated23[12]}), .c ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, new_AGEMA_signal_2975, sum_rotated[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_13_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810, sum_rotated01[13]}), .a ({new_AGEMA_signal_2872, new_AGEMA_signal_2871, new_AGEMA_signal_2870, sum_rotated23[13]}), .c ({new_AGEMA_signal_2980, new_AGEMA_signal_2979, new_AGEMA_signal_2978, sum_rotated[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_14_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2938, new_AGEMA_signal_2937, new_AGEMA_signal_2936, sum_rotated01[14]}), .a ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, new_AGEMA_signal_2873, sum_rotated23[14]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3107, sum_rotated[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_15_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, new_AGEMA_signal_2570, sum_rotated01[15]}), .a ({new_AGEMA_signal_2944, new_AGEMA_signal_2943, new_AGEMA_signal_2942, sum_rotated23[15]}), .c ({new_AGEMA_signal_3112, new_AGEMA_signal_3111, new_AGEMA_signal_3110, sum_rotated[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_17_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, new_AGEMA_signal_2648, sum_rotated01[17]}), .a ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, sum_rotated23[17]}), .c ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, new_AGEMA_signal_2921, sum_rotated[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_18_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, new_AGEMA_signal_2651, sum_rotated01[18]}), .a ({new_AGEMA_signal_2878, new_AGEMA_signal_2877, new_AGEMA_signal_2876, sum_rotated23[18]}), .c ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, new_AGEMA_signal_2981, sum_rotated[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_19_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, new_AGEMA_signal_2654, sum_rotated01[19]}), .a ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, new_AGEMA_signal_2879, sum_rotated23[19]}), .c ({new_AGEMA_signal_2986, new_AGEMA_signal_2985, new_AGEMA_signal_2984, sum_rotated[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_20_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, new_AGEMA_signal_2657, sum_rotated01[20]}), .a ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, new_AGEMA_signal_2882, sum_rotated23[20]}), .c ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, new_AGEMA_signal_2987, sum_rotated[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_21_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, new_AGEMA_signal_2660, sum_rotated01[21]}), .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, new_AGEMA_signal_2885, sum_rotated23[21]}), .c ({new_AGEMA_signal_2992, new_AGEMA_signal_2991, new_AGEMA_signal_2990, sum_rotated[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_22_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, new_AGEMA_signal_2663, sum_rotated01[22]}), .a ({new_AGEMA_signal_2890, new_AGEMA_signal_2889, new_AGEMA_signal_2888, sum_rotated23[22]}), .c ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, new_AGEMA_signal_2993, sum_rotated[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_23_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, new_AGEMA_signal_2717, sum_rotated01[23]}), .a ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, new_AGEMA_signal_2891, sum_rotated23[23]}), .c ({new_AGEMA_signal_2998, new_AGEMA_signal_2997, new_AGEMA_signal_2996, sum_rotated[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_24_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, sum_rotated01[24]}), .a ({new_AGEMA_signal_2896, new_AGEMA_signal_2895, new_AGEMA_signal_2894, sum_rotated23[24]}), .c ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, new_AGEMA_signal_2999, sum_rotated[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_25_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, new_AGEMA_signal_2813, sum_rotated01[25]}), .a ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, new_AGEMA_signal_2897, sum_rotated23[25]}), .c ({new_AGEMA_signal_3004, new_AGEMA_signal_3003, new_AGEMA_signal_3002, sum_rotated[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_26_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, new_AGEMA_signal_2816, sum_rotated01[26]}), .a ({new_AGEMA_signal_2902, new_AGEMA_signal_2901, new_AGEMA_signal_2900, sum_rotated23[26]}), .c ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, new_AGEMA_signal_3005, sum_rotated[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_27_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, new_AGEMA_signal_2819, sum_rotated01[27]}), .a ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, new_AGEMA_signal_2903, sum_rotated23[27]}), .c ({new_AGEMA_signal_3010, new_AGEMA_signal_3009, new_AGEMA_signal_3008, sum_rotated[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_28_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, new_AGEMA_signal_2822, sum_rotated01[28]}), .a ({new_AGEMA_signal_2908, new_AGEMA_signal_2907, new_AGEMA_signal_2906, sum_rotated23[28]}), .c ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, new_AGEMA_signal_3011, sum_rotated[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_29_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, new_AGEMA_signal_2825, sum_rotated01[29]}), .a ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, new_AGEMA_signal_2909, sum_rotated23[29]}), .c ({new_AGEMA_signal_3016, new_AGEMA_signal_3015, new_AGEMA_signal_3014, sum_rotated[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_30_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, new_AGEMA_signal_2828, sum_rotated01[30]}), .a ({new_AGEMA_signal_2914, new_AGEMA_signal_2913, new_AGEMA_signal_2912, sum_rotated23[30]}), .c ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, new_AGEMA_signal_3017, sum_rotated[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) M6_mux_inst_31_U1 ( .s (round[1]), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, new_AGEMA_signal_2831, sum_rotated01[31]}), .a ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, new_AGEMA_signal_2915, sum_rotated23[31]}), .c ({new_AGEMA_signal_3022, new_AGEMA_signal_3021, new_AGEMA_signal_3020, sum_rotated[31]}) ) ;

endmodule
