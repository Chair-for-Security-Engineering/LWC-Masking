/* modified netlist. Source: module RoundFunction in file ./test/RoundFunction.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module RoundFunction_HPC2_ClockGating_d1 (ROUND_KEY_s0, /*ROUND_KEY,*/ ROUND_IN_s0, CONST_IN, clk, ROUND_KEY_s1, ROUND_IN_s1, Fresh, /*rst,*/ ROUND_OUT_s0, ROUND_OUT_s1/*, Synch*/);
    input [383:0] ROUND_KEY_s0 ;
    //input [319:0] ROUND_KEY ;
    input [127:0] ROUND_IN_s0 ;
    input [5:0] CONST_IN ;
    input clk ;
    input [383:0] ROUND_KEY_s1 ;
    input [127:0] ROUND_IN_s1 ;
    //input rst ;
    input [127:0] Fresh ;
    output [127:0] ROUND_OUT_s0 ;
    output [127:0] ROUND_OUT_s1 ;
    //output Synch ;
    wire SUBSTITUTION_89 ;
    wire SUBSTITUTION_88 ;
    wire SUBSTITUTION_57 ;
    wire n405 ;
    wire n406 ;
    wire n407 ;
    wire n408 ;
    wire n409 ;
    wire n410 ;
    wire n411 ;
    wire n412 ;
    wire n413 ;
    wire n414 ;
    wire n415 ;
    wire n416 ;
    wire n417 ;
    wire n418 ;
    wire n419 ;
    wire n420 ;
    wire n421 ;
    wire n422 ;
    wire n423 ;
    wire n424 ;
    wire n425 ;
    wire n426 ;
    wire n427 ;
    wire n428 ;
    wire n429 ;
    wire n430 ;
    wire n431 ;
    wire n432 ;
    wire n433 ;
    wire n434 ;
    wire n435 ;
    wire n436 ;
    wire n437 ;
    wire n438 ;
    wire n439 ;
    wire n440 ;
    wire n441 ;
    wire n442 ;
    wire n443 ;
    wire n444 ;
    wire n445 ;
    wire n446 ;
    wire n447 ;
    wire n448 ;
    wire n449 ;
    wire n450 ;
    wire n451 ;
    wire n452 ;
    wire n453 ;
    wire n454 ;
    wire n455 ;
    wire n456 ;
    wire n457 ;
    wire n458 ;
    wire n459 ;
    wire n460 ;
    wire n461 ;
    wire n462 ;
    wire n463 ;
    wire n464 ;
    wire n465 ;
    wire n466 ;
    wire n467 ;
    wire n468 ;
    wire n469 ;
    wire n470 ;
    wire n471 ;
    wire n472 ;
    wire n473 ;
    wire n474 ;
    wire n475 ;
    wire n476 ;
    wire n477 ;
    wire n478 ;
    wire n479 ;
    wire n480 ;
    wire n481 ;
    wire n482 ;
    wire n483 ;
    wire n484 ;
    wire n485 ;
    wire n486 ;
    wire n487 ;
    wire n488 ;
    wire n489 ;
    wire n490 ;
    wire n491 ;
    wire n492 ;
    wire n493 ;
    wire n494 ;
    wire n495 ;
    wire n496 ;
    wire n497 ;
    wire n498 ;
    wire n499 ;
    wire n500 ;
    wire n501 ;
    wire n502 ;
    wire n503 ;
    wire n504 ;
    wire n505 ;
    wire n506 ;
    wire n507 ;
    wire n508 ;
    wire n509 ;
    wire n510 ;
    wire n511 ;
    wire n512 ;
    wire n513 ;
    wire n514 ;
    wire n515 ;
    wire n516 ;
    wire n517 ;
    wire n518 ;
    wire n519 ;
    wire n520 ;
    wire n521 ;
    wire n522 ;
    wire n523 ;
    wire n524 ;
    wire n525 ;
    wire n526 ;
    wire n527 ;
    wire n528 ;
    wire n529 ;
    wire n530 ;
    wire n531 ;
    wire n532 ;
    wire n533 ;
    wire n534 ;
    wire n535 ;
    wire n536 ;
    wire n537 ;
    wire n538 ;
    wire [123:120] SUBSTITUTION ;
    wire [127:64] CONST_ADDITION ;
    wire [95:0] SHIFTROWS ;
    wire [3:0] S_0_R2 ;
    wire [3:0] S_0_R1 ;
    wire [3:0] S_1_R2 ;
    wire [3:0] S_1_R1 ;
    wire [3:0] S_2_R2 ;
    wire [3:0] S_2_R1 ;
    wire [3:0] S_3_R2 ;
    wire [3:0] S_3_R1 ;
    wire [3:0] S_4_R2 ;
    wire [3:0] S_4_R1 ;
    wire [3:0] S_5_R2 ;
    wire [3:0] S_5_R1 ;
    wire [3:0] S_6_R2 ;
    wire [3:0] S_6_R1 ;
    wire [3:0] S_7_R2 ;
    wire [3:0] S_7_R1 ;
    wire [3:0] S_8_R2 ;
    wire [3:0] S_8_R1 ;
    wire [3:0] S_9_R2 ;
    wire [3:0] S_9_R1 ;
    wire [3:0] S_10_R2 ;
    wire [3:0] S_10_R1 ;
    wire [3:0] S_11_R2 ;
    wire [3:0] S_11_R1 ;
    wire [3:0] S_12_R2 ;
    wire [3:0] S_12_R1 ;
    wire [3:0] S_13_R2 ;
    wire [3:0] S_13_R1 ;
    wire [3:0] S_14_R2 ;
    wire [3:0] S_14_R1 ;
    wire [3:0] S_15_R2 ;
    wire [3:0] S_15_R1 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1938 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) U400 ( .a ({ROUND_KEY_s1[227], ROUND_KEY_s0[227]}), .b ({ROUND_KEY_s1[99], ROUND_KEY_s0[99]}), .c ({new_AGEMA_signal_1084, n406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U403 ( .a ({ROUND_KEY_s1[226], ROUND_KEY_s0[226]}), .b ({ROUND_KEY_s1[98], ROUND_KEY_s0[98]}), .c ({new_AGEMA_signal_1087, n408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U406 ( .a ({ROUND_KEY_s1[225], ROUND_KEY_s0[225]}), .b ({ROUND_KEY_s1[97], ROUND_KEY_s0[97]}), .c ({new_AGEMA_signal_1090, n410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U409 ( .a ({ROUND_KEY_s1[224], ROUND_KEY_s0[224]}), .b ({ROUND_KEY_s1[96], ROUND_KEY_s0[96]}), .c ({new_AGEMA_signal_1093, n412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U412 ( .a ({ROUND_KEY_s1[223], ROUND_KEY_s0[223]}), .b ({ROUND_KEY_s1[95], ROUND_KEY_s0[95]}), .c ({new_AGEMA_signal_1096, n414}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U415 ( .a ({ROUND_KEY_s1[222], ROUND_KEY_s0[222]}), .b ({ROUND_KEY_s1[94], ROUND_KEY_s0[94]}), .c ({new_AGEMA_signal_1099, n416}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U418 ( .a ({ROUND_KEY_s1[221], ROUND_KEY_s0[221]}), .b ({ROUND_KEY_s1[93], ROUND_KEY_s0[93]}), .c ({new_AGEMA_signal_1102, n418}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U421 ( .a ({ROUND_KEY_s1[220], ROUND_KEY_s0[220]}), .b ({ROUND_KEY_s1[92], ROUND_KEY_s0[92]}), .c ({new_AGEMA_signal_1105, n420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U424 ( .a ({ROUND_KEY_s1[219], ROUND_KEY_s0[219]}), .b ({ROUND_KEY_s1[91], ROUND_KEY_s0[91]}), .c ({new_AGEMA_signal_1108, n422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U427 ( .a ({ROUND_KEY_s1[218], ROUND_KEY_s0[218]}), .b ({ROUND_KEY_s1[90], ROUND_KEY_s0[90]}), .c ({new_AGEMA_signal_1111, n424}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U430 ( .a ({ROUND_KEY_s1[217], ROUND_KEY_s0[217]}), .b ({ROUND_KEY_s1[89], ROUND_KEY_s0[89]}), .c ({new_AGEMA_signal_1114, n426}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U434 ( .a ({ROUND_KEY_s1[216], ROUND_KEY_s0[216]}), .b ({ROUND_KEY_s1[88], ROUND_KEY_s0[88]}), .c ({new_AGEMA_signal_1117, n429}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U438 ( .a ({ROUND_KEY_s1[215], ROUND_KEY_s0[215]}), .b ({ROUND_KEY_s1[87], ROUND_KEY_s0[87]}), .c ({new_AGEMA_signal_1120, n432}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U441 ( .a ({ROUND_KEY_s1[214], ROUND_KEY_s0[214]}), .b ({ROUND_KEY_s1[86], ROUND_KEY_s0[86]}), .c ({new_AGEMA_signal_1123, n434}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U444 ( .a ({ROUND_KEY_s1[213], ROUND_KEY_s0[213]}), .b ({ROUND_KEY_s1[85], ROUND_KEY_s0[85]}), .c ({new_AGEMA_signal_1126, n436}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U447 ( .a ({ROUND_KEY_s1[212], ROUND_KEY_s0[212]}), .b ({ROUND_KEY_s1[84], ROUND_KEY_s0[84]}), .c ({new_AGEMA_signal_1129, n438}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U450 ( .a ({ROUND_KEY_s1[211], ROUND_KEY_s0[211]}), .b ({ROUND_KEY_s1[83], ROUND_KEY_s0[83]}), .c ({new_AGEMA_signal_1132, n440}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U453 ( .a ({ROUND_KEY_s1[210], ROUND_KEY_s0[210]}), .b ({ROUND_KEY_s1[82], ROUND_KEY_s0[82]}), .c ({new_AGEMA_signal_1135, n442}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U456 ( .a ({ROUND_KEY_s1[209], ROUND_KEY_s0[209]}), .b ({ROUND_KEY_s1[81], ROUND_KEY_s0[81]}), .c ({new_AGEMA_signal_1138, n444}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U459 ( .a ({ROUND_KEY_s1[208], ROUND_KEY_s0[208]}), .b ({ROUND_KEY_s1[80], ROUND_KEY_s0[80]}), .c ({new_AGEMA_signal_1141, n446}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U462 ( .a ({ROUND_KEY_s1[207], ROUND_KEY_s0[207]}), .b ({ROUND_KEY_s1[79], ROUND_KEY_s0[79]}), .c ({new_AGEMA_signal_1144, n448}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U465 ( .a ({ROUND_KEY_s1[206], ROUND_KEY_s0[206]}), .b ({ROUND_KEY_s1[78], ROUND_KEY_s0[78]}), .c ({new_AGEMA_signal_1147, n450}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U468 ( .a ({ROUND_KEY_s1[205], ROUND_KEY_s0[205]}), .b ({ROUND_KEY_s1[77], ROUND_KEY_s0[77]}), .c ({new_AGEMA_signal_1150, n452}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U471 ( .a ({ROUND_KEY_s1[204], ROUND_KEY_s0[204]}), .b ({ROUND_KEY_s1[76], ROUND_KEY_s0[76]}), .c ({new_AGEMA_signal_1153, n454}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U474 ( .a ({ROUND_KEY_s1[203], ROUND_KEY_s0[203]}), .b ({ROUND_KEY_s1[75], ROUND_KEY_s0[75]}), .c ({new_AGEMA_signal_1156, n456}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U477 ( .a ({ROUND_KEY_s1[202], ROUND_KEY_s0[202]}), .b ({ROUND_KEY_s1[74], ROUND_KEY_s0[74]}), .c ({new_AGEMA_signal_1159, n458}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U480 ( .a ({ROUND_KEY_s1[201], ROUND_KEY_s0[201]}), .b ({ROUND_KEY_s1[73], ROUND_KEY_s0[73]}), .c ({new_AGEMA_signal_1162, n460}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U483 ( .a ({ROUND_KEY_s1[200], ROUND_KEY_s0[200]}), .b ({ROUND_KEY_s1[72], ROUND_KEY_s0[72]}), .c ({new_AGEMA_signal_1165, n462}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U486 ( .a ({ROUND_KEY_s1[199], ROUND_KEY_s0[199]}), .b ({ROUND_KEY_s1[71], ROUND_KEY_s0[71]}), .c ({new_AGEMA_signal_1168, n464}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U489 ( .a ({ROUND_KEY_s1[198], ROUND_KEY_s0[198]}), .b ({ROUND_KEY_s1[70], ROUND_KEY_s0[70]}), .c ({new_AGEMA_signal_1171, n466}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U492 ( .a ({ROUND_KEY_s1[197], ROUND_KEY_s0[197]}), .b ({ROUND_KEY_s1[69], ROUND_KEY_s0[69]}), .c ({new_AGEMA_signal_1174, n468}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U495 ( .a ({ROUND_KEY_s1[196], ROUND_KEY_s0[196]}), .b ({ROUND_KEY_s1[68], ROUND_KEY_s0[68]}), .c ({new_AGEMA_signal_1177, n470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U498 ( .a ({ROUND_KEY_s1[195], ROUND_KEY_s0[195]}), .b ({ROUND_KEY_s1[67], ROUND_KEY_s0[67]}), .c ({new_AGEMA_signal_1180, n472}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U501 ( .a ({ROUND_KEY_s1[194], ROUND_KEY_s0[194]}), .b ({ROUND_KEY_s1[66], ROUND_KEY_s0[66]}), .c ({new_AGEMA_signal_1183, n474}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U504 ( .a ({ROUND_KEY_s1[193], ROUND_KEY_s0[193]}), .b ({ROUND_KEY_s1[65], ROUND_KEY_s0[65]}), .c ({new_AGEMA_signal_1186, n476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U507 ( .a ({ROUND_KEY_s1[192], ROUND_KEY_s0[192]}), .b ({ROUND_KEY_s1[64], ROUND_KEY_s0[64]}), .c ({new_AGEMA_signal_1189, n478}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U510 ( .a ({ROUND_KEY_s1[127], ROUND_KEY_s0[127]}), .b ({ROUND_KEY_s1[255], ROUND_KEY_s0[255]}), .c ({new_AGEMA_signal_1192, n480}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U513 ( .a ({ROUND_KEY_s1[126], ROUND_KEY_s0[126]}), .b ({ROUND_KEY_s1[254], ROUND_KEY_s0[254]}), .c ({new_AGEMA_signal_1195, n482}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U516 ( .a ({ROUND_KEY_s1[125], ROUND_KEY_s0[125]}), .b ({ROUND_KEY_s1[253], ROUND_KEY_s0[253]}), .c ({new_AGEMA_signal_1198, n484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U519 ( .a ({ROUND_KEY_s1[124], ROUND_KEY_s0[124]}), .b ({ROUND_KEY_s1[252], ROUND_KEY_s0[252]}), .c ({new_AGEMA_signal_1201, n486}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U522 ( .a ({ROUND_KEY_s1[123], ROUND_KEY_s0[123]}), .b ({ROUND_KEY_s1[251], ROUND_KEY_s0[251]}), .c ({new_AGEMA_signal_1204, n488}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U526 ( .a ({ROUND_KEY_s1[122], ROUND_KEY_s0[122]}), .b ({ROUND_KEY_s1[250], ROUND_KEY_s0[250]}), .c ({new_AGEMA_signal_1207, n491}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U530 ( .a ({ROUND_KEY_s1[121], ROUND_KEY_s0[121]}), .b ({ROUND_KEY_s1[249], ROUND_KEY_s0[249]}), .c ({new_AGEMA_signal_1210, n494}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U534 ( .a ({ROUND_KEY_s1[120], ROUND_KEY_s0[120]}), .b ({ROUND_KEY_s1[248], ROUND_KEY_s0[248]}), .c ({new_AGEMA_signal_1213, n497}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U538 ( .a ({ROUND_KEY_s1[119], ROUND_KEY_s0[119]}), .b ({ROUND_KEY_s1[247], ROUND_KEY_s0[247]}), .c ({new_AGEMA_signal_1216, n500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U541 ( .a ({ROUND_KEY_s1[118], ROUND_KEY_s0[118]}), .b ({ROUND_KEY_s1[246], ROUND_KEY_s0[246]}), .c ({new_AGEMA_signal_1219, n502}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U544 ( .a ({ROUND_KEY_s1[117], ROUND_KEY_s0[117]}), .b ({ROUND_KEY_s1[245], ROUND_KEY_s0[245]}), .c ({new_AGEMA_signal_1222, n504}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U547 ( .a ({ROUND_KEY_s1[116], ROUND_KEY_s0[116]}), .b ({ROUND_KEY_s1[244], ROUND_KEY_s0[244]}), .c ({new_AGEMA_signal_1225, n506}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U550 ( .a ({ROUND_KEY_s1[115], ROUND_KEY_s0[115]}), .b ({ROUND_KEY_s1[243], ROUND_KEY_s0[243]}), .c ({new_AGEMA_signal_1228, n508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U553 ( .a ({ROUND_KEY_s1[114], ROUND_KEY_s0[114]}), .b ({ROUND_KEY_s1[242], ROUND_KEY_s0[242]}), .c ({new_AGEMA_signal_1231, n510}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U556 ( .a ({ROUND_KEY_s1[113], ROUND_KEY_s0[113]}), .b ({ROUND_KEY_s1[241], ROUND_KEY_s0[241]}), .c ({new_AGEMA_signal_1234, n512}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U559 ( .a ({ROUND_KEY_s1[112], ROUND_KEY_s0[112]}), .b ({ROUND_KEY_s1[240], ROUND_KEY_s0[240]}), .c ({new_AGEMA_signal_1237, n514}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U562 ( .a ({ROUND_KEY_s1[111], ROUND_KEY_s0[111]}), .b ({ROUND_KEY_s1[239], ROUND_KEY_s0[239]}), .c ({new_AGEMA_signal_1240, n516}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U565 ( .a ({ROUND_KEY_s1[110], ROUND_KEY_s0[110]}), .b ({ROUND_KEY_s1[238], ROUND_KEY_s0[238]}), .c ({new_AGEMA_signal_1243, n518}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U568 ( .a ({ROUND_KEY_s1[109], ROUND_KEY_s0[109]}), .b ({ROUND_KEY_s1[237], ROUND_KEY_s0[237]}), .c ({new_AGEMA_signal_1246, n520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U571 ( .a ({ROUND_KEY_s1[108], ROUND_KEY_s0[108]}), .b ({ROUND_KEY_s1[236], ROUND_KEY_s0[236]}), .c ({new_AGEMA_signal_1249, n522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U574 ( .a ({ROUND_KEY_s1[107], ROUND_KEY_s0[107]}), .b ({ROUND_KEY_s1[235], ROUND_KEY_s0[235]}), .c ({new_AGEMA_signal_1252, n524}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U577 ( .a ({ROUND_KEY_s1[106], ROUND_KEY_s0[106]}), .b ({ROUND_KEY_s1[234], ROUND_KEY_s0[234]}), .c ({new_AGEMA_signal_1255, n526}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U580 ( .a ({ROUND_KEY_s1[105], ROUND_KEY_s0[105]}), .b ({ROUND_KEY_s1[233], ROUND_KEY_s0[233]}), .c ({new_AGEMA_signal_1258, n528}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U583 ( .a ({ROUND_KEY_s1[104], ROUND_KEY_s0[104]}), .b ({ROUND_KEY_s1[232], ROUND_KEY_s0[232]}), .c ({new_AGEMA_signal_1261, n530}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U586 ( .a ({ROUND_KEY_s1[103], ROUND_KEY_s0[103]}), .b ({ROUND_KEY_s1[231], ROUND_KEY_s0[231]}), .c ({new_AGEMA_signal_1264, n532}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U589 ( .a ({ROUND_KEY_s1[102], ROUND_KEY_s0[102]}), .b ({ROUND_KEY_s1[230], ROUND_KEY_s0[230]}), .c ({new_AGEMA_signal_1267, n534}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U592 ( .a ({ROUND_KEY_s1[101], ROUND_KEY_s0[101]}), .b ({ROUND_KEY_s1[229], ROUND_KEY_s0[229]}), .c ({new_AGEMA_signal_1270, n536}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U595 ( .a ({ROUND_KEY_s1[100], ROUND_KEY_s0[100]}), .b ({ROUND_KEY_s1[228], ROUND_KEY_s0[228]}), .c ({new_AGEMA_signal_1273, n538}) ) ;
    //ClockGatingController #(8) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U404 ( .a ({ROUND_KEY_s1[354], ROUND_KEY_s0[354]}), .b ({new_AGEMA_signal_1462, CONST_ADDITION[98]}), .c ({new_AGEMA_signal_1483, n407}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U405 ( .a ({new_AGEMA_signal_1087, n408}), .b ({new_AGEMA_signal_1483, n407}), .c ({ROUND_OUT_s1[66], ROUND_OUT_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U416 ( .a ({ROUND_KEY_s1[350], ROUND_KEY_s0[350]}), .b ({new_AGEMA_signal_1461, CONST_ADDITION[94]}), .c ({new_AGEMA_signal_1485, n415}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U417 ( .a ({new_AGEMA_signal_1099, n416}), .b ({new_AGEMA_signal_1485, n415}), .c ({new_AGEMA_signal_1563, SHIFTROWS[86]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U419 ( .a ({ROUND_KEY_s1[349], ROUND_KEY_s0[349]}), .b ({new_AGEMA_signal_1459, CONST_ADDITION[93]}), .c ({new_AGEMA_signal_1487, n417}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U420 ( .a ({new_AGEMA_signal_1102, n418}), .b ({new_AGEMA_signal_1487, n417}), .c ({new_AGEMA_signal_1564, SHIFTROWS[85]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U428 ( .a ({ROUND_KEY_s1[346], ROUND_KEY_s0[346]}), .b ({new_AGEMA_signal_1457, CONST_ADDITION[90]}), .c ({new_AGEMA_signal_1489, n423}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U429 ( .a ({new_AGEMA_signal_1111, n424}), .b ({new_AGEMA_signal_1489, n423}), .c ({new_AGEMA_signal_1565, SHIFTROWS[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U442 ( .a ({ROUND_KEY_s1[342], ROUND_KEY_s0[342]}), .b ({new_AGEMA_signal_1456, CONST_ADDITION[86]}), .c ({new_AGEMA_signal_1491, n433}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U443 ( .a ({new_AGEMA_signal_1123, n434}), .b ({new_AGEMA_signal_1491, n433}), .c ({new_AGEMA_signal_1566, SHIFTROWS[78]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U445 ( .a ({ROUND_KEY_s1[341], ROUND_KEY_s0[341]}), .b ({new_AGEMA_signal_1454, CONST_ADDITION[85]}), .c ({new_AGEMA_signal_1493, n435}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U446 ( .a ({new_AGEMA_signal_1126, n436}), .b ({new_AGEMA_signal_1493, n435}), .c ({new_AGEMA_signal_1567, SHIFTROWS[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U454 ( .a ({ROUND_KEY_s1[338], ROUND_KEY_s0[338]}), .b ({new_AGEMA_signal_1452, CONST_ADDITION[82]}), .c ({new_AGEMA_signal_1495, n441}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U455 ( .a ({new_AGEMA_signal_1135, n442}), .b ({new_AGEMA_signal_1495, n441}), .c ({new_AGEMA_signal_1568, SHIFTROWS[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U466 ( .a ({ROUND_KEY_s1[334], ROUND_KEY_s0[334]}), .b ({new_AGEMA_signal_1451, CONST_ADDITION[78]}), .c ({new_AGEMA_signal_1497, n449}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U467 ( .a ({new_AGEMA_signal_1147, n450}), .b ({new_AGEMA_signal_1497, n449}), .c ({new_AGEMA_signal_1569, SHIFTROWS[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U469 ( .a ({ROUND_KEY_s1[333], ROUND_KEY_s0[333]}), .b ({new_AGEMA_signal_1449, CONST_ADDITION[77]}), .c ({new_AGEMA_signal_1499, n451}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U470 ( .a ({new_AGEMA_signal_1150, n452}), .b ({new_AGEMA_signal_1499, n451}), .c ({new_AGEMA_signal_1570, SHIFTROWS[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U478 ( .a ({ROUND_KEY_s1[330], ROUND_KEY_s0[330]}), .b ({new_AGEMA_signal_1447, CONST_ADDITION[74]}), .c ({new_AGEMA_signal_1501, n457}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U479 ( .a ({new_AGEMA_signal_1159, n458}), .b ({new_AGEMA_signal_1501, n457}), .c ({new_AGEMA_signal_1571, SHIFTROWS[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U490 ( .a ({ROUND_KEY_s1[326], ROUND_KEY_s0[326]}), .b ({new_AGEMA_signal_1446, CONST_ADDITION[70]}), .c ({new_AGEMA_signal_1503, n465}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U491 ( .a ({new_AGEMA_signal_1171, n466}), .b ({new_AGEMA_signal_1503, n465}), .c ({new_AGEMA_signal_1572, SHIFTROWS[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U493 ( .a ({ROUND_KEY_s1[325], ROUND_KEY_s0[325]}), .b ({new_AGEMA_signal_1444, CONST_ADDITION[69]}), .c ({new_AGEMA_signal_1505, n467}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U494 ( .a ({new_AGEMA_signal_1174, n468}), .b ({new_AGEMA_signal_1505, n467}), .c ({new_AGEMA_signal_1573, SHIFTROWS[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U502 ( .a ({ROUND_KEY_s1[322], ROUND_KEY_s0[322]}), .b ({new_AGEMA_signal_1442, CONST_ADDITION[66]}), .c ({new_AGEMA_signal_1507, n473}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U503 ( .a ({new_AGEMA_signal_1183, n474}), .b ({new_AGEMA_signal_1507, n473}), .c ({new_AGEMA_signal_1574, SHIFTROWS[90]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U514 ( .a ({ROUND_KEY_s1[382], ROUND_KEY_s0[382]}), .b ({new_AGEMA_signal_1481, CONST_ADDITION[126]}), .c ({new_AGEMA_signal_1509, n481}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U515 ( .a ({new_AGEMA_signal_1195, n482}), .b ({new_AGEMA_signal_1509, n481}), .c ({ROUND_OUT_s1[94], ROUND_OUT_s0[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U517 ( .a ({ROUND_KEY_s1[381], ROUND_KEY_s0[381]}), .b ({new_AGEMA_signal_1479, CONST_ADDITION[125]}), .c ({new_AGEMA_signal_1511, n483}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U518 ( .a ({new_AGEMA_signal_1198, n484}), .b ({new_AGEMA_signal_1511, n483}), .c ({ROUND_OUT_s1[93], ROUND_OUT_s0[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U527 ( .a ({new_AGEMA_signal_1477, SUBSTITUTION[122]}), .b ({ROUND_KEY_s1[378], ROUND_KEY_s0[378]}), .c ({new_AGEMA_signal_1513, n490}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U528 ( .a ({new_AGEMA_signal_1207, n491}), .b ({new_AGEMA_signal_1513, n490}), .c ({new_AGEMA_signal_1577, n492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U529 ( .a ({1'b0, CONST_IN[2]}), .b ({new_AGEMA_signal_1577, n492}), .c ({ROUND_OUT_s1[90], ROUND_OUT_s0[90]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U542 ( .a ({ROUND_KEY_s1[374], ROUND_KEY_s0[374]}), .b ({new_AGEMA_signal_1476, CONST_ADDITION[118]}), .c ({new_AGEMA_signal_1515, n501}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U543 ( .a ({new_AGEMA_signal_1219, n502}), .b ({new_AGEMA_signal_1515, n501}), .c ({ROUND_OUT_s1[86], ROUND_OUT_s0[86]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U545 ( .a ({ROUND_KEY_s1[373], ROUND_KEY_s0[373]}), .b ({new_AGEMA_signal_1474, CONST_ADDITION[117]}), .c ({new_AGEMA_signal_1517, n503}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U546 ( .a ({new_AGEMA_signal_1222, n504}), .b ({new_AGEMA_signal_1517, n503}), .c ({ROUND_OUT_s1[85], ROUND_OUT_s0[85]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U554 ( .a ({ROUND_KEY_s1[370], ROUND_KEY_s0[370]}), .b ({new_AGEMA_signal_1472, CONST_ADDITION[114]}), .c ({new_AGEMA_signal_1519, n509}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U555 ( .a ({new_AGEMA_signal_1231, n510}), .b ({new_AGEMA_signal_1519, n509}), .c ({ROUND_OUT_s1[82], ROUND_OUT_s0[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U566 ( .a ({ROUND_KEY_s1[366], ROUND_KEY_s0[366]}), .b ({new_AGEMA_signal_1471, CONST_ADDITION[110]}), .c ({new_AGEMA_signal_1521, n517}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U567 ( .a ({new_AGEMA_signal_1243, n518}), .b ({new_AGEMA_signal_1521, n517}), .c ({ROUND_OUT_s1[78], ROUND_OUT_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U569 ( .a ({ROUND_KEY_s1[365], ROUND_KEY_s0[365]}), .b ({new_AGEMA_signal_1469, CONST_ADDITION[109]}), .c ({new_AGEMA_signal_1523, n519}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U570 ( .a ({new_AGEMA_signal_1246, n520}), .b ({new_AGEMA_signal_1523, n519}), .c ({ROUND_OUT_s1[77], ROUND_OUT_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U578 ( .a ({ROUND_KEY_s1[362], ROUND_KEY_s0[362]}), .b ({new_AGEMA_signal_1467, CONST_ADDITION[106]}), .c ({new_AGEMA_signal_1525, n525}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U579 ( .a ({new_AGEMA_signal_1255, n526}), .b ({new_AGEMA_signal_1525, n525}), .c ({ROUND_OUT_s1[74], ROUND_OUT_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U590 ( .a ({ROUND_KEY_s1[358], ROUND_KEY_s0[358]}), .b ({new_AGEMA_signal_1466, CONST_ADDITION[102]}), .c ({new_AGEMA_signal_1527, n533}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U591 ( .a ({new_AGEMA_signal_1267, n534}), .b ({new_AGEMA_signal_1527, n533}), .c ({ROUND_OUT_s1[70], ROUND_OUT_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U593 ( .a ({ROUND_KEY_s1[357], ROUND_KEY_s0[357]}), .b ({new_AGEMA_signal_1464, CONST_ADDITION[101]}), .c ({new_AGEMA_signal_1529, n535}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U594 ( .a ({new_AGEMA_signal_1270, n536}), .b ({new_AGEMA_signal_1529, n535}), .c ({ROUND_OUT_s1[69], ROUND_OUT_s0[69]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_0_U6 ( .a ({new_AGEMA_signal_1281, S_0_R1[1]}), .b ({ROUND_IN_s1[6], ROUND_IN_s0[6]}), .c ({new_AGEMA_signal_1402, SHIFTROWS[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_0_U3 ( .a ({new_AGEMA_signal_1279, S_0_R2[0]}), .b ({ROUND_IN_s1[0], ROUND_IN_s0[0]}), .c ({new_AGEMA_signal_1404, SHIFTROWS[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_0_U2 ( .a ({new_AGEMA_signal_1276, S_0_R1[0]}), .b ({ROUND_IN_s1[4], ROUND_IN_s0[4]}), .c ({new_AGEMA_signal_1406, SHIFTROWS[14]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_0_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[6], ROUND_IN_s0[6]}), .b ({ROUND_IN_s1[7], ROUND_IN_s0[7]}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_1276, S_0_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_0_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[2], ROUND_IN_s0[2]}), .b ({ROUND_IN_s1[3], ROUND_IN_s0[3]}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_1279, S_0_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_0_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[1], ROUND_IN_s0[1]}), .b ({ROUND_IN_s1[2], ROUND_IN_s0[2]}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_1281, S_0_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_1_U6 ( .a ({new_AGEMA_signal_1289, S_1_R1[1]}), .b ({ROUND_IN_s1[14], ROUND_IN_s0[14]}), .c ({new_AGEMA_signal_1407, SHIFTROWS[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_1_U3 ( .a ({new_AGEMA_signal_1287, S_1_R2[0]}), .b ({ROUND_IN_s1[8], ROUND_IN_s0[8]}), .c ({new_AGEMA_signal_1409, SHIFTROWS[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_1_U2 ( .a ({new_AGEMA_signal_1284, S_1_R1[0]}), .b ({ROUND_IN_s1[12], ROUND_IN_s0[12]}), .c ({new_AGEMA_signal_1411, SHIFTROWS[22]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_1_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[14], ROUND_IN_s0[14]}), .b ({ROUND_IN_s1[15], ROUND_IN_s0[15]}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_1284, S_1_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_1_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[10], ROUND_IN_s0[10]}), .b ({ROUND_IN_s1[11], ROUND_IN_s0[11]}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_1287, S_1_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_1_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[9], ROUND_IN_s0[9]}), .b ({ROUND_IN_s1[10], ROUND_IN_s0[10]}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_1289, S_1_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_2_U6 ( .a ({new_AGEMA_signal_1297, S_2_R1[1]}), .b ({ROUND_IN_s1[22], ROUND_IN_s0[22]}), .c ({new_AGEMA_signal_1412, SHIFTROWS[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_2_U3 ( .a ({new_AGEMA_signal_1295, S_2_R2[0]}), .b ({ROUND_IN_s1[16], ROUND_IN_s0[16]}), .c ({new_AGEMA_signal_1414, SHIFTROWS[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_2_U2 ( .a ({new_AGEMA_signal_1292, S_2_R1[0]}), .b ({ROUND_IN_s1[20], ROUND_IN_s0[20]}), .c ({new_AGEMA_signal_1416, SHIFTROWS[30]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_2_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[22], ROUND_IN_s0[22]}), .b ({ROUND_IN_s1[23], ROUND_IN_s0[23]}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_1292, S_2_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_2_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[18], ROUND_IN_s0[18]}), .b ({ROUND_IN_s1[19], ROUND_IN_s0[19]}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_1295, S_2_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_2_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[17], ROUND_IN_s0[17]}), .b ({ROUND_IN_s1[18], ROUND_IN_s0[18]}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_1297, S_2_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_3_U6 ( .a ({new_AGEMA_signal_1305, S_3_R1[1]}), .b ({ROUND_IN_s1[30], ROUND_IN_s0[30]}), .c ({new_AGEMA_signal_1417, SHIFTROWS[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_3_U3 ( .a ({new_AGEMA_signal_1303, S_3_R2[0]}), .b ({ROUND_IN_s1[24], ROUND_IN_s0[24]}), .c ({new_AGEMA_signal_1419, SHIFTROWS[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_3_U2 ( .a ({new_AGEMA_signal_1300, S_3_R1[0]}), .b ({ROUND_IN_s1[28], ROUND_IN_s0[28]}), .c ({new_AGEMA_signal_1421, SHIFTROWS[6]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_3_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[30], ROUND_IN_s0[30]}), .b ({ROUND_IN_s1[31], ROUND_IN_s0[31]}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_1300, S_3_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_3_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[26], ROUND_IN_s0[26]}), .b ({ROUND_IN_s1[27], ROUND_IN_s0[27]}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_1303, S_3_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_3_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[25], ROUND_IN_s0[25]}), .b ({ROUND_IN_s1[26], ROUND_IN_s0[26]}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_1305, S_3_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_4_U6 ( .a ({new_AGEMA_signal_1313, S_4_R1[1]}), .b ({ROUND_IN_s1[38], ROUND_IN_s0[38]}), .c ({new_AGEMA_signal_1422, SHIFTROWS[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_4_U3 ( .a ({new_AGEMA_signal_1311, S_4_R2[0]}), .b ({ROUND_IN_s1[32], ROUND_IN_s0[32]}), .c ({new_AGEMA_signal_1424, SHIFTROWS[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_4_U2 ( .a ({new_AGEMA_signal_1308, S_4_R1[0]}), .b ({ROUND_IN_s1[36], ROUND_IN_s0[36]}), .c ({new_AGEMA_signal_1426, SHIFTROWS[54]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_4_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[38], ROUND_IN_s0[38]}), .b ({ROUND_IN_s1[39], ROUND_IN_s0[39]}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_1308, S_4_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_4_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[34], ROUND_IN_s0[34]}), .b ({ROUND_IN_s1[35], ROUND_IN_s0[35]}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_1311, S_4_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_4_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[33], ROUND_IN_s0[33]}), .b ({ROUND_IN_s1[34], ROUND_IN_s0[34]}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_1313, S_4_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_5_U6 ( .a ({new_AGEMA_signal_1321, S_5_R1[1]}), .b ({ROUND_IN_s1[46], ROUND_IN_s0[46]}), .c ({new_AGEMA_signal_1427, SHIFTROWS[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_5_U3 ( .a ({new_AGEMA_signal_1319, S_5_R2[0]}), .b ({ROUND_IN_s1[40], ROUND_IN_s0[40]}), .c ({new_AGEMA_signal_1429, SHIFTROWS[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_5_U2 ( .a ({new_AGEMA_signal_1316, S_5_R1[0]}), .b ({ROUND_IN_s1[44], ROUND_IN_s0[44]}), .c ({new_AGEMA_signal_1431, SHIFTROWS[62]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_5_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[46], ROUND_IN_s0[46]}), .b ({ROUND_IN_s1[47], ROUND_IN_s0[47]}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_1316, S_5_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_5_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[42], ROUND_IN_s0[42]}), .b ({ROUND_IN_s1[43], ROUND_IN_s0[43]}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_1319, S_5_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_5_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[41], ROUND_IN_s0[41]}), .b ({ROUND_IN_s1[42], ROUND_IN_s0[42]}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_1321, S_5_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_6_U6 ( .a ({new_AGEMA_signal_1329, S_6_R1[1]}), .b ({ROUND_IN_s1[54], ROUND_IN_s0[54]}), .c ({new_AGEMA_signal_1432, SHIFTROWS[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_6_U3 ( .a ({new_AGEMA_signal_1327, S_6_R2[0]}), .b ({ROUND_IN_s1[48], ROUND_IN_s0[48]}), .c ({new_AGEMA_signal_1434, SHIFTROWS[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_6_U2 ( .a ({new_AGEMA_signal_1324, S_6_R1[0]}), .b ({ROUND_IN_s1[52], ROUND_IN_s0[52]}), .c ({new_AGEMA_signal_1436, SHIFTROWS[38]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_6_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[54], ROUND_IN_s0[54]}), .b ({ROUND_IN_s1[55], ROUND_IN_s0[55]}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_1324, S_6_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_6_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[50], ROUND_IN_s0[50]}), .b ({ROUND_IN_s1[51], ROUND_IN_s0[51]}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_1327, S_6_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_6_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[49], ROUND_IN_s0[49]}), .b ({ROUND_IN_s1[50], ROUND_IN_s0[50]}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_1329, S_6_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_7_U6 ( .a ({new_AGEMA_signal_1337, S_7_R1[1]}), .b ({ROUND_IN_s1[62], ROUND_IN_s0[62]}), .c ({new_AGEMA_signal_1437, SHIFTROWS[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_7_U3 ( .a ({new_AGEMA_signal_1335, S_7_R2[0]}), .b ({ROUND_IN_s1[56], ROUND_IN_s0[56]}), .c ({new_AGEMA_signal_1439, SHIFTROWS[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_7_U2 ( .a ({new_AGEMA_signal_1332, S_7_R1[0]}), .b ({ROUND_IN_s1[60], ROUND_IN_s0[60]}), .c ({new_AGEMA_signal_1441, SHIFTROWS[46]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_7_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[62], ROUND_IN_s0[62]}), .b ({ROUND_IN_s1[63], ROUND_IN_s0[63]}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_1332, S_7_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_7_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[58], ROUND_IN_s0[58]}), .b ({ROUND_IN_s1[59], ROUND_IN_s0[59]}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_1335, S_7_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_7_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[57], ROUND_IN_s0[57]}), .b ({ROUND_IN_s1[58], ROUND_IN_s0[58]}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_1337, S_7_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_8_U6 ( .a ({new_AGEMA_signal_1345, S_8_R1[1]}), .b ({ROUND_IN_s1[70], ROUND_IN_s0[70]}), .c ({new_AGEMA_signal_1442, CONST_ADDITION[66]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_8_U3 ( .a ({new_AGEMA_signal_1343, S_8_R2[0]}), .b ({ROUND_IN_s1[64], ROUND_IN_s0[64]}), .c ({new_AGEMA_signal_1444, CONST_ADDITION[69]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_8_U2 ( .a ({new_AGEMA_signal_1340, S_8_R1[0]}), .b ({ROUND_IN_s1[68], ROUND_IN_s0[68]}), .c ({new_AGEMA_signal_1446, CONST_ADDITION[70]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_8_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[70], ROUND_IN_s0[70]}), .b ({ROUND_IN_s1[71], ROUND_IN_s0[71]}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_1340, S_8_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_8_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[66], ROUND_IN_s0[66]}), .b ({ROUND_IN_s1[67], ROUND_IN_s0[67]}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_1343, S_8_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_8_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[65], ROUND_IN_s0[65]}), .b ({ROUND_IN_s1[66], ROUND_IN_s0[66]}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_1345, S_8_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_9_U6 ( .a ({new_AGEMA_signal_1353, S_9_R1[1]}), .b ({ROUND_IN_s1[78], ROUND_IN_s0[78]}), .c ({new_AGEMA_signal_1447, CONST_ADDITION[74]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_9_U3 ( .a ({new_AGEMA_signal_1351, S_9_R2[0]}), .b ({ROUND_IN_s1[72], ROUND_IN_s0[72]}), .c ({new_AGEMA_signal_1449, CONST_ADDITION[77]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_9_U2 ( .a ({new_AGEMA_signal_1348, S_9_R1[0]}), .b ({ROUND_IN_s1[76], ROUND_IN_s0[76]}), .c ({new_AGEMA_signal_1451, CONST_ADDITION[78]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_9_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[78], ROUND_IN_s0[78]}), .b ({ROUND_IN_s1[79], ROUND_IN_s0[79]}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_1348, S_9_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_9_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[74], ROUND_IN_s0[74]}), .b ({ROUND_IN_s1[75], ROUND_IN_s0[75]}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_1351, S_9_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_9_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[73], ROUND_IN_s0[73]}), .b ({ROUND_IN_s1[74], ROUND_IN_s0[74]}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_1353, S_9_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_10_U6 ( .a ({new_AGEMA_signal_1361, S_10_R1[1]}), .b ({ROUND_IN_s1[86], ROUND_IN_s0[86]}), .c ({new_AGEMA_signal_1452, CONST_ADDITION[82]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_10_U3 ( .a ({new_AGEMA_signal_1359, S_10_R2[0]}), .b ({ROUND_IN_s1[80], ROUND_IN_s0[80]}), .c ({new_AGEMA_signal_1454, CONST_ADDITION[85]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_10_U2 ( .a ({new_AGEMA_signal_1356, S_10_R1[0]}), .b ({ROUND_IN_s1[84], ROUND_IN_s0[84]}), .c ({new_AGEMA_signal_1456, CONST_ADDITION[86]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_10_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[86], ROUND_IN_s0[86]}), .b ({ROUND_IN_s1[87], ROUND_IN_s0[87]}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_1356, S_10_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_10_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[82], ROUND_IN_s0[82]}), .b ({ROUND_IN_s1[83], ROUND_IN_s0[83]}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_1359, S_10_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_10_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[81], ROUND_IN_s0[81]}), .b ({ROUND_IN_s1[82], ROUND_IN_s0[82]}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_1361, S_10_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_11_U6 ( .a ({new_AGEMA_signal_1369, S_11_R1[1]}), .b ({ROUND_IN_s1[94], ROUND_IN_s0[94]}), .c ({new_AGEMA_signal_1457, CONST_ADDITION[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_11_U3 ( .a ({new_AGEMA_signal_1367, S_11_R2[0]}), .b ({ROUND_IN_s1[88], ROUND_IN_s0[88]}), .c ({new_AGEMA_signal_1459, CONST_ADDITION[93]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_11_U2 ( .a ({new_AGEMA_signal_1364, S_11_R1[0]}), .b ({ROUND_IN_s1[92], ROUND_IN_s0[92]}), .c ({new_AGEMA_signal_1461, CONST_ADDITION[94]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_11_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[94], ROUND_IN_s0[94]}), .b ({ROUND_IN_s1[95], ROUND_IN_s0[95]}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_1364, S_11_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_11_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[90], ROUND_IN_s0[90]}), .b ({ROUND_IN_s1[91], ROUND_IN_s0[91]}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_1367, S_11_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_11_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[89], ROUND_IN_s0[89]}), .b ({ROUND_IN_s1[90], ROUND_IN_s0[90]}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_1369, S_11_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_12_U6 ( .a ({new_AGEMA_signal_1377, S_12_R1[1]}), .b ({ROUND_IN_s1[102], ROUND_IN_s0[102]}), .c ({new_AGEMA_signal_1462, CONST_ADDITION[98]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_12_U3 ( .a ({new_AGEMA_signal_1375, S_12_R2[0]}), .b ({ROUND_IN_s1[96], ROUND_IN_s0[96]}), .c ({new_AGEMA_signal_1464, CONST_ADDITION[101]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_12_U2 ( .a ({new_AGEMA_signal_1372, S_12_R1[0]}), .b ({ROUND_IN_s1[100], ROUND_IN_s0[100]}), .c ({new_AGEMA_signal_1466, CONST_ADDITION[102]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_12_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[102], ROUND_IN_s0[102]}), .b ({ROUND_IN_s1[103], ROUND_IN_s0[103]}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_1372, S_12_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_12_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[98], ROUND_IN_s0[98]}), .b ({ROUND_IN_s1[99], ROUND_IN_s0[99]}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_1375, S_12_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_12_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[97], ROUND_IN_s0[97]}), .b ({ROUND_IN_s1[98], ROUND_IN_s0[98]}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_1377, S_12_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_13_U6 ( .a ({new_AGEMA_signal_1385, S_13_R1[1]}), .b ({ROUND_IN_s1[110], ROUND_IN_s0[110]}), .c ({new_AGEMA_signal_1467, CONST_ADDITION[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_13_U3 ( .a ({new_AGEMA_signal_1383, S_13_R2[0]}), .b ({ROUND_IN_s1[104], ROUND_IN_s0[104]}), .c ({new_AGEMA_signal_1469, CONST_ADDITION[109]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_13_U2 ( .a ({new_AGEMA_signal_1380, S_13_R1[0]}), .b ({ROUND_IN_s1[108], ROUND_IN_s0[108]}), .c ({new_AGEMA_signal_1471, CONST_ADDITION[110]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_13_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[110], ROUND_IN_s0[110]}), .b ({ROUND_IN_s1[111], ROUND_IN_s0[111]}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_1380, S_13_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_13_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[106], ROUND_IN_s0[106]}), .b ({ROUND_IN_s1[107], ROUND_IN_s0[107]}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_1383, S_13_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_13_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[105], ROUND_IN_s0[105]}), .b ({ROUND_IN_s1[106], ROUND_IN_s0[106]}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_1385, S_13_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_14_U6 ( .a ({new_AGEMA_signal_1393, S_14_R1[1]}), .b ({ROUND_IN_s1[118], ROUND_IN_s0[118]}), .c ({new_AGEMA_signal_1472, CONST_ADDITION[114]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_14_U3 ( .a ({new_AGEMA_signal_1391, S_14_R2[0]}), .b ({ROUND_IN_s1[112], ROUND_IN_s0[112]}), .c ({new_AGEMA_signal_1474, CONST_ADDITION[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_14_U2 ( .a ({new_AGEMA_signal_1388, S_14_R1[0]}), .b ({ROUND_IN_s1[116], ROUND_IN_s0[116]}), .c ({new_AGEMA_signal_1476, CONST_ADDITION[118]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_14_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[118], ROUND_IN_s0[118]}), .b ({ROUND_IN_s1[119], ROUND_IN_s0[119]}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_1388, S_14_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_14_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[114], ROUND_IN_s0[114]}), .b ({ROUND_IN_s1[115], ROUND_IN_s0[115]}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_1391, S_14_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_14_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[113], ROUND_IN_s0[113]}), .b ({ROUND_IN_s1[114], ROUND_IN_s0[114]}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_1393, S_14_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_15_U6 ( .a ({new_AGEMA_signal_1401, S_15_R1[1]}), .b ({ROUND_IN_s1[126], ROUND_IN_s0[126]}), .c ({new_AGEMA_signal_1477, SUBSTITUTION[122]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_15_U3 ( .a ({new_AGEMA_signal_1399, S_15_R2[0]}), .b ({ROUND_IN_s1[120], ROUND_IN_s0[120]}), .c ({new_AGEMA_signal_1479, CONST_ADDITION[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_15_U2 ( .a ({new_AGEMA_signal_1396, S_15_R1[0]}), .b ({ROUND_IN_s1[124], ROUND_IN_s0[124]}), .c ({new_AGEMA_signal_1481, CONST_ADDITION[126]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_15_NOR1Inst_0_U1 ( .a ({ROUND_IN_s1[126], ROUND_IN_s0[126]}), .b ({ROUND_IN_s1[127], ROUND_IN_s0[127]}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_1396, S_15_R1[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_15_NOR2Inst_0_U1 ( .a ({ROUND_IN_s1[122], ROUND_IN_s0[122]}), .b ({ROUND_IN_s1[123], ROUND_IN_s0[123]}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_1399, S_15_R2[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_15_NOR1Inst_1_U1 ( .a ({ROUND_IN_s1[121], ROUND_IN_s0[121]}), .b ({ROUND_IN_s1[122], ROUND_IN_s0[122]}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_1401, S_15_R1[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U92 ( .a ({new_AGEMA_signal_1416, SHIFTROWS[30]}), .b ({ROUND_OUT_s1[30], ROUND_OUT_s0[30]}), .c ({ROUND_OUT_s1[126], ROUND_OUT_s0[126]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U91 ( .a ({ROUND_OUT_s1[94], ROUND_OUT_s0[94]}), .b ({new_AGEMA_signal_1431, SHIFTROWS[62]}), .c ({ROUND_OUT_s1[30], ROUND_OUT_s0[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U80 ( .a ({new_AGEMA_signal_1406, SHIFTROWS[14]}), .b ({ROUND_OUT_s1[14], ROUND_OUT_s0[14]}), .c ({ROUND_OUT_s1[110], ROUND_OUT_s0[110]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U79 ( .a ({ROUND_OUT_s1[78], ROUND_OUT_s0[78]}), .b ({new_AGEMA_signal_1441, SHIFTROWS[46]}), .c ({ROUND_OUT_s1[14], ROUND_OUT_s0[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U78 ( .a ({new_AGEMA_signal_1404, SHIFTROWS[13]}), .b ({ROUND_OUT_s1[13], ROUND_OUT_s0[13]}), .c ({ROUND_OUT_s1[109], ROUND_OUT_s0[109]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U77 ( .a ({ROUND_OUT_s1[77], ROUND_OUT_s0[77]}), .b ({new_AGEMA_signal_1439, SHIFTROWS[45]}), .c ({ROUND_OUT_s1[13], ROUND_OUT_s0[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U74 ( .a ({new_AGEMA_signal_1411, SHIFTROWS[22]}), .b ({ROUND_OUT_s1[22], ROUND_OUT_s0[22]}), .c ({ROUND_OUT_s1[118], ROUND_OUT_s0[118]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U73 ( .a ({ROUND_OUT_s1[86], ROUND_OUT_s0[86]}), .b ({new_AGEMA_signal_1426, SHIFTROWS[54]}), .c ({ROUND_OUT_s1[22], ROUND_OUT_s0[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U68 ( .a ({new_AGEMA_signal_1409, SHIFTROWS[21]}), .b ({ROUND_OUT_s1[21], ROUND_OUT_s0[21]}), .c ({ROUND_OUT_s1[117], ROUND_OUT_s0[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U67 ( .a ({ROUND_OUT_s1[85], ROUND_OUT_s0[85]}), .b ({new_AGEMA_signal_1424, SHIFTROWS[53]}), .c ({ROUND_OUT_s1[21], ROUND_OUT_s0[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U66 ( .a ({new_AGEMA_signal_1402, SHIFTROWS[10]}), .b ({ROUND_OUT_s1[10], ROUND_OUT_s0[10]}), .c ({ROUND_OUT_s1[106], ROUND_OUT_s0[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U65 ( .a ({ROUND_OUT_s1[74], ROUND_OUT_s0[74]}), .b ({new_AGEMA_signal_1437, SHIFTROWS[42]}), .c ({ROUND_OUT_s1[10], ROUND_OUT_s0[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U62 ( .a ({new_AGEMA_signal_1414, SHIFTROWS[29]}), .b ({ROUND_OUT_s1[29], ROUND_OUT_s0[29]}), .c ({ROUND_OUT_s1[125], ROUND_OUT_s0[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U61 ( .a ({ROUND_OUT_s1[93], ROUND_OUT_s0[93]}), .b ({new_AGEMA_signal_1429, SHIFTROWS[61]}), .c ({ROUND_OUT_s1[29], ROUND_OUT_s0[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U60 ( .a ({new_AGEMA_signal_1412, SHIFTROWS[26]}), .b ({ROUND_OUT_s1[26], ROUND_OUT_s0[26]}), .c ({ROUND_OUT_s1[122], ROUND_OUT_s0[122]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U59 ( .a ({ROUND_OUT_s1[90], ROUND_OUT_s0[90]}), .b ({new_AGEMA_signal_1427, SHIFTROWS[58]}), .c ({ROUND_OUT_s1[26], ROUND_OUT_s0[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U50 ( .a ({new_AGEMA_signal_1421, SHIFTROWS[6]}), .b ({ROUND_OUT_s1[6], ROUND_OUT_s0[6]}), .c ({ROUND_OUT_s1[102], ROUND_OUT_s0[102]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U49 ( .a ({ROUND_OUT_s1[70], ROUND_OUT_s0[70]}), .b ({new_AGEMA_signal_1436, SHIFTROWS[38]}), .c ({ROUND_OUT_s1[6], ROUND_OUT_s0[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U48 ( .a ({new_AGEMA_signal_1419, SHIFTROWS[5]}), .b ({ROUND_OUT_s1[5], ROUND_OUT_s0[5]}), .c ({ROUND_OUT_s1[101], ROUND_OUT_s0[101]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U47 ( .a ({ROUND_OUT_s1[69], ROUND_OUT_s0[69]}), .b ({new_AGEMA_signal_1434, SHIFTROWS[37]}), .c ({ROUND_OUT_s1[5], ROUND_OUT_s0[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U44 ( .a ({new_AGEMA_signal_1407, SHIFTROWS[18]}), .b ({ROUND_OUT_s1[18], ROUND_OUT_s0[18]}), .c ({ROUND_OUT_s1[114], ROUND_OUT_s0[114]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U43 ( .a ({ROUND_OUT_s1[82], ROUND_OUT_s0[82]}), .b ({new_AGEMA_signal_1422, SHIFTROWS[50]}), .c ({ROUND_OUT_s1[18], ROUND_OUT_s0[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U36 ( .a ({new_AGEMA_signal_1417, SHIFTROWS[2]}), .b ({ROUND_OUT_s1[2], ROUND_OUT_s0[2]}), .c ({ROUND_OUT_s1[98], ROUND_OUT_s0[98]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U35 ( .a ({ROUND_OUT_s1[66], ROUND_OUT_s0[66]}), .b ({new_AGEMA_signal_1432, SHIFTROWS[34]}), .c ({ROUND_OUT_s1[2], ROUND_OUT_s0[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U30 ( .a ({new_AGEMA_signal_1432, SHIFTROWS[34]}), .b ({new_AGEMA_signal_1571, SHIFTROWS[66]}), .c ({ROUND_OUT_s1[34], ROUND_OUT_s0[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U27 ( .a ({new_AGEMA_signal_1434, SHIFTROWS[37]}), .b ({new_AGEMA_signal_1570, SHIFTROWS[69]}), .c ({ROUND_OUT_s1[37], ROUND_OUT_s0[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U26 ( .a ({new_AGEMA_signal_1436, SHIFTROWS[38]}), .b ({new_AGEMA_signal_1569, SHIFTROWS[70]}), .c ({ROUND_OUT_s1[38], ROUND_OUT_s0[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U22 ( .a ({new_AGEMA_signal_1437, SHIFTROWS[42]}), .b ({new_AGEMA_signal_1568, SHIFTROWS[74]}), .c ({ROUND_OUT_s1[42], ROUND_OUT_s0[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U19 ( .a ({new_AGEMA_signal_1439, SHIFTROWS[45]}), .b ({new_AGEMA_signal_1567, SHIFTROWS[77]}), .c ({ROUND_OUT_s1[45], ROUND_OUT_s0[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U18 ( .a ({new_AGEMA_signal_1441, SHIFTROWS[46]}), .b ({new_AGEMA_signal_1566, SHIFTROWS[78]}), .c ({ROUND_OUT_s1[46], ROUND_OUT_s0[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U14 ( .a ({new_AGEMA_signal_1422, SHIFTROWS[50]}), .b ({new_AGEMA_signal_1565, SHIFTROWS[82]}), .c ({ROUND_OUT_s1[50], ROUND_OUT_s0[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U11 ( .a ({new_AGEMA_signal_1424, SHIFTROWS[53]}), .b ({new_AGEMA_signal_1564, SHIFTROWS[85]}), .c ({ROUND_OUT_s1[53], ROUND_OUT_s0[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U10 ( .a ({new_AGEMA_signal_1426, SHIFTROWS[54]}), .b ({new_AGEMA_signal_1563, SHIFTROWS[86]}), .c ({ROUND_OUT_s1[54], ROUND_OUT_s0[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U6 ( .a ({new_AGEMA_signal_1427, SHIFTROWS[58]}), .b ({new_AGEMA_signal_1574, SHIFTROWS[90]}), .c ({ROUND_OUT_s1[58], ROUND_OUT_s0[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U3 ( .a ({new_AGEMA_signal_1429, SHIFTROWS[61]}), .b ({new_AGEMA_signal_1573, SHIFTROWS[93]}), .c ({ROUND_OUT_s1[61], ROUND_OUT_s0[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U2 ( .a ({new_AGEMA_signal_1431, SHIFTROWS[62]}), .b ({new_AGEMA_signal_1572, SHIFTROWS[94]}), .c ({ROUND_OUT_s1[62], ROUND_OUT_s0[62]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U401 ( .a ({ROUND_KEY_s1[355], ROUND_KEY_s0[355]}), .b ({new_AGEMA_signal_1622, CONST_ADDITION[99]}), .c ({new_AGEMA_signal_1635, n405}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U402 ( .a ({new_AGEMA_signal_1084, n406}), .b ({new_AGEMA_signal_1635, n405}), .c ({ROUND_OUT_s1[67], ROUND_OUT_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U413 ( .a ({ROUND_KEY_s1[351], ROUND_KEY_s0[351]}), .b ({new_AGEMA_signal_1621, CONST_ADDITION[95]}), .c ({new_AGEMA_signal_1637, n413}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U414 ( .a ({new_AGEMA_signal_1096, n414}), .b ({new_AGEMA_signal_1637, n413}), .c ({new_AGEMA_signal_1723, SHIFTROWS[87]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U425 ( .a ({ROUND_KEY_s1[347], ROUND_KEY_s0[347]}), .b ({new_AGEMA_signal_1619, CONST_ADDITION[91]}), .c ({new_AGEMA_signal_1639, n421}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U426 ( .a ({new_AGEMA_signal_1108, n422}), .b ({new_AGEMA_signal_1639, n421}), .c ({new_AGEMA_signal_1724, SHIFTROWS[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U439 ( .a ({ROUND_KEY_s1[343], ROUND_KEY_s0[343]}), .b ({new_AGEMA_signal_1618, CONST_ADDITION[87]}), .c ({new_AGEMA_signal_1641, n431}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U440 ( .a ({new_AGEMA_signal_1120, n432}), .b ({new_AGEMA_signal_1641, n431}), .c ({new_AGEMA_signal_1725, SHIFTROWS[79]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U451 ( .a ({ROUND_KEY_s1[339], ROUND_KEY_s0[339]}), .b ({new_AGEMA_signal_1616, CONST_ADDITION[83]}), .c ({new_AGEMA_signal_1643, n439}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U452 ( .a ({new_AGEMA_signal_1132, n440}), .b ({new_AGEMA_signal_1643, n439}), .c ({new_AGEMA_signal_1726, SHIFTROWS[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U463 ( .a ({ROUND_KEY_s1[335], ROUND_KEY_s0[335]}), .b ({new_AGEMA_signal_1615, CONST_ADDITION[79]}), .c ({new_AGEMA_signal_1645, n447}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U464 ( .a ({new_AGEMA_signal_1144, n448}), .b ({new_AGEMA_signal_1645, n447}), .c ({new_AGEMA_signal_1727, SHIFTROWS[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U475 ( .a ({ROUND_KEY_s1[331], ROUND_KEY_s0[331]}), .b ({new_AGEMA_signal_1613, CONST_ADDITION[75]}), .c ({new_AGEMA_signal_1647, n455}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U476 ( .a ({new_AGEMA_signal_1156, n456}), .b ({new_AGEMA_signal_1647, n455}), .c ({new_AGEMA_signal_1728, SHIFTROWS[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U487 ( .a ({ROUND_KEY_s1[327], ROUND_KEY_s0[327]}), .b ({new_AGEMA_signal_1612, CONST_ADDITION[71]}), .c ({new_AGEMA_signal_1649, n463}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U488 ( .a ({new_AGEMA_signal_1168, n464}), .b ({new_AGEMA_signal_1649, n463}), .c ({new_AGEMA_signal_1729, SHIFTROWS[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U499 ( .a ({ROUND_KEY_s1[323], ROUND_KEY_s0[323]}), .b ({new_AGEMA_signal_1610, CONST_ADDITION[67]}), .c ({new_AGEMA_signal_1651, n471}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U500 ( .a ({new_AGEMA_signal_1180, n472}), .b ({new_AGEMA_signal_1651, n471}), .c ({new_AGEMA_signal_1730, SHIFTROWS[91]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U511 ( .a ({ROUND_KEY_s1[383], ROUND_KEY_s0[383]}), .b ({new_AGEMA_signal_1633, CONST_ADDITION[127]}), .c ({new_AGEMA_signal_1653, n479}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U512 ( .a ({new_AGEMA_signal_1192, n480}), .b ({new_AGEMA_signal_1653, n479}), .c ({ROUND_OUT_s1[95], ROUND_OUT_s0[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U523 ( .a ({new_AGEMA_signal_1631, SUBSTITUTION[123]}), .b ({ROUND_KEY_s1[379], ROUND_KEY_s0[379]}), .c ({new_AGEMA_signal_1655, n487}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U524 ( .a ({new_AGEMA_signal_1204, n488}), .b ({new_AGEMA_signal_1655, n487}), .c ({new_AGEMA_signal_1732, n489}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U525 ( .a ({1'b0, CONST_IN[3]}), .b ({new_AGEMA_signal_1732, n489}), .c ({ROUND_OUT_s1[91], ROUND_OUT_s0[91]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U539 ( .a ({ROUND_KEY_s1[375], ROUND_KEY_s0[375]}), .b ({new_AGEMA_signal_1630, CONST_ADDITION[119]}), .c ({new_AGEMA_signal_1658, n499}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U540 ( .a ({new_AGEMA_signal_1216, n500}), .b ({new_AGEMA_signal_1658, n499}), .c ({ROUND_OUT_s1[87], ROUND_OUT_s0[87]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U551 ( .a ({ROUND_KEY_s1[371], ROUND_KEY_s0[371]}), .b ({new_AGEMA_signal_1628, CONST_ADDITION[115]}), .c ({new_AGEMA_signal_1660, n507}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U552 ( .a ({new_AGEMA_signal_1228, n508}), .b ({new_AGEMA_signal_1660, n507}), .c ({ROUND_OUT_s1[83], ROUND_OUT_s0[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U563 ( .a ({ROUND_KEY_s1[367], ROUND_KEY_s0[367]}), .b ({new_AGEMA_signal_1627, CONST_ADDITION[111]}), .c ({new_AGEMA_signal_1662, n515}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U564 ( .a ({new_AGEMA_signal_1240, n516}), .b ({new_AGEMA_signal_1662, n515}), .c ({ROUND_OUT_s1[79], ROUND_OUT_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U575 ( .a ({ROUND_KEY_s1[363], ROUND_KEY_s0[363]}), .b ({new_AGEMA_signal_1625, CONST_ADDITION[107]}), .c ({new_AGEMA_signal_1664, n523}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U576 ( .a ({new_AGEMA_signal_1252, n524}), .b ({new_AGEMA_signal_1664, n523}), .c ({ROUND_OUT_s1[75], ROUND_OUT_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U587 ( .a ({ROUND_KEY_s1[359], ROUND_KEY_s0[359]}), .b ({new_AGEMA_signal_1624, CONST_ADDITION[103]}), .c ({new_AGEMA_signal_1666, n531}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U588 ( .a ({new_AGEMA_signal_1264, n532}), .b ({new_AGEMA_signal_1666, n531}), .c ({ROUND_OUT_s1[71], ROUND_OUT_s0[71]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_0_U5 ( .a ({new_AGEMA_signal_1531, S_0_R1[2]}), .b ({ROUND_IN_s1[1], ROUND_IN_s0[1]}), .c ({new_AGEMA_signal_1586, SHIFTROWS[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_0_U1 ( .a ({new_AGEMA_signal_1530, S_0_R2[1]}), .b ({ROUND_IN_s1[5], ROUND_IN_s0[5]}), .c ({new_AGEMA_signal_1588, SHIFTROWS[15]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_0_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1404, SHIFTROWS[13]}), .b ({new_AGEMA_signal_1406, SHIFTROWS[14]}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_1530, S_0_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_0_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[3], ROUND_IN_s0[3]}), .b ({new_AGEMA_signal_1404, SHIFTROWS[13]}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_1531, S_0_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_1_U5 ( .a ({new_AGEMA_signal_1533, S_1_R1[2]}), .b ({ROUND_IN_s1[9], ROUND_IN_s0[9]}), .c ({new_AGEMA_signal_1589, SHIFTROWS[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_1_U1 ( .a ({new_AGEMA_signal_1532, S_1_R2[1]}), .b ({ROUND_IN_s1[13], ROUND_IN_s0[13]}), .c ({new_AGEMA_signal_1591, SHIFTROWS[23]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_1_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1409, SHIFTROWS[21]}), .b ({new_AGEMA_signal_1411, SHIFTROWS[22]}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_1532, S_1_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_1_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[11], ROUND_IN_s0[11]}), .b ({new_AGEMA_signal_1409, SHIFTROWS[21]}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_1533, S_1_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_2_U5 ( .a ({new_AGEMA_signal_1535, S_2_R1[2]}), .b ({ROUND_IN_s1[17], ROUND_IN_s0[17]}), .c ({new_AGEMA_signal_1592, SHIFTROWS[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_2_U1 ( .a ({new_AGEMA_signal_1534, S_2_R2[1]}), .b ({ROUND_IN_s1[21], ROUND_IN_s0[21]}), .c ({new_AGEMA_signal_1594, SHIFTROWS[31]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_2_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1414, SHIFTROWS[29]}), .b ({new_AGEMA_signal_1416, SHIFTROWS[30]}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_1534, S_2_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_2_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[19], ROUND_IN_s0[19]}), .b ({new_AGEMA_signal_1414, SHIFTROWS[29]}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_1535, S_2_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_3_U5 ( .a ({new_AGEMA_signal_1537, S_3_R1[2]}), .b ({ROUND_IN_s1[25], ROUND_IN_s0[25]}), .c ({new_AGEMA_signal_1595, SHIFTROWS[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_3_U1 ( .a ({new_AGEMA_signal_1536, S_3_R2[1]}), .b ({ROUND_IN_s1[29], ROUND_IN_s0[29]}), .c ({new_AGEMA_signal_1597, SHIFTROWS[7]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_3_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1419, SHIFTROWS[5]}), .b ({new_AGEMA_signal_1421, SHIFTROWS[6]}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_1536, S_3_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_3_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[27], ROUND_IN_s0[27]}), .b ({new_AGEMA_signal_1419, SHIFTROWS[5]}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_1537, S_3_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_4_U5 ( .a ({new_AGEMA_signal_1539, S_4_R1[2]}), .b ({ROUND_IN_s1[33], ROUND_IN_s0[33]}), .c ({new_AGEMA_signal_1598, SHIFTROWS[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_4_U1 ( .a ({new_AGEMA_signal_1538, S_4_R2[1]}), .b ({ROUND_IN_s1[37], ROUND_IN_s0[37]}), .c ({new_AGEMA_signal_1600, SHIFTROWS[55]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_4_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1424, SHIFTROWS[53]}), .b ({new_AGEMA_signal_1426, SHIFTROWS[54]}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_1538, S_4_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_4_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[35], ROUND_IN_s0[35]}), .b ({new_AGEMA_signal_1424, SHIFTROWS[53]}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_1539, S_4_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_5_U5 ( .a ({new_AGEMA_signal_1541, S_5_R1[2]}), .b ({ROUND_IN_s1[41], ROUND_IN_s0[41]}), .c ({new_AGEMA_signal_1601, SHIFTROWS[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_5_U1 ( .a ({new_AGEMA_signal_1540, S_5_R2[1]}), .b ({ROUND_IN_s1[45], ROUND_IN_s0[45]}), .c ({new_AGEMA_signal_1603, SHIFTROWS[63]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_5_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1429, SHIFTROWS[61]}), .b ({new_AGEMA_signal_1431, SHIFTROWS[62]}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_1540, S_5_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_5_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[43], ROUND_IN_s0[43]}), .b ({new_AGEMA_signal_1429, SHIFTROWS[61]}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_1541, S_5_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_6_U5 ( .a ({new_AGEMA_signal_1543, S_6_R1[2]}), .b ({ROUND_IN_s1[49], ROUND_IN_s0[49]}), .c ({new_AGEMA_signal_1604, SHIFTROWS[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_6_U1 ( .a ({new_AGEMA_signal_1542, S_6_R2[1]}), .b ({ROUND_IN_s1[53], ROUND_IN_s0[53]}), .c ({new_AGEMA_signal_1606, SHIFTROWS[39]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_6_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1434, SHIFTROWS[37]}), .b ({new_AGEMA_signal_1436, SHIFTROWS[38]}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_1542, S_6_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_6_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[51], ROUND_IN_s0[51]}), .b ({new_AGEMA_signal_1434, SHIFTROWS[37]}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_1543, S_6_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_7_U5 ( .a ({new_AGEMA_signal_1545, S_7_R1[2]}), .b ({ROUND_IN_s1[57], ROUND_IN_s0[57]}), .c ({new_AGEMA_signal_1607, SHIFTROWS[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_7_U1 ( .a ({new_AGEMA_signal_1544, S_7_R2[1]}), .b ({ROUND_IN_s1[61], ROUND_IN_s0[61]}), .c ({new_AGEMA_signal_1609, SHIFTROWS[47]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_7_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1439, SHIFTROWS[45]}), .b ({new_AGEMA_signal_1441, SHIFTROWS[46]}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_1544, S_7_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_7_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[59], ROUND_IN_s0[59]}), .b ({new_AGEMA_signal_1439, SHIFTROWS[45]}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_1545, S_7_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_8_U5 ( .a ({new_AGEMA_signal_1547, S_8_R1[2]}), .b ({ROUND_IN_s1[65], ROUND_IN_s0[65]}), .c ({new_AGEMA_signal_1610, CONST_ADDITION[67]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_8_U1 ( .a ({new_AGEMA_signal_1546, S_8_R2[1]}), .b ({ROUND_IN_s1[69], ROUND_IN_s0[69]}), .c ({new_AGEMA_signal_1612, CONST_ADDITION[71]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_8_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1444, CONST_ADDITION[69]}), .b ({new_AGEMA_signal_1446, CONST_ADDITION[70]}), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_1546, S_8_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_8_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[67], ROUND_IN_s0[67]}), .b ({new_AGEMA_signal_1444, CONST_ADDITION[69]}), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_1547, S_8_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_9_U5 ( .a ({new_AGEMA_signal_1549, S_9_R1[2]}), .b ({ROUND_IN_s1[73], ROUND_IN_s0[73]}), .c ({new_AGEMA_signal_1613, CONST_ADDITION[75]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_9_U1 ( .a ({new_AGEMA_signal_1548, S_9_R2[1]}), .b ({ROUND_IN_s1[77], ROUND_IN_s0[77]}), .c ({new_AGEMA_signal_1615, CONST_ADDITION[79]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_9_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1449, CONST_ADDITION[77]}), .b ({new_AGEMA_signal_1451, CONST_ADDITION[78]}), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_1548, S_9_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_9_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[75], ROUND_IN_s0[75]}), .b ({new_AGEMA_signal_1449, CONST_ADDITION[77]}), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_1549, S_9_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_10_U5 ( .a ({new_AGEMA_signal_1551, S_10_R1[2]}), .b ({ROUND_IN_s1[81], ROUND_IN_s0[81]}), .c ({new_AGEMA_signal_1616, CONST_ADDITION[83]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_10_U1 ( .a ({new_AGEMA_signal_1550, S_10_R2[1]}), .b ({ROUND_IN_s1[85], ROUND_IN_s0[85]}), .c ({new_AGEMA_signal_1618, CONST_ADDITION[87]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_10_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1454, CONST_ADDITION[85]}), .b ({new_AGEMA_signal_1456, CONST_ADDITION[86]}), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_1550, S_10_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_10_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[83], ROUND_IN_s0[83]}), .b ({new_AGEMA_signal_1454, CONST_ADDITION[85]}), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_1551, S_10_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_11_U5 ( .a ({new_AGEMA_signal_1553, S_11_R1[2]}), .b ({ROUND_IN_s1[89], ROUND_IN_s0[89]}), .c ({new_AGEMA_signal_1619, CONST_ADDITION[91]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_11_U1 ( .a ({new_AGEMA_signal_1552, S_11_R2[1]}), .b ({ROUND_IN_s1[93], ROUND_IN_s0[93]}), .c ({new_AGEMA_signal_1621, CONST_ADDITION[95]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_11_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1459, CONST_ADDITION[93]}), .b ({new_AGEMA_signal_1461, CONST_ADDITION[94]}), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_1552, S_11_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_11_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[91], ROUND_IN_s0[91]}), .b ({new_AGEMA_signal_1459, CONST_ADDITION[93]}), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_1553, S_11_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_12_U5 ( .a ({new_AGEMA_signal_1555, S_12_R1[2]}), .b ({ROUND_IN_s1[97], ROUND_IN_s0[97]}), .c ({new_AGEMA_signal_1622, CONST_ADDITION[99]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_12_U1 ( .a ({new_AGEMA_signal_1554, S_12_R2[1]}), .b ({ROUND_IN_s1[101], ROUND_IN_s0[101]}), .c ({new_AGEMA_signal_1624, CONST_ADDITION[103]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_12_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1464, CONST_ADDITION[101]}), .b ({new_AGEMA_signal_1466, CONST_ADDITION[102]}), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_1554, S_12_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_12_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[99], ROUND_IN_s0[99]}), .b ({new_AGEMA_signal_1464, CONST_ADDITION[101]}), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_1555, S_12_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_13_U5 ( .a ({new_AGEMA_signal_1557, S_13_R1[2]}), .b ({ROUND_IN_s1[105], ROUND_IN_s0[105]}), .c ({new_AGEMA_signal_1625, CONST_ADDITION[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_13_U1 ( .a ({new_AGEMA_signal_1556, S_13_R2[1]}), .b ({ROUND_IN_s1[109], ROUND_IN_s0[109]}), .c ({new_AGEMA_signal_1627, CONST_ADDITION[111]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_13_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1469, CONST_ADDITION[109]}), .b ({new_AGEMA_signal_1471, CONST_ADDITION[110]}), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_1556, S_13_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_13_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[107], ROUND_IN_s0[107]}), .b ({new_AGEMA_signal_1469, CONST_ADDITION[109]}), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_1557, S_13_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_14_U5 ( .a ({new_AGEMA_signal_1559, S_14_R1[2]}), .b ({ROUND_IN_s1[113], ROUND_IN_s0[113]}), .c ({new_AGEMA_signal_1628, CONST_ADDITION[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_14_U1 ( .a ({new_AGEMA_signal_1558, S_14_R2[1]}), .b ({ROUND_IN_s1[117], ROUND_IN_s0[117]}), .c ({new_AGEMA_signal_1630, CONST_ADDITION[119]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_14_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1474, CONST_ADDITION[117]}), .b ({new_AGEMA_signal_1476, CONST_ADDITION[118]}), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_1558, S_14_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_14_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[115], ROUND_IN_s0[115]}), .b ({new_AGEMA_signal_1474, CONST_ADDITION[117]}), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_1559, S_14_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_15_U5 ( .a ({new_AGEMA_signal_1561, S_15_R1[2]}), .b ({ROUND_IN_s1[121], ROUND_IN_s0[121]}), .c ({new_AGEMA_signal_1631, SUBSTITUTION[123]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_15_U1 ( .a ({new_AGEMA_signal_1560, S_15_R2[1]}), .b ({ROUND_IN_s1[125], ROUND_IN_s0[125]}), .c ({new_AGEMA_signal_1633, CONST_ADDITION[127]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_15_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_1479, CONST_ADDITION[125]}), .b ({new_AGEMA_signal_1481, CONST_ADDITION[126]}), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_1560, S_15_R2[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_15_NOR1Inst_2_U1 ( .a ({ROUND_IN_s1[123], ROUND_IN_s0[123]}), .b ({new_AGEMA_signal_1479, CONST_ADDITION[125]}), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_1561, S_15_R1[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U96 ( .a ({new_AGEMA_signal_1594, SHIFTROWS[31]}), .b ({ROUND_OUT_s1[31], ROUND_OUT_s0[31]}), .c ({ROUND_OUT_s1[127], ROUND_OUT_s0[127]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U95 ( .a ({ROUND_OUT_s1[95], ROUND_OUT_s0[95]}), .b ({new_AGEMA_signal_1603, SHIFTROWS[63]}), .c ({ROUND_OUT_s1[31], ROUND_OUT_s0[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U84 ( .a ({new_AGEMA_signal_1588, SHIFTROWS[15]}), .b ({ROUND_OUT_s1[15], ROUND_OUT_s0[15]}), .c ({ROUND_OUT_s1[111], ROUND_OUT_s0[111]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U83 ( .a ({ROUND_OUT_s1[79], ROUND_OUT_s0[79]}), .b ({new_AGEMA_signal_1609, SHIFTROWS[47]}), .c ({ROUND_OUT_s1[15], ROUND_OUT_s0[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U82 ( .a ({new_AGEMA_signal_1591, SHIFTROWS[23]}), .b ({ROUND_OUT_s1[23], ROUND_OUT_s0[23]}), .c ({ROUND_OUT_s1[119], ROUND_OUT_s0[119]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U81 ( .a ({ROUND_OUT_s1[87], ROUND_OUT_s0[87]}), .b ({new_AGEMA_signal_1600, SHIFTROWS[55]}), .c ({ROUND_OUT_s1[23], ROUND_OUT_s0[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U76 ( .a ({new_AGEMA_signal_1592, SHIFTROWS[27]}), .b ({ROUND_OUT_s1[27], ROUND_OUT_s0[27]}), .c ({ROUND_OUT_s1[123], ROUND_OUT_s0[123]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U75 ( .a ({ROUND_OUT_s1[91], ROUND_OUT_s0[91]}), .b ({new_AGEMA_signal_1601, SHIFTROWS[59]}), .c ({ROUND_OUT_s1[27], ROUND_OUT_s0[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U70 ( .a ({new_AGEMA_signal_1586, SHIFTROWS[11]}), .b ({ROUND_OUT_s1[11], ROUND_OUT_s0[11]}), .c ({ROUND_OUT_s1[107], ROUND_OUT_s0[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U69 ( .a ({ROUND_OUT_s1[75], ROUND_OUT_s0[75]}), .b ({new_AGEMA_signal_1607, SHIFTROWS[43]}), .c ({ROUND_OUT_s1[11], ROUND_OUT_s0[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U54 ( .a ({new_AGEMA_signal_1597, SHIFTROWS[7]}), .b ({ROUND_OUT_s1[7], ROUND_OUT_s0[7]}), .c ({ROUND_OUT_s1[103], ROUND_OUT_s0[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U53 ( .a ({ROUND_OUT_s1[71], ROUND_OUT_s0[71]}), .b ({new_AGEMA_signal_1606, SHIFTROWS[39]}), .c ({ROUND_OUT_s1[7], ROUND_OUT_s0[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U52 ( .a ({new_AGEMA_signal_1589, SHIFTROWS[19]}), .b ({ROUND_OUT_s1[19], ROUND_OUT_s0[19]}), .c ({ROUND_OUT_s1[115], ROUND_OUT_s0[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U51 ( .a ({ROUND_OUT_s1[83], ROUND_OUT_s0[83]}), .b ({new_AGEMA_signal_1598, SHIFTROWS[51]}), .c ({ROUND_OUT_s1[19], ROUND_OUT_s0[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U40 ( .a ({new_AGEMA_signal_1595, SHIFTROWS[3]}), .b ({ROUND_OUT_s1[3], ROUND_OUT_s0[3]}), .c ({ROUND_OUT_s1[99], ROUND_OUT_s0[99]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U39 ( .a ({ROUND_OUT_s1[67], ROUND_OUT_s0[67]}), .b ({new_AGEMA_signal_1604, SHIFTROWS[35]}), .c ({ROUND_OUT_s1[3], ROUND_OUT_s0[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U29 ( .a ({new_AGEMA_signal_1604, SHIFTROWS[35]}), .b ({new_AGEMA_signal_1728, SHIFTROWS[67]}), .c ({ROUND_OUT_s1[35], ROUND_OUT_s0[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U25 ( .a ({new_AGEMA_signal_1606, SHIFTROWS[39]}), .b ({new_AGEMA_signal_1727, SHIFTROWS[71]}), .c ({ROUND_OUT_s1[39], ROUND_OUT_s0[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U21 ( .a ({new_AGEMA_signal_1607, SHIFTROWS[43]}), .b ({new_AGEMA_signal_1726, SHIFTROWS[75]}), .c ({ROUND_OUT_s1[43], ROUND_OUT_s0[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U17 ( .a ({new_AGEMA_signal_1609, SHIFTROWS[47]}), .b ({new_AGEMA_signal_1725, SHIFTROWS[79]}), .c ({ROUND_OUT_s1[47], ROUND_OUT_s0[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U13 ( .a ({new_AGEMA_signal_1598, SHIFTROWS[51]}), .b ({new_AGEMA_signal_1724, SHIFTROWS[83]}), .c ({ROUND_OUT_s1[51], ROUND_OUT_s0[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U9 ( .a ({new_AGEMA_signal_1600, SHIFTROWS[55]}), .b ({new_AGEMA_signal_1723, SHIFTROWS[87]}), .c ({ROUND_OUT_s1[55], ROUND_OUT_s0[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U5 ( .a ({new_AGEMA_signal_1601, SHIFTROWS[59]}), .b ({new_AGEMA_signal_1730, SHIFTROWS[91]}), .c ({ROUND_OUT_s1[59], ROUND_OUT_s0[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U1 ( .a ({new_AGEMA_signal_1603, SHIFTROWS[63]}), .b ({new_AGEMA_signal_1729, SHIFTROWS[95]}), .c ({ROUND_OUT_s1[63], ROUND_OUT_s0[63]}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    not_masked #(.security_order(1), .pipeline(0)) U399 ( .a ({new_AGEMA_signal_1752, SUBSTITUTION_57}), .b ({new_AGEMA_signal_1782, SHIFTROWS[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U407 ( .a ({ROUND_KEY_s1[353], ROUND_KEY_s0[353]}), .b ({new_AGEMA_signal_1762, CONST_ADDITION[97]}), .c ({new_AGEMA_signal_1784, n409}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U408 ( .a ({new_AGEMA_signal_1090, n410}), .b ({new_AGEMA_signal_1784, n409}), .c ({ROUND_OUT_s1[65], ROUND_OUT_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U422 ( .a ({ROUND_KEY_s1[348], ROUND_KEY_s0[348]}), .b ({new_AGEMA_signal_1761, CONST_ADDITION[92]}), .c ({new_AGEMA_signal_1786, n419}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U423 ( .a ({new_AGEMA_signal_1105, n420}), .b ({new_AGEMA_signal_1786, n419}), .c ({new_AGEMA_signal_1849, SHIFTROWS[84]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U431 ( .a ({new_AGEMA_signal_1760, SUBSTITUTION_89}), .b ({ROUND_KEY_s1[345], ROUND_KEY_s0[345]}), .c ({new_AGEMA_signal_1788, n425}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U432 ( .a ({new_AGEMA_signal_1114, n426}), .b ({new_AGEMA_signal_1788, n425}), .c ({new_AGEMA_signal_1850, n427}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U433 ( .a ({1'b0, CONST_IN[5]}), .b ({new_AGEMA_signal_1850, n427}), .c ({new_AGEMA_signal_1890, SHIFTROWS[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U448 ( .a ({ROUND_KEY_s1[340], ROUND_KEY_s0[340]}), .b ({new_AGEMA_signal_1759, CONST_ADDITION[84]}), .c ({new_AGEMA_signal_1790, n437}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U449 ( .a ({new_AGEMA_signal_1129, n438}), .b ({new_AGEMA_signal_1790, n437}), .c ({new_AGEMA_signal_1851, SHIFTROWS[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U457 ( .a ({ROUND_KEY_s1[337], ROUND_KEY_s0[337]}), .b ({new_AGEMA_signal_1758, CONST_ADDITION[81]}), .c ({new_AGEMA_signal_1792, n443}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U458 ( .a ({new_AGEMA_signal_1138, n444}), .b ({new_AGEMA_signal_1792, n443}), .c ({new_AGEMA_signal_1852, SHIFTROWS[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U472 ( .a ({ROUND_KEY_s1[332], ROUND_KEY_s0[332]}), .b ({new_AGEMA_signal_1757, CONST_ADDITION[76]}), .c ({new_AGEMA_signal_1794, n453}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U473 ( .a ({new_AGEMA_signal_1153, n454}), .b ({new_AGEMA_signal_1794, n453}), .c ({new_AGEMA_signal_1853, SHIFTROWS[68]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U481 ( .a ({ROUND_KEY_s1[329], ROUND_KEY_s0[329]}), .b ({new_AGEMA_signal_1756, CONST_ADDITION[73]}), .c ({new_AGEMA_signal_1796, n459}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U482 ( .a ({new_AGEMA_signal_1162, n460}), .b ({new_AGEMA_signal_1796, n459}), .c ({new_AGEMA_signal_1854, SHIFTROWS[65]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U496 ( .a ({ROUND_KEY_s1[324], ROUND_KEY_s0[324]}), .b ({new_AGEMA_signal_1755, CONST_ADDITION[68]}), .c ({new_AGEMA_signal_1798, n469}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U497 ( .a ({new_AGEMA_signal_1177, n470}), .b ({new_AGEMA_signal_1798, n469}), .c ({new_AGEMA_signal_1855, SHIFTROWS[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U505 ( .a ({ROUND_KEY_s1[321], ROUND_KEY_s0[321]}), .b ({new_AGEMA_signal_1754, CONST_ADDITION[65]}), .c ({new_AGEMA_signal_1800, n475}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U506 ( .a ({new_AGEMA_signal_1186, n476}), .b ({new_AGEMA_signal_1800, n475}), .c ({new_AGEMA_signal_1856, SHIFTROWS[89]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U520 ( .a ({ROUND_KEY_s1[380], ROUND_KEY_s0[380]}), .b ({new_AGEMA_signal_1769, CONST_ADDITION[124]}), .c ({new_AGEMA_signal_1802, n485}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U521 ( .a ({new_AGEMA_signal_1201, n486}), .b ({new_AGEMA_signal_1802, n485}), .c ({ROUND_OUT_s1[92], ROUND_OUT_s0[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U531 ( .a ({new_AGEMA_signal_1768, SUBSTITUTION[121]}), .b ({ROUND_KEY_s1[377], ROUND_KEY_s0[377]}), .c ({new_AGEMA_signal_1805, n493}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U532 ( .a ({new_AGEMA_signal_1210, n494}), .b ({new_AGEMA_signal_1805, n493}), .c ({new_AGEMA_signal_1858, n495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U533 ( .a ({1'b0, CONST_IN[1]}), .b ({new_AGEMA_signal_1858, n495}), .c ({ROUND_OUT_s1[89], ROUND_OUT_s0[89]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U548 ( .a ({ROUND_KEY_s1[372], ROUND_KEY_s0[372]}), .b ({new_AGEMA_signal_1767, CONST_ADDITION[116]}), .c ({new_AGEMA_signal_1807, n505}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U549 ( .a ({new_AGEMA_signal_1225, n506}), .b ({new_AGEMA_signal_1807, n505}), .c ({ROUND_OUT_s1[84], ROUND_OUT_s0[84]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U557 ( .a ({ROUND_KEY_s1[369], ROUND_KEY_s0[369]}), .b ({new_AGEMA_signal_1766, CONST_ADDITION[113]}), .c ({new_AGEMA_signal_1809, n511}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U558 ( .a ({new_AGEMA_signal_1234, n512}), .b ({new_AGEMA_signal_1809, n511}), .c ({ROUND_OUT_s1[81], ROUND_OUT_s0[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U572 ( .a ({ROUND_KEY_s1[364], ROUND_KEY_s0[364]}), .b ({new_AGEMA_signal_1765, CONST_ADDITION[108]}), .c ({new_AGEMA_signal_1811, n521}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U573 ( .a ({new_AGEMA_signal_1249, n522}), .b ({new_AGEMA_signal_1811, n521}), .c ({ROUND_OUT_s1[76], ROUND_OUT_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U581 ( .a ({ROUND_KEY_s1[361], ROUND_KEY_s0[361]}), .b ({new_AGEMA_signal_1764, CONST_ADDITION[105]}), .c ({new_AGEMA_signal_1813, n527}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U582 ( .a ({new_AGEMA_signal_1258, n528}), .b ({new_AGEMA_signal_1813, n527}), .c ({ROUND_OUT_s1[73], ROUND_OUT_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U596 ( .a ({ROUND_KEY_s1[356], ROUND_KEY_s0[356]}), .b ({new_AGEMA_signal_1763, CONST_ADDITION[100]}), .c ({new_AGEMA_signal_1815, n537}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U597 ( .a ({new_AGEMA_signal_1273, n538}), .b ({new_AGEMA_signal_1815, n537}), .c ({ROUND_OUT_s1[68], ROUND_OUT_s0[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_0_U7 ( .a ({new_AGEMA_signal_1667, S_0_R2[2]}), .b ({ROUND_IN_s1[7], ROUND_IN_s0[7]}), .c ({new_AGEMA_signal_1738, SHIFTROWS[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_0_U4 ( .a ({new_AGEMA_signal_1668, S_0_R1[3]}), .b ({ROUND_IN_s1[3], ROUND_IN_s0[3]}), .c ({new_AGEMA_signal_1739, SHIFTROWS[12]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_0_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1588, SHIFTROWS[15]}), .b ({new_AGEMA_signal_1402, SHIFTROWS[10]}), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_1667, S_0_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_0_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1406, SHIFTROWS[14]}), .b ({new_AGEMA_signal_1588, SHIFTROWS[15]}), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_1668, S_0_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_1_U7 ( .a ({new_AGEMA_signal_1669, S_1_R2[2]}), .b ({ROUND_IN_s1[15], ROUND_IN_s0[15]}), .c ({new_AGEMA_signal_1740, SHIFTROWS[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_1_U4 ( .a ({new_AGEMA_signal_1670, S_1_R1[3]}), .b ({ROUND_IN_s1[11], ROUND_IN_s0[11]}), .c ({new_AGEMA_signal_1741, SHIFTROWS[20]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_1_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1591, SHIFTROWS[23]}), .b ({new_AGEMA_signal_1407, SHIFTROWS[18]}), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_1669, S_1_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_1_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1411, SHIFTROWS[22]}), .b ({new_AGEMA_signal_1591, SHIFTROWS[23]}), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_1670, S_1_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_2_U7 ( .a ({new_AGEMA_signal_1671, S_2_R2[2]}), .b ({ROUND_IN_s1[23], ROUND_IN_s0[23]}), .c ({new_AGEMA_signal_1742, SHIFTROWS[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_2_U4 ( .a ({new_AGEMA_signal_1672, S_2_R1[3]}), .b ({ROUND_IN_s1[19], ROUND_IN_s0[19]}), .c ({new_AGEMA_signal_1743, SHIFTROWS[28]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_2_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1594, SHIFTROWS[31]}), .b ({new_AGEMA_signal_1412, SHIFTROWS[26]}), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_1671, S_2_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_2_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1416, SHIFTROWS[30]}), .b ({new_AGEMA_signal_1594, SHIFTROWS[31]}), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_1672, S_2_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_3_U7 ( .a ({new_AGEMA_signal_1673, S_3_R2[2]}), .b ({ROUND_IN_s1[31], ROUND_IN_s0[31]}), .c ({new_AGEMA_signal_1744, SHIFTROWS[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_3_U4 ( .a ({new_AGEMA_signal_1674, S_3_R1[3]}), .b ({ROUND_IN_s1[27], ROUND_IN_s0[27]}), .c ({new_AGEMA_signal_1745, SHIFTROWS[4]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_3_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1597, SHIFTROWS[7]}), .b ({new_AGEMA_signal_1417, SHIFTROWS[2]}), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_1673, S_3_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_3_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1421, SHIFTROWS[6]}), .b ({new_AGEMA_signal_1597, SHIFTROWS[7]}), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_1674, S_3_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_4_U7 ( .a ({new_AGEMA_signal_1675, S_4_R2[2]}), .b ({ROUND_IN_s1[39], ROUND_IN_s0[39]}), .c ({new_AGEMA_signal_1746, SHIFTROWS[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_4_U4 ( .a ({new_AGEMA_signal_1676, S_4_R1[3]}), .b ({ROUND_IN_s1[35], ROUND_IN_s0[35]}), .c ({new_AGEMA_signal_1747, SHIFTROWS[52]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_4_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1600, SHIFTROWS[55]}), .b ({new_AGEMA_signal_1422, SHIFTROWS[50]}), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_1675, S_4_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_4_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1426, SHIFTROWS[54]}), .b ({new_AGEMA_signal_1600, SHIFTROWS[55]}), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_1676, S_4_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_5_U7 ( .a ({new_AGEMA_signal_1677, S_5_R2[2]}), .b ({ROUND_IN_s1[47], ROUND_IN_s0[47]}), .c ({new_AGEMA_signal_1748, SHIFTROWS[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_5_U4 ( .a ({new_AGEMA_signal_1678, S_5_R1[3]}), .b ({ROUND_IN_s1[43], ROUND_IN_s0[43]}), .c ({new_AGEMA_signal_1749, SHIFTROWS[60]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_5_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1603, SHIFTROWS[63]}), .b ({new_AGEMA_signal_1427, SHIFTROWS[58]}), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_1677, S_5_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_5_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1431, SHIFTROWS[62]}), .b ({new_AGEMA_signal_1603, SHIFTROWS[63]}), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_1678, S_5_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_6_U7 ( .a ({new_AGEMA_signal_1679, S_6_R2[2]}), .b ({ROUND_IN_s1[55], ROUND_IN_s0[55]}), .c ({new_AGEMA_signal_1750, SHIFTROWS[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_6_U4 ( .a ({new_AGEMA_signal_1680, S_6_R1[3]}), .b ({ROUND_IN_s1[51], ROUND_IN_s0[51]}), .c ({new_AGEMA_signal_1751, SHIFTROWS[36]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_6_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1606, SHIFTROWS[39]}), .b ({new_AGEMA_signal_1432, SHIFTROWS[34]}), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_1679, S_6_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_6_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1436, SHIFTROWS[38]}), .b ({new_AGEMA_signal_1606, SHIFTROWS[39]}), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_1680, S_6_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_7_U7 ( .a ({new_AGEMA_signal_1681, S_7_R2[2]}), .b ({ROUND_IN_s1[63], ROUND_IN_s0[63]}), .c ({new_AGEMA_signal_1752, SUBSTITUTION_57}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_7_U4 ( .a ({new_AGEMA_signal_1682, S_7_R1[3]}), .b ({ROUND_IN_s1[59], ROUND_IN_s0[59]}), .c ({new_AGEMA_signal_1753, SHIFTROWS[44]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_7_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1609, SHIFTROWS[47]}), .b ({new_AGEMA_signal_1437, SHIFTROWS[42]}), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_1681, S_7_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_7_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1441, SHIFTROWS[46]}), .b ({new_AGEMA_signal_1609, SHIFTROWS[47]}), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_1682, S_7_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_8_U7 ( .a ({new_AGEMA_signal_1683, S_8_R2[2]}), .b ({ROUND_IN_s1[71], ROUND_IN_s0[71]}), .c ({new_AGEMA_signal_1754, CONST_ADDITION[65]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_8_U4 ( .a ({new_AGEMA_signal_1684, S_8_R1[3]}), .b ({ROUND_IN_s1[67], ROUND_IN_s0[67]}), .c ({new_AGEMA_signal_1755, CONST_ADDITION[68]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_8_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1612, CONST_ADDITION[71]}), .b ({new_AGEMA_signal_1442, CONST_ADDITION[66]}), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_1683, S_8_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_8_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1446, CONST_ADDITION[70]}), .b ({new_AGEMA_signal_1612, CONST_ADDITION[71]}), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_1684, S_8_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_9_U7 ( .a ({new_AGEMA_signal_1685, S_9_R2[2]}), .b ({ROUND_IN_s1[79], ROUND_IN_s0[79]}), .c ({new_AGEMA_signal_1756, CONST_ADDITION[73]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_9_U4 ( .a ({new_AGEMA_signal_1686, S_9_R1[3]}), .b ({ROUND_IN_s1[75], ROUND_IN_s0[75]}), .c ({new_AGEMA_signal_1757, CONST_ADDITION[76]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_9_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1615, CONST_ADDITION[79]}), .b ({new_AGEMA_signal_1447, CONST_ADDITION[74]}), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_1685, S_9_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_9_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1451, CONST_ADDITION[78]}), .b ({new_AGEMA_signal_1615, CONST_ADDITION[79]}), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_1686, S_9_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_10_U7 ( .a ({new_AGEMA_signal_1687, S_10_R2[2]}), .b ({ROUND_IN_s1[87], ROUND_IN_s0[87]}), .c ({new_AGEMA_signal_1758, CONST_ADDITION[81]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_10_U4 ( .a ({new_AGEMA_signal_1688, S_10_R1[3]}), .b ({ROUND_IN_s1[83], ROUND_IN_s0[83]}), .c ({new_AGEMA_signal_1759, CONST_ADDITION[84]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_10_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1618, CONST_ADDITION[87]}), .b ({new_AGEMA_signal_1452, CONST_ADDITION[82]}), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_1687, S_10_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_10_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1456, CONST_ADDITION[86]}), .b ({new_AGEMA_signal_1618, CONST_ADDITION[87]}), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_1688, S_10_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_11_U7 ( .a ({new_AGEMA_signal_1689, S_11_R2[2]}), .b ({ROUND_IN_s1[95], ROUND_IN_s0[95]}), .c ({new_AGEMA_signal_1760, SUBSTITUTION_89}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_11_U4 ( .a ({new_AGEMA_signal_1690, S_11_R1[3]}), .b ({ROUND_IN_s1[91], ROUND_IN_s0[91]}), .c ({new_AGEMA_signal_1761, CONST_ADDITION[92]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_11_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1621, CONST_ADDITION[95]}), .b ({new_AGEMA_signal_1457, CONST_ADDITION[90]}), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_1689, S_11_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_11_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1461, CONST_ADDITION[94]}), .b ({new_AGEMA_signal_1621, CONST_ADDITION[95]}), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_1690, S_11_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_12_U7 ( .a ({new_AGEMA_signal_1691, S_12_R2[2]}), .b ({ROUND_IN_s1[103], ROUND_IN_s0[103]}), .c ({new_AGEMA_signal_1762, CONST_ADDITION[97]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_12_U4 ( .a ({new_AGEMA_signal_1692, S_12_R1[3]}), .b ({ROUND_IN_s1[99], ROUND_IN_s0[99]}), .c ({new_AGEMA_signal_1763, CONST_ADDITION[100]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_12_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1624, CONST_ADDITION[103]}), .b ({new_AGEMA_signal_1462, CONST_ADDITION[98]}), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_1691, S_12_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_12_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1466, CONST_ADDITION[102]}), .b ({new_AGEMA_signal_1624, CONST_ADDITION[103]}), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_1692, S_12_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_13_U7 ( .a ({new_AGEMA_signal_1693, S_13_R2[2]}), .b ({ROUND_IN_s1[111], ROUND_IN_s0[111]}), .c ({new_AGEMA_signal_1764, CONST_ADDITION[105]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_13_U4 ( .a ({new_AGEMA_signal_1694, S_13_R1[3]}), .b ({ROUND_IN_s1[107], ROUND_IN_s0[107]}), .c ({new_AGEMA_signal_1765, CONST_ADDITION[108]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_13_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1627, CONST_ADDITION[111]}), .b ({new_AGEMA_signal_1467, CONST_ADDITION[106]}), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_1693, S_13_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_13_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1471, CONST_ADDITION[110]}), .b ({new_AGEMA_signal_1627, CONST_ADDITION[111]}), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_1694, S_13_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_14_U7 ( .a ({new_AGEMA_signal_1695, S_14_R2[2]}), .b ({ROUND_IN_s1[119], ROUND_IN_s0[119]}), .c ({new_AGEMA_signal_1766, CONST_ADDITION[113]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_14_U4 ( .a ({new_AGEMA_signal_1696, S_14_R1[3]}), .b ({ROUND_IN_s1[115], ROUND_IN_s0[115]}), .c ({new_AGEMA_signal_1767, CONST_ADDITION[116]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_14_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1630, CONST_ADDITION[119]}), .b ({new_AGEMA_signal_1472, CONST_ADDITION[114]}), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_1695, S_14_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_14_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1476, CONST_ADDITION[118]}), .b ({new_AGEMA_signal_1630, CONST_ADDITION[119]}), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_1696, S_14_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_15_U7 ( .a ({new_AGEMA_signal_1697, S_15_R2[2]}), .b ({ROUND_IN_s1[127], ROUND_IN_s0[127]}), .c ({new_AGEMA_signal_1768, SUBSTITUTION[121]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_15_U4 ( .a ({new_AGEMA_signal_1698, S_15_R1[3]}), .b ({ROUND_IN_s1[123], ROUND_IN_s0[123]}), .c ({new_AGEMA_signal_1769, CONST_ADDITION[124]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_15_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_1633, CONST_ADDITION[127]}), .b ({new_AGEMA_signal_1477, SUBSTITUTION[122]}), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_1697, S_15_R2[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_15_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_1481, CONST_ADDITION[126]}), .b ({new_AGEMA_signal_1633, CONST_ADDITION[127]}), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_1698, S_15_R1[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U90 ( .a ({new_AGEMA_signal_1743, SHIFTROWS[28]}), .b ({ROUND_OUT_s1[28], ROUND_OUT_s0[28]}), .c ({ROUND_OUT_s1[124], ROUND_OUT_s0[124]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U89 ( .a ({ROUND_OUT_s1[92], ROUND_OUT_s0[92]}), .b ({new_AGEMA_signal_1749, SHIFTROWS[60]}), .c ({ROUND_OUT_s1[28], ROUND_OUT_s0[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U72 ( .a ({new_AGEMA_signal_1739, SHIFTROWS[12]}), .b ({ROUND_OUT_s1[12], ROUND_OUT_s0[12]}), .c ({ROUND_OUT_s1[108], ROUND_OUT_s0[108]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U71 ( .a ({ROUND_OUT_s1[76], ROUND_OUT_s0[76]}), .b ({new_AGEMA_signal_1753, SHIFTROWS[44]}), .c ({ROUND_OUT_s1[12], ROUND_OUT_s0[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U64 ( .a ({new_AGEMA_signal_1738, SHIFTROWS[9]}), .b ({ROUND_OUT_s1[9], ROUND_OUT_s0[9]}), .c ({ROUND_OUT_s1[105], ROUND_OUT_s0[105]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U63 ( .a ({ROUND_OUT_s1[73], ROUND_OUT_s0[73]}), .b ({new_AGEMA_signal_1782, SHIFTROWS[41]}), .c ({ROUND_OUT_s1[9], ROUND_OUT_s0[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U58 ( .a ({new_AGEMA_signal_1741, SHIFTROWS[20]}), .b ({ROUND_OUT_s1[20], ROUND_OUT_s0[20]}), .c ({ROUND_OUT_s1[116], ROUND_OUT_s0[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U57 ( .a ({ROUND_OUT_s1[84], ROUND_OUT_s0[84]}), .b ({new_AGEMA_signal_1747, SHIFTROWS[52]}), .c ({ROUND_OUT_s1[20], ROUND_OUT_s0[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U46 ( .a ({new_AGEMA_signal_1742, SHIFTROWS[25]}), .b ({ROUND_OUT_s1[25], ROUND_OUT_s0[25]}), .c ({ROUND_OUT_s1[121], ROUND_OUT_s0[121]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U45 ( .a ({ROUND_OUT_s1[89], ROUND_OUT_s0[89]}), .b ({new_AGEMA_signal_1748, SHIFTROWS[57]}), .c ({ROUND_OUT_s1[25], ROUND_OUT_s0[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U42 ( .a ({new_AGEMA_signal_1745, SHIFTROWS[4]}), .b ({ROUND_OUT_s1[4], ROUND_OUT_s0[4]}), .c ({ROUND_OUT_s1[100], ROUND_OUT_s0[100]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U41 ( .a ({ROUND_OUT_s1[68], ROUND_OUT_s0[68]}), .b ({new_AGEMA_signal_1751, SHIFTROWS[36]}), .c ({ROUND_OUT_s1[4], ROUND_OUT_s0[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U38 ( .a ({new_AGEMA_signal_1740, SHIFTROWS[17]}), .b ({ROUND_OUT_s1[17], ROUND_OUT_s0[17]}), .c ({ROUND_OUT_s1[113], ROUND_OUT_s0[113]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U37 ( .a ({ROUND_OUT_s1[81], ROUND_OUT_s0[81]}), .b ({new_AGEMA_signal_1746, SHIFTROWS[49]}), .c ({ROUND_OUT_s1[17], ROUND_OUT_s0[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U34 ( .a ({new_AGEMA_signal_1744, SHIFTROWS[1]}), .b ({ROUND_OUT_s1[1], ROUND_OUT_s0[1]}), .c ({ROUND_OUT_s1[97], ROUND_OUT_s0[97]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U33 ( .a ({ROUND_OUT_s1[65], ROUND_OUT_s0[65]}), .b ({new_AGEMA_signal_1750, SHIFTROWS[33]}), .c ({ROUND_OUT_s1[1], ROUND_OUT_s0[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U31 ( .a ({new_AGEMA_signal_1750, SHIFTROWS[33]}), .b ({new_AGEMA_signal_1854, SHIFTROWS[65]}), .c ({ROUND_OUT_s1[33], ROUND_OUT_s0[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U28 ( .a ({new_AGEMA_signal_1751, SHIFTROWS[36]}), .b ({new_AGEMA_signal_1853, SHIFTROWS[68]}), .c ({ROUND_OUT_s1[36], ROUND_OUT_s0[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U23 ( .a ({new_AGEMA_signal_1782, SHIFTROWS[41]}), .b ({new_AGEMA_signal_1852, SHIFTROWS[73]}), .c ({ROUND_OUT_s1[41], ROUND_OUT_s0[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U20 ( .a ({new_AGEMA_signal_1753, SHIFTROWS[44]}), .b ({new_AGEMA_signal_1851, SHIFTROWS[76]}), .c ({ROUND_OUT_s1[44], ROUND_OUT_s0[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U15 ( .a ({new_AGEMA_signal_1746, SHIFTROWS[49]}), .b ({new_AGEMA_signal_1890, SHIFTROWS[81]}), .c ({ROUND_OUT_s1[49], ROUND_OUT_s0[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U12 ( .a ({new_AGEMA_signal_1747, SHIFTROWS[52]}), .b ({new_AGEMA_signal_1849, SHIFTROWS[84]}), .c ({ROUND_OUT_s1[52], ROUND_OUT_s0[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U7 ( .a ({new_AGEMA_signal_1748, SHIFTROWS[57]}), .b ({new_AGEMA_signal_1856, SHIFTROWS[89]}), .c ({ROUND_OUT_s1[57], ROUND_OUT_s0[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U4 ( .a ({new_AGEMA_signal_1749, SHIFTROWS[60]}), .b ({new_AGEMA_signal_1855, SHIFTROWS[92]}), .c ({ROUND_OUT_s1[60], ROUND_OUT_s0[60]}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U410 ( .a ({ROUND_KEY_s1[352], ROUND_KEY_s0[352]}), .b ({new_AGEMA_signal_1876, CONST_ADDITION[96]}), .c ({new_AGEMA_signal_1889, n411}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U411 ( .a ({new_AGEMA_signal_1093, n412}), .b ({new_AGEMA_signal_1889, n411}), .c ({ROUND_OUT_s1[64], ROUND_OUT_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U435 ( .a ({new_AGEMA_signal_1875, SUBSTITUTION_88}), .b ({ROUND_KEY_s1[344], ROUND_KEY_s0[344]}), .c ({new_AGEMA_signal_1892, n428}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U436 ( .a ({new_AGEMA_signal_1117, n429}), .b ({new_AGEMA_signal_1892, n428}), .c ({new_AGEMA_signal_1922, n430}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U437 ( .a ({1'b0, CONST_IN[4]}), .b ({new_AGEMA_signal_1922, n430}), .c ({new_AGEMA_signal_1938, SHIFTROWS[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U460 ( .a ({ROUND_KEY_s1[336], ROUND_KEY_s0[336]}), .b ({new_AGEMA_signal_1874, CONST_ADDITION[80]}), .c ({new_AGEMA_signal_1894, n445}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U461 ( .a ({new_AGEMA_signal_1141, n446}), .b ({new_AGEMA_signal_1894, n445}), .c ({new_AGEMA_signal_1923, SHIFTROWS[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U484 ( .a ({ROUND_KEY_s1[328], ROUND_KEY_s0[328]}), .b ({new_AGEMA_signal_1873, CONST_ADDITION[72]}), .c ({new_AGEMA_signal_1896, n461}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U485 ( .a ({new_AGEMA_signal_1165, n462}), .b ({new_AGEMA_signal_1896, n461}), .c ({new_AGEMA_signal_1924, SHIFTROWS[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U508 ( .a ({ROUND_KEY_s1[320], ROUND_KEY_s0[320]}), .b ({new_AGEMA_signal_1872, CONST_ADDITION[64]}), .c ({new_AGEMA_signal_1898, n477}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U509 ( .a ({new_AGEMA_signal_1189, n478}), .b ({new_AGEMA_signal_1898, n477}), .c ({new_AGEMA_signal_1925, SHIFTROWS[88]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U535 ( .a ({new_AGEMA_signal_1879, SUBSTITUTION[120]}), .b ({ROUND_KEY_s1[376], ROUND_KEY_s0[376]}), .c ({new_AGEMA_signal_1901, n496}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U536 ( .a ({new_AGEMA_signal_1213, n497}), .b ({new_AGEMA_signal_1901, n496}), .c ({new_AGEMA_signal_1926, n498}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) U537 ( .a ({1'b0, CONST_IN[0]}), .b ({new_AGEMA_signal_1926, n498}), .c ({ROUND_OUT_s1[88], ROUND_OUT_s0[88]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U560 ( .a ({ROUND_KEY_s1[368], ROUND_KEY_s0[368]}), .b ({new_AGEMA_signal_1878, CONST_ADDITION[112]}), .c ({new_AGEMA_signal_1903, n513}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U561 ( .a ({new_AGEMA_signal_1237, n514}), .b ({new_AGEMA_signal_1903, n513}), .c ({ROUND_OUT_s1[80], ROUND_OUT_s0[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U584 ( .a ({ROUND_KEY_s1[360], ROUND_KEY_s0[360]}), .b ({new_AGEMA_signal_1877, CONST_ADDITION[104]}), .c ({new_AGEMA_signal_1905, n529}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) U585 ( .a ({new_AGEMA_signal_1261, n530}), .b ({new_AGEMA_signal_1905, n529}), .c ({ROUND_OUT_s1[72], ROUND_OUT_s0[72]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_0_U8 ( .a ({new_AGEMA_signal_1816, S_0_R2[3]}), .b ({ROUND_IN_s1[2], ROUND_IN_s0[2]}), .c ({new_AGEMA_signal_1864, SHIFTROWS[8]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_0_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1738, SHIFTROWS[9]}), .b ({new_AGEMA_signal_1586, SHIFTROWS[11]}), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_1816, S_0_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_1_U8 ( .a ({new_AGEMA_signal_1817, S_1_R2[3]}), .b ({ROUND_IN_s1[10], ROUND_IN_s0[10]}), .c ({new_AGEMA_signal_1865, SHIFTROWS[16]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_1_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1740, SHIFTROWS[17]}), .b ({new_AGEMA_signal_1589, SHIFTROWS[19]}), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_1817, S_1_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_2_U8 ( .a ({new_AGEMA_signal_1818, S_2_R2[3]}), .b ({ROUND_IN_s1[18], ROUND_IN_s0[18]}), .c ({new_AGEMA_signal_1866, SHIFTROWS[24]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_2_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1742, SHIFTROWS[25]}), .b ({new_AGEMA_signal_1592, SHIFTROWS[27]}), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_1818, S_2_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_3_U8 ( .a ({new_AGEMA_signal_1819, S_3_R2[3]}), .b ({ROUND_IN_s1[26], ROUND_IN_s0[26]}), .c ({new_AGEMA_signal_1867, SHIFTROWS[0]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_3_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1744, SHIFTROWS[1]}), .b ({new_AGEMA_signal_1595, SHIFTROWS[3]}), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_1819, S_3_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_4_U8 ( .a ({new_AGEMA_signal_1820, S_4_R2[3]}), .b ({ROUND_IN_s1[34], ROUND_IN_s0[34]}), .c ({new_AGEMA_signal_1868, SHIFTROWS[48]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_4_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1746, SHIFTROWS[49]}), .b ({new_AGEMA_signal_1598, SHIFTROWS[51]}), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_1820, S_4_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_5_U8 ( .a ({new_AGEMA_signal_1821, S_5_R2[3]}), .b ({ROUND_IN_s1[42], ROUND_IN_s0[42]}), .c ({new_AGEMA_signal_1869, SHIFTROWS[56]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_5_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1748, SHIFTROWS[57]}), .b ({new_AGEMA_signal_1601, SHIFTROWS[59]}), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_1821, S_5_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_6_U8 ( .a ({new_AGEMA_signal_1822, S_6_R2[3]}), .b ({ROUND_IN_s1[50], ROUND_IN_s0[50]}), .c ({new_AGEMA_signal_1870, SHIFTROWS[32]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_6_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1750, SHIFTROWS[33]}), .b ({new_AGEMA_signal_1604, SHIFTROWS[35]}), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_1822, S_6_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_7_U8 ( .a ({new_AGEMA_signal_1823, S_7_R2[3]}), .b ({ROUND_IN_s1[58], ROUND_IN_s0[58]}), .c ({new_AGEMA_signal_1871, SHIFTROWS[40]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_7_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1752, SUBSTITUTION_57}), .b ({new_AGEMA_signal_1607, SHIFTROWS[43]}), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_1823, S_7_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_8_U8 ( .a ({new_AGEMA_signal_1824, S_8_R2[3]}), .b ({ROUND_IN_s1[66], ROUND_IN_s0[66]}), .c ({new_AGEMA_signal_1872, CONST_ADDITION[64]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_8_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1754, CONST_ADDITION[65]}), .b ({new_AGEMA_signal_1610, CONST_ADDITION[67]}), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_1824, S_8_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_9_U8 ( .a ({new_AGEMA_signal_1825, S_9_R2[3]}), .b ({ROUND_IN_s1[74], ROUND_IN_s0[74]}), .c ({new_AGEMA_signal_1873, CONST_ADDITION[72]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_9_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1756, CONST_ADDITION[73]}), .b ({new_AGEMA_signal_1613, CONST_ADDITION[75]}), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_1825, S_9_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_10_U8 ( .a ({new_AGEMA_signal_1826, S_10_R2[3]}), .b ({ROUND_IN_s1[82], ROUND_IN_s0[82]}), .c ({new_AGEMA_signal_1874, CONST_ADDITION[80]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_10_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1758, CONST_ADDITION[81]}), .b ({new_AGEMA_signal_1616, CONST_ADDITION[83]}), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_1826, S_10_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_11_U8 ( .a ({new_AGEMA_signal_1827, S_11_R2[3]}), .b ({ROUND_IN_s1[90], ROUND_IN_s0[90]}), .c ({new_AGEMA_signal_1875, SUBSTITUTION_88}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_11_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1760, SUBSTITUTION_89}), .b ({new_AGEMA_signal_1619, CONST_ADDITION[91]}), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_1827, S_11_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_12_U8 ( .a ({new_AGEMA_signal_1828, S_12_R2[3]}), .b ({ROUND_IN_s1[98], ROUND_IN_s0[98]}), .c ({new_AGEMA_signal_1876, CONST_ADDITION[96]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_12_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1762, CONST_ADDITION[97]}), .b ({new_AGEMA_signal_1622, CONST_ADDITION[99]}), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_1828, S_12_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_13_U8 ( .a ({new_AGEMA_signal_1829, S_13_R2[3]}), .b ({ROUND_IN_s1[106], ROUND_IN_s0[106]}), .c ({new_AGEMA_signal_1877, CONST_ADDITION[104]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_13_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1764, CONST_ADDITION[105]}), .b ({new_AGEMA_signal_1625, CONST_ADDITION[107]}), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_1829, S_13_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_14_U8 ( .a ({new_AGEMA_signal_1830, S_14_R2[3]}), .b ({ROUND_IN_s1[114], ROUND_IN_s0[114]}), .c ({new_AGEMA_signal_1878, CONST_ADDITION[112]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_14_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1766, CONST_ADDITION[113]}), .b ({new_AGEMA_signal_1628, CONST_ADDITION[115]}), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_1830, S_14_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) S_15_U8 ( .a ({new_AGEMA_signal_1831, S_15_R2[3]}), .b ({ROUND_IN_s1[122], ROUND_IN_s0[122]}), .c ({new_AGEMA_signal_1879, SUBSTITUTION[120]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(0)) S_15_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_1768, SUBSTITUTION[121]}), .b ({new_AGEMA_signal_1631, SUBSTITUTION[123]}), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_1831, S_15_R2[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U94 ( .a ({new_AGEMA_signal_1867, SHIFTROWS[0]}), .b ({ROUND_OUT_s1[0], ROUND_OUT_s0[0]}), .c ({ROUND_OUT_s1[96], ROUND_OUT_s0[96]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U93 ( .a ({ROUND_OUT_s1[64], ROUND_OUT_s0[64]}), .b ({new_AGEMA_signal_1870, SHIFTROWS[32]}), .c ({ROUND_OUT_s1[0], ROUND_OUT_s0[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U88 ( .a ({new_AGEMA_signal_1866, SHIFTROWS[24]}), .b ({ROUND_OUT_s1[24], ROUND_OUT_s0[24]}), .c ({ROUND_OUT_s1[120], ROUND_OUT_s0[120]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U87 ( .a ({ROUND_OUT_s1[88], ROUND_OUT_s0[88]}), .b ({new_AGEMA_signal_1869, SHIFTROWS[56]}), .c ({ROUND_OUT_s1[24], ROUND_OUT_s0[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U86 ( .a ({new_AGEMA_signal_1865, SHIFTROWS[16]}), .b ({ROUND_OUT_s1[16], ROUND_OUT_s0[16]}), .c ({ROUND_OUT_s1[112], ROUND_OUT_s0[112]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U85 ( .a ({ROUND_OUT_s1[80], ROUND_OUT_s0[80]}), .b ({new_AGEMA_signal_1868, SHIFTROWS[48]}), .c ({ROUND_OUT_s1[16], ROUND_OUT_s0[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U56 ( .a ({new_AGEMA_signal_1864, SHIFTROWS[8]}), .b ({ROUND_OUT_s1[8], ROUND_OUT_s0[8]}), .c ({ROUND_OUT_s1[104], ROUND_OUT_s0[104]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U55 ( .a ({ROUND_OUT_s1[72], ROUND_OUT_s0[72]}), .b ({new_AGEMA_signal_1871, SHIFTROWS[40]}), .c ({ROUND_OUT_s1[8], ROUND_OUT_s0[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U32 ( .a ({new_AGEMA_signal_1870, SHIFTROWS[32]}), .b ({new_AGEMA_signal_1924, SHIFTROWS[64]}), .c ({ROUND_OUT_s1[32], ROUND_OUT_s0[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U24 ( .a ({new_AGEMA_signal_1871, SHIFTROWS[40]}), .b ({new_AGEMA_signal_1923, SHIFTROWS[72]}), .c ({ROUND_OUT_s1[40], ROUND_OUT_s0[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U16 ( .a ({new_AGEMA_signal_1868, SHIFTROWS[48]}), .b ({new_AGEMA_signal_1938, SHIFTROWS[80]}), .c ({ROUND_OUT_s1[48], ROUND_OUT_s0[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) MC_U8 ( .a ({new_AGEMA_signal_1869, SHIFTROWS[56]}), .b ({new_AGEMA_signal_1925, SHIFTROWS[88]}), .c ({ROUND_OUT_s1[56], ROUND_OUT_s0[56]}) ) ;

endmodule
