/* modified netlist. Source: module RoundFunction in file ./test/RoundFunction.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module RoundFunction_HPC2_ClockGating_d3 (ROUND_KEY_s0, /*ROUND_KEY,*/ ROUND_IN_s0, CONST_IN, clk, ROUND_KEY_s1, ROUND_KEY_s2, ROUND_KEY_s3, ROUND_IN_s1, ROUND_IN_s2, ROUND_IN_s3, Fresh, /*rst,*/ ROUND_OUT_s0, ROUND_OUT_s1, ROUND_OUT_s2, ROUND_OUT_s3/*, Synch*/);
    input [383:0] ROUND_KEY_s0 ;
    //input [319:0] ROUND_KEY ;
    input [127:0] ROUND_IN_s0 ;
    input [5:0] CONST_IN ;
    input clk ;
    input [383:0] ROUND_KEY_s1 ;
    input [383:0] ROUND_KEY_s2 ;
    input [383:0] ROUND_KEY_s3 ;
    input [127:0] ROUND_IN_s1 ;
    input [127:0] ROUND_IN_s2 ;
    input [127:0] ROUND_IN_s3 ;
    //input rst ;
    input [767:0] Fresh ;
    output [127:0] ROUND_OUT_s0 ;
    output [127:0] ROUND_OUT_s1 ;
    output [127:0] ROUND_OUT_s2 ;
    output [127:0] ROUND_OUT_s3 ;
    //output Synch ;
    wire SUBSTITUTION_89 ;
    wire SUBSTITUTION_88 ;
    wire SUBSTITUTION_57 ;
    wire n405 ;
    wire n406 ;
    wire n407 ;
    wire n408 ;
    wire n409 ;
    wire n410 ;
    wire n411 ;
    wire n412 ;
    wire n413 ;
    wire n414 ;
    wire n415 ;
    wire n416 ;
    wire n417 ;
    wire n418 ;
    wire n419 ;
    wire n420 ;
    wire n421 ;
    wire n422 ;
    wire n423 ;
    wire n424 ;
    wire n425 ;
    wire n426 ;
    wire n427 ;
    wire n428 ;
    wire n429 ;
    wire n430 ;
    wire n431 ;
    wire n432 ;
    wire n433 ;
    wire n434 ;
    wire n435 ;
    wire n436 ;
    wire n437 ;
    wire n438 ;
    wire n439 ;
    wire n440 ;
    wire n441 ;
    wire n442 ;
    wire n443 ;
    wire n444 ;
    wire n445 ;
    wire n446 ;
    wire n447 ;
    wire n448 ;
    wire n449 ;
    wire n450 ;
    wire n451 ;
    wire n452 ;
    wire n453 ;
    wire n454 ;
    wire n455 ;
    wire n456 ;
    wire n457 ;
    wire n458 ;
    wire n459 ;
    wire n460 ;
    wire n461 ;
    wire n462 ;
    wire n463 ;
    wire n464 ;
    wire n465 ;
    wire n466 ;
    wire n467 ;
    wire n468 ;
    wire n469 ;
    wire n470 ;
    wire n471 ;
    wire n472 ;
    wire n473 ;
    wire n474 ;
    wire n475 ;
    wire n476 ;
    wire n477 ;
    wire n478 ;
    wire n479 ;
    wire n480 ;
    wire n481 ;
    wire n482 ;
    wire n483 ;
    wire n484 ;
    wire n485 ;
    wire n486 ;
    wire n487 ;
    wire n488 ;
    wire n489 ;
    wire n490 ;
    wire n491 ;
    wire n492 ;
    wire n493 ;
    wire n494 ;
    wire n495 ;
    wire n496 ;
    wire n497 ;
    wire n498 ;
    wire n499 ;
    wire n500 ;
    wire n501 ;
    wire n502 ;
    wire n503 ;
    wire n504 ;
    wire n505 ;
    wire n506 ;
    wire n507 ;
    wire n508 ;
    wire n509 ;
    wire n510 ;
    wire n511 ;
    wire n512 ;
    wire n513 ;
    wire n514 ;
    wire n515 ;
    wire n516 ;
    wire n517 ;
    wire n518 ;
    wire n519 ;
    wire n520 ;
    wire n521 ;
    wire n522 ;
    wire n523 ;
    wire n524 ;
    wire n525 ;
    wire n526 ;
    wire n527 ;
    wire n528 ;
    wire n529 ;
    wire n530 ;
    wire n531 ;
    wire n532 ;
    wire n533 ;
    wire n534 ;
    wire n535 ;
    wire n536 ;
    wire n537 ;
    wire n538 ;
    wire [123:120] SUBSTITUTION ;
    wire [127:64] CONST_ADDITION ;
    wire [95:0] SHIFTROWS ;
    wire [3:0] S_0_R2 ;
    wire [3:0] S_0_R1 ;
    wire [3:0] S_1_R2 ;
    wire [3:0] S_1_R1 ;
    wire [3:0] S_2_R2 ;
    wire [3:0] S_2_R1 ;
    wire [3:0] S_3_R2 ;
    wire [3:0] S_3_R1 ;
    wire [3:0] S_4_R2 ;
    wire [3:0] S_4_R1 ;
    wire [3:0] S_5_R2 ;
    wire [3:0] S_5_R1 ;
    wire [3:0] S_6_R2 ;
    wire [3:0] S_6_R1 ;
    wire [3:0] S_7_R2 ;
    wire [3:0] S_7_R1 ;
    wire [3:0] S_8_R2 ;
    wire [3:0] S_8_R1 ;
    wire [3:0] S_9_R2 ;
    wire [3:0] S_9_R1 ;
    wire [3:0] S_10_R2 ;
    wire [3:0] S_10_R1 ;
    wire [3:0] S_11_R2 ;
    wire [3:0] S_11_R1 ;
    wire [3:0] S_12_R2 ;
    wire [3:0] S_12_R1 ;
    wire [3:0] S_13_R2 ;
    wire [3:0] S_13_R1 ;
    wire [3:0] S_14_R2 ;
    wire [3:0] S_14_R1 ;
    wire [3:0] S_15_R2 ;
    wire [3:0] S_15_R1 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) U400 ( .a ({ROUND_KEY_s3[227], ROUND_KEY_s2[227], ROUND_KEY_s1[227], ROUND_KEY_s0[227]}), .b ({ROUND_KEY_s3[99], ROUND_KEY_s2[99], ROUND_KEY_s1[99], ROUND_KEY_s0[99]}), .c ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, new_AGEMA_signal_1088, n406}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U403 ( .a ({ROUND_KEY_s3[226], ROUND_KEY_s2[226], ROUND_KEY_s1[226], ROUND_KEY_s0[226]}), .b ({ROUND_KEY_s3[98], ROUND_KEY_s2[98], ROUND_KEY_s1[98], ROUND_KEY_s0[98]}), .c ({new_AGEMA_signal_1099, new_AGEMA_signal_1098, new_AGEMA_signal_1097, n408}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U406 ( .a ({ROUND_KEY_s3[225], ROUND_KEY_s2[225], ROUND_KEY_s1[225], ROUND_KEY_s0[225]}), .b ({ROUND_KEY_s3[97], ROUND_KEY_s2[97], ROUND_KEY_s1[97], ROUND_KEY_s0[97]}), .c ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, n410}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U409 ( .a ({ROUND_KEY_s3[224], ROUND_KEY_s2[224], ROUND_KEY_s1[224], ROUND_KEY_s0[224]}), .b ({ROUND_KEY_s3[96], ROUND_KEY_s2[96], ROUND_KEY_s1[96], ROUND_KEY_s0[96]}), .c ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, new_AGEMA_signal_1115, n412}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U412 ( .a ({ROUND_KEY_s3[223], ROUND_KEY_s2[223], ROUND_KEY_s1[223], ROUND_KEY_s0[223]}), .b ({ROUND_KEY_s3[95], ROUND_KEY_s2[95], ROUND_KEY_s1[95], ROUND_KEY_s0[95]}), .c ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, new_AGEMA_signal_1124, n414}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U415 ( .a ({ROUND_KEY_s3[222], ROUND_KEY_s2[222], ROUND_KEY_s1[222], ROUND_KEY_s0[222]}), .b ({ROUND_KEY_s3[94], ROUND_KEY_s2[94], ROUND_KEY_s1[94], ROUND_KEY_s0[94]}), .c ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, new_AGEMA_signal_1133, n416}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U418 ( .a ({ROUND_KEY_s3[221], ROUND_KEY_s2[221], ROUND_KEY_s1[221], ROUND_KEY_s0[221]}), .b ({ROUND_KEY_s3[93], ROUND_KEY_s2[93], ROUND_KEY_s1[93], ROUND_KEY_s0[93]}), .c ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, new_AGEMA_signal_1142, n418}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U421 ( .a ({ROUND_KEY_s3[220], ROUND_KEY_s2[220], ROUND_KEY_s1[220], ROUND_KEY_s0[220]}), .b ({ROUND_KEY_s3[92], ROUND_KEY_s2[92], ROUND_KEY_s1[92], ROUND_KEY_s0[92]}), .c ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, n420}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U424 ( .a ({ROUND_KEY_s3[219], ROUND_KEY_s2[219], ROUND_KEY_s1[219], ROUND_KEY_s0[219]}), .b ({ROUND_KEY_s3[91], ROUND_KEY_s2[91], ROUND_KEY_s1[91], ROUND_KEY_s0[91]}), .c ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, new_AGEMA_signal_1160, n422}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U427 ( .a ({ROUND_KEY_s3[218], ROUND_KEY_s2[218], ROUND_KEY_s1[218], ROUND_KEY_s0[218]}), .b ({ROUND_KEY_s3[90], ROUND_KEY_s2[90], ROUND_KEY_s1[90], ROUND_KEY_s0[90]}), .c ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, new_AGEMA_signal_1169, n424}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U430 ( .a ({ROUND_KEY_s3[217], ROUND_KEY_s2[217], ROUND_KEY_s1[217], ROUND_KEY_s0[217]}), .b ({ROUND_KEY_s3[89], ROUND_KEY_s2[89], ROUND_KEY_s1[89], ROUND_KEY_s0[89]}), .c ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, n426}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U434 ( .a ({ROUND_KEY_s3[216], ROUND_KEY_s2[216], ROUND_KEY_s1[216], ROUND_KEY_s0[216]}), .b ({ROUND_KEY_s3[88], ROUND_KEY_s2[88], ROUND_KEY_s1[88], ROUND_KEY_s0[88]}), .c ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, new_AGEMA_signal_1187, n429}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U438 ( .a ({ROUND_KEY_s3[215], ROUND_KEY_s2[215], ROUND_KEY_s1[215], ROUND_KEY_s0[215]}), .b ({ROUND_KEY_s3[87], ROUND_KEY_s2[87], ROUND_KEY_s1[87], ROUND_KEY_s0[87]}), .c ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, new_AGEMA_signal_1196, n432}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U441 ( .a ({ROUND_KEY_s3[214], ROUND_KEY_s2[214], ROUND_KEY_s1[214], ROUND_KEY_s0[214]}), .b ({ROUND_KEY_s3[86], ROUND_KEY_s2[86], ROUND_KEY_s1[86], ROUND_KEY_s0[86]}), .c ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, new_AGEMA_signal_1205, n434}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U444 ( .a ({ROUND_KEY_s3[213], ROUND_KEY_s2[213], ROUND_KEY_s1[213], ROUND_KEY_s0[213]}), .b ({ROUND_KEY_s3[85], ROUND_KEY_s2[85], ROUND_KEY_s1[85], ROUND_KEY_s0[85]}), .c ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, new_AGEMA_signal_1214, n436}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U447 ( .a ({ROUND_KEY_s3[212], ROUND_KEY_s2[212], ROUND_KEY_s1[212], ROUND_KEY_s0[212]}), .b ({ROUND_KEY_s3[84], ROUND_KEY_s2[84], ROUND_KEY_s1[84], ROUND_KEY_s0[84]}), .c ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, n438}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U450 ( .a ({ROUND_KEY_s3[211], ROUND_KEY_s2[211], ROUND_KEY_s1[211], ROUND_KEY_s0[211]}), .b ({ROUND_KEY_s3[83], ROUND_KEY_s2[83], ROUND_KEY_s1[83], ROUND_KEY_s0[83]}), .c ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, new_AGEMA_signal_1232, n440}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U453 ( .a ({ROUND_KEY_s3[210], ROUND_KEY_s2[210], ROUND_KEY_s1[210], ROUND_KEY_s0[210]}), .b ({ROUND_KEY_s3[82], ROUND_KEY_s2[82], ROUND_KEY_s1[82], ROUND_KEY_s0[82]}), .c ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, new_AGEMA_signal_1241, n442}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U456 ( .a ({ROUND_KEY_s3[209], ROUND_KEY_s2[209], ROUND_KEY_s1[209], ROUND_KEY_s0[209]}), .b ({ROUND_KEY_s3[81], ROUND_KEY_s2[81], ROUND_KEY_s1[81], ROUND_KEY_s0[81]}), .c ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, new_AGEMA_signal_1250, n444}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U459 ( .a ({ROUND_KEY_s3[208], ROUND_KEY_s2[208], ROUND_KEY_s1[208], ROUND_KEY_s0[208]}), .b ({ROUND_KEY_s3[80], ROUND_KEY_s2[80], ROUND_KEY_s1[80], ROUND_KEY_s0[80]}), .c ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, new_AGEMA_signal_1259, n446}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U462 ( .a ({ROUND_KEY_s3[207], ROUND_KEY_s2[207], ROUND_KEY_s1[207], ROUND_KEY_s0[207]}), .b ({ROUND_KEY_s3[79], ROUND_KEY_s2[79], ROUND_KEY_s1[79], ROUND_KEY_s0[79]}), .c ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, new_AGEMA_signal_1268, n448}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U465 ( .a ({ROUND_KEY_s3[206], ROUND_KEY_s2[206], ROUND_KEY_s1[206], ROUND_KEY_s0[206]}), .b ({ROUND_KEY_s3[78], ROUND_KEY_s2[78], ROUND_KEY_s1[78], ROUND_KEY_s0[78]}), .c ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, new_AGEMA_signal_1277, n450}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U468 ( .a ({ROUND_KEY_s3[205], ROUND_KEY_s2[205], ROUND_KEY_s1[205], ROUND_KEY_s0[205]}), .b ({ROUND_KEY_s3[77], ROUND_KEY_s2[77], ROUND_KEY_s1[77], ROUND_KEY_s0[77]}), .c ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, n452}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U471 ( .a ({ROUND_KEY_s3[204], ROUND_KEY_s2[204], ROUND_KEY_s1[204], ROUND_KEY_s0[204]}), .b ({ROUND_KEY_s3[76], ROUND_KEY_s2[76], ROUND_KEY_s1[76], ROUND_KEY_s0[76]}), .c ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, new_AGEMA_signal_1295, n454}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U474 ( .a ({ROUND_KEY_s3[203], ROUND_KEY_s2[203], ROUND_KEY_s1[203], ROUND_KEY_s0[203]}), .b ({ROUND_KEY_s3[75], ROUND_KEY_s2[75], ROUND_KEY_s1[75], ROUND_KEY_s0[75]}), .c ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, new_AGEMA_signal_1304, n456}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U477 ( .a ({ROUND_KEY_s3[202], ROUND_KEY_s2[202], ROUND_KEY_s1[202], ROUND_KEY_s0[202]}), .b ({ROUND_KEY_s3[74], ROUND_KEY_s2[74], ROUND_KEY_s1[74], ROUND_KEY_s0[74]}), .c ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, new_AGEMA_signal_1313, n458}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U480 ( .a ({ROUND_KEY_s3[201], ROUND_KEY_s2[201], ROUND_KEY_s1[201], ROUND_KEY_s0[201]}), .b ({ROUND_KEY_s3[73], ROUND_KEY_s2[73], ROUND_KEY_s1[73], ROUND_KEY_s0[73]}), .c ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, n460}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U483 ( .a ({ROUND_KEY_s3[200], ROUND_KEY_s2[200], ROUND_KEY_s1[200], ROUND_KEY_s0[200]}), .b ({ROUND_KEY_s3[72], ROUND_KEY_s2[72], ROUND_KEY_s1[72], ROUND_KEY_s0[72]}), .c ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, n462}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U486 ( .a ({ROUND_KEY_s3[199], ROUND_KEY_s2[199], ROUND_KEY_s1[199], ROUND_KEY_s0[199]}), .b ({ROUND_KEY_s3[71], ROUND_KEY_s2[71], ROUND_KEY_s1[71], ROUND_KEY_s0[71]}), .c ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, new_AGEMA_signal_1340, n464}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U489 ( .a ({ROUND_KEY_s3[198], ROUND_KEY_s2[198], ROUND_KEY_s1[198], ROUND_KEY_s0[198]}), .b ({ROUND_KEY_s3[70], ROUND_KEY_s2[70], ROUND_KEY_s1[70], ROUND_KEY_s0[70]}), .c ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, new_AGEMA_signal_1349, n466}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U492 ( .a ({ROUND_KEY_s3[197], ROUND_KEY_s2[197], ROUND_KEY_s1[197], ROUND_KEY_s0[197]}), .b ({ROUND_KEY_s3[69], ROUND_KEY_s2[69], ROUND_KEY_s1[69], ROUND_KEY_s0[69]}), .c ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, new_AGEMA_signal_1358, n468}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U495 ( .a ({ROUND_KEY_s3[196], ROUND_KEY_s2[196], ROUND_KEY_s1[196], ROUND_KEY_s0[196]}), .b ({ROUND_KEY_s3[68], ROUND_KEY_s2[68], ROUND_KEY_s1[68], ROUND_KEY_s0[68]}), .c ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, n470}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U498 ( .a ({ROUND_KEY_s3[195], ROUND_KEY_s2[195], ROUND_KEY_s1[195], ROUND_KEY_s0[195]}), .b ({ROUND_KEY_s3[67], ROUND_KEY_s2[67], ROUND_KEY_s1[67], ROUND_KEY_s0[67]}), .c ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, new_AGEMA_signal_1376, n472}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U501 ( .a ({ROUND_KEY_s3[194], ROUND_KEY_s2[194], ROUND_KEY_s1[194], ROUND_KEY_s0[194]}), .b ({ROUND_KEY_s3[66], ROUND_KEY_s2[66], ROUND_KEY_s1[66], ROUND_KEY_s0[66]}), .c ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, new_AGEMA_signal_1385, n474}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U504 ( .a ({ROUND_KEY_s3[193], ROUND_KEY_s2[193], ROUND_KEY_s1[193], ROUND_KEY_s0[193]}), .b ({ROUND_KEY_s3[65], ROUND_KEY_s2[65], ROUND_KEY_s1[65], ROUND_KEY_s0[65]}), .c ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, n476}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U507 ( .a ({ROUND_KEY_s3[192], ROUND_KEY_s2[192], ROUND_KEY_s1[192], ROUND_KEY_s0[192]}), .b ({ROUND_KEY_s3[64], ROUND_KEY_s2[64], ROUND_KEY_s1[64], ROUND_KEY_s0[64]}), .c ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, new_AGEMA_signal_1403, n478}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U510 ( .a ({ROUND_KEY_s3[127], ROUND_KEY_s2[127], ROUND_KEY_s1[127], ROUND_KEY_s0[127]}), .b ({ROUND_KEY_s3[255], ROUND_KEY_s2[255], ROUND_KEY_s1[255], ROUND_KEY_s0[255]}), .c ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, new_AGEMA_signal_1412, n480}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U513 ( .a ({ROUND_KEY_s3[126], ROUND_KEY_s2[126], ROUND_KEY_s1[126], ROUND_KEY_s0[126]}), .b ({ROUND_KEY_s3[254], ROUND_KEY_s2[254], ROUND_KEY_s1[254], ROUND_KEY_s0[254]}), .c ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, new_AGEMA_signal_1421, n482}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U516 ( .a ({ROUND_KEY_s3[125], ROUND_KEY_s2[125], ROUND_KEY_s1[125], ROUND_KEY_s0[125]}), .b ({ROUND_KEY_s3[253], ROUND_KEY_s2[253], ROUND_KEY_s1[253], ROUND_KEY_s0[253]}), .c ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, new_AGEMA_signal_1430, n484}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U519 ( .a ({ROUND_KEY_s3[124], ROUND_KEY_s2[124], ROUND_KEY_s1[124], ROUND_KEY_s0[124]}), .b ({ROUND_KEY_s3[252], ROUND_KEY_s2[252], ROUND_KEY_s1[252], ROUND_KEY_s0[252]}), .c ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, n486}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U522 ( .a ({ROUND_KEY_s3[123], ROUND_KEY_s2[123], ROUND_KEY_s1[123], ROUND_KEY_s0[123]}), .b ({ROUND_KEY_s3[251], ROUND_KEY_s2[251], ROUND_KEY_s1[251], ROUND_KEY_s0[251]}), .c ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, new_AGEMA_signal_1448, n488}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U526 ( .a ({ROUND_KEY_s3[122], ROUND_KEY_s2[122], ROUND_KEY_s1[122], ROUND_KEY_s0[122]}), .b ({ROUND_KEY_s3[250], ROUND_KEY_s2[250], ROUND_KEY_s1[250], ROUND_KEY_s0[250]}), .c ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, new_AGEMA_signal_1457, n491}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U530 ( .a ({ROUND_KEY_s3[121], ROUND_KEY_s2[121], ROUND_KEY_s1[121], ROUND_KEY_s0[121]}), .b ({ROUND_KEY_s3[249], ROUND_KEY_s2[249], ROUND_KEY_s1[249], ROUND_KEY_s0[249]}), .c ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, new_AGEMA_signal_1466, n494}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U534 ( .a ({ROUND_KEY_s3[120], ROUND_KEY_s2[120], ROUND_KEY_s1[120], ROUND_KEY_s0[120]}), .b ({ROUND_KEY_s3[248], ROUND_KEY_s2[248], ROUND_KEY_s1[248], ROUND_KEY_s0[248]}), .c ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, new_AGEMA_signal_1475, n497}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U538 ( .a ({ROUND_KEY_s3[119], ROUND_KEY_s2[119], ROUND_KEY_s1[119], ROUND_KEY_s0[119]}), .b ({ROUND_KEY_s3[247], ROUND_KEY_s2[247], ROUND_KEY_s1[247], ROUND_KEY_s0[247]}), .c ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, new_AGEMA_signal_1484, n500}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U541 ( .a ({ROUND_KEY_s3[118], ROUND_KEY_s2[118], ROUND_KEY_s1[118], ROUND_KEY_s0[118]}), .b ({ROUND_KEY_s3[246], ROUND_KEY_s2[246], ROUND_KEY_s1[246], ROUND_KEY_s0[246]}), .c ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, new_AGEMA_signal_1493, n502}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U544 ( .a ({ROUND_KEY_s3[117], ROUND_KEY_s2[117], ROUND_KEY_s1[117], ROUND_KEY_s0[117]}), .b ({ROUND_KEY_s3[245], ROUND_KEY_s2[245], ROUND_KEY_s1[245], ROUND_KEY_s0[245]}), .c ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, new_AGEMA_signal_1502, n504}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U547 ( .a ({ROUND_KEY_s3[116], ROUND_KEY_s2[116], ROUND_KEY_s1[116], ROUND_KEY_s0[116]}), .b ({ROUND_KEY_s3[244], ROUND_KEY_s2[244], ROUND_KEY_s1[244], ROUND_KEY_s0[244]}), .c ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, new_AGEMA_signal_1511, n506}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U550 ( .a ({ROUND_KEY_s3[115], ROUND_KEY_s2[115], ROUND_KEY_s1[115], ROUND_KEY_s0[115]}), .b ({ROUND_KEY_s3[243], ROUND_KEY_s2[243], ROUND_KEY_s1[243], ROUND_KEY_s0[243]}), .c ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, new_AGEMA_signal_1520, n508}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U553 ( .a ({ROUND_KEY_s3[114], ROUND_KEY_s2[114], ROUND_KEY_s1[114], ROUND_KEY_s0[114]}), .b ({ROUND_KEY_s3[242], ROUND_KEY_s2[242], ROUND_KEY_s1[242], ROUND_KEY_s0[242]}), .c ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, new_AGEMA_signal_1529, n510}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U556 ( .a ({ROUND_KEY_s3[113], ROUND_KEY_s2[113], ROUND_KEY_s1[113], ROUND_KEY_s0[113]}), .b ({ROUND_KEY_s3[241], ROUND_KEY_s2[241], ROUND_KEY_s1[241], ROUND_KEY_s0[241]}), .c ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, new_AGEMA_signal_1538, n512}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U559 ( .a ({ROUND_KEY_s3[112], ROUND_KEY_s2[112], ROUND_KEY_s1[112], ROUND_KEY_s0[112]}), .b ({ROUND_KEY_s3[240], ROUND_KEY_s2[240], ROUND_KEY_s1[240], ROUND_KEY_s0[240]}), .c ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, new_AGEMA_signal_1547, n514}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U562 ( .a ({ROUND_KEY_s3[111], ROUND_KEY_s2[111], ROUND_KEY_s1[111], ROUND_KEY_s0[111]}), .b ({ROUND_KEY_s3[239], ROUND_KEY_s2[239], ROUND_KEY_s1[239], ROUND_KEY_s0[239]}), .c ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, new_AGEMA_signal_1556, n516}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U565 ( .a ({ROUND_KEY_s3[110], ROUND_KEY_s2[110], ROUND_KEY_s1[110], ROUND_KEY_s0[110]}), .b ({ROUND_KEY_s3[238], ROUND_KEY_s2[238], ROUND_KEY_s1[238], ROUND_KEY_s0[238]}), .c ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, new_AGEMA_signal_1565, n518}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U568 ( .a ({ROUND_KEY_s3[109], ROUND_KEY_s2[109], ROUND_KEY_s1[109], ROUND_KEY_s0[109]}), .b ({ROUND_KEY_s3[237], ROUND_KEY_s2[237], ROUND_KEY_s1[237], ROUND_KEY_s0[237]}), .c ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1574, n520}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U571 ( .a ({ROUND_KEY_s3[108], ROUND_KEY_s2[108], ROUND_KEY_s1[108], ROUND_KEY_s0[108]}), .b ({ROUND_KEY_s3[236], ROUND_KEY_s2[236], ROUND_KEY_s1[236], ROUND_KEY_s0[236]}), .c ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, new_AGEMA_signal_1583, n522}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U574 ( .a ({ROUND_KEY_s3[107], ROUND_KEY_s2[107], ROUND_KEY_s1[107], ROUND_KEY_s0[107]}), .b ({ROUND_KEY_s3[235], ROUND_KEY_s2[235], ROUND_KEY_s1[235], ROUND_KEY_s0[235]}), .c ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, new_AGEMA_signal_1592, n524}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U577 ( .a ({ROUND_KEY_s3[106], ROUND_KEY_s2[106], ROUND_KEY_s1[106], ROUND_KEY_s0[106]}), .b ({ROUND_KEY_s3[234], ROUND_KEY_s2[234], ROUND_KEY_s1[234], ROUND_KEY_s0[234]}), .c ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, new_AGEMA_signal_1601, n526}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U580 ( .a ({ROUND_KEY_s3[105], ROUND_KEY_s2[105], ROUND_KEY_s1[105], ROUND_KEY_s0[105]}), .b ({ROUND_KEY_s3[233], ROUND_KEY_s2[233], ROUND_KEY_s1[233], ROUND_KEY_s0[233]}), .c ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1610, n528}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U583 ( .a ({ROUND_KEY_s3[104], ROUND_KEY_s2[104], ROUND_KEY_s1[104], ROUND_KEY_s0[104]}), .b ({ROUND_KEY_s3[232], ROUND_KEY_s2[232], ROUND_KEY_s1[232], ROUND_KEY_s0[232]}), .c ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, new_AGEMA_signal_1619, n530}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U586 ( .a ({ROUND_KEY_s3[103], ROUND_KEY_s2[103], ROUND_KEY_s1[103], ROUND_KEY_s0[103]}), .b ({ROUND_KEY_s3[231], ROUND_KEY_s2[231], ROUND_KEY_s1[231], ROUND_KEY_s0[231]}), .c ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, new_AGEMA_signal_1628, n532}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U589 ( .a ({ROUND_KEY_s3[102], ROUND_KEY_s2[102], ROUND_KEY_s1[102], ROUND_KEY_s0[102]}), .b ({ROUND_KEY_s3[230], ROUND_KEY_s2[230], ROUND_KEY_s1[230], ROUND_KEY_s0[230]}), .c ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, new_AGEMA_signal_1637, n534}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U592 ( .a ({ROUND_KEY_s3[101], ROUND_KEY_s2[101], ROUND_KEY_s1[101], ROUND_KEY_s0[101]}), .b ({ROUND_KEY_s3[229], ROUND_KEY_s2[229], ROUND_KEY_s1[229], ROUND_KEY_s0[229]}), .c ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1646, n536}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U595 ( .a ({ROUND_KEY_s3[100], ROUND_KEY_s2[100], ROUND_KEY_s1[100], ROUND_KEY_s0[100]}), .b ({ROUND_KEY_s3[228], ROUND_KEY_s2[228], ROUND_KEY_s1[228], ROUND_KEY_s0[228]}), .c ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, new_AGEMA_signal_1655, n538}) ) ;
    //ClockGatingController #(8) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U404 ( .a ({ROUND_KEY_s3[354], ROUND_KEY_s2[354], ROUND_KEY_s1[354], ROUND_KEY_s0[354]}), .b ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, CONST_ADDITION[98]}), .c ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, new_AGEMA_signal_2285, n407}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U405 ( .a ({new_AGEMA_signal_1099, new_AGEMA_signal_1098, new_AGEMA_signal_1097, n408}), .b ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, new_AGEMA_signal_2285, n407}), .c ({ROUND_OUT_s3[66], ROUND_OUT_s2[66], ROUND_OUT_s1[66], ROUND_OUT_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U416 ( .a ({ROUND_KEY_s3[350], ROUND_KEY_s2[350], ROUND_KEY_s1[350], ROUND_KEY_s0[350]}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, new_AGEMA_signal_2219, CONST_ADDITION[94]}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, new_AGEMA_signal_2291, n415}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U417 ( .a ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, new_AGEMA_signal_1133, n416}), .b ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, new_AGEMA_signal_2291, n415}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, new_AGEMA_signal_2525, SHIFTROWS[86]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U419 ( .a ({ROUND_KEY_s3[349], ROUND_KEY_s2[349], ROUND_KEY_s1[349], ROUND_KEY_s0[349]}), .b ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, new_AGEMA_signal_2213, CONST_ADDITION[93]}), .c ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, new_AGEMA_signal_2297, n417}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U420 ( .a ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, new_AGEMA_signal_1142, n418}), .b ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, new_AGEMA_signal_2297, n417}), .c ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, new_AGEMA_signal_2528, SHIFTROWS[85]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U428 ( .a ({ROUND_KEY_s3[346], ROUND_KEY_s2[346], ROUND_KEY_s1[346], ROUND_KEY_s0[346]}), .b ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, new_AGEMA_signal_2207, CONST_ADDITION[90]}), .c ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, new_AGEMA_signal_2303, n423}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U429 ( .a ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, new_AGEMA_signal_1169, n424}), .b ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, new_AGEMA_signal_2303, n423}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, new_AGEMA_signal_2531, SHIFTROWS[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U442 ( .a ({ROUND_KEY_s3[342], ROUND_KEY_s2[342], ROUND_KEY_s1[342], ROUND_KEY_s0[342]}), .b ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, new_AGEMA_signal_2204, CONST_ADDITION[86]}), .c ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, new_AGEMA_signal_2309, n433}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U443 ( .a ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, new_AGEMA_signal_1205, n434}), .b ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, new_AGEMA_signal_2309, n433}), .c ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, new_AGEMA_signal_2534, SHIFTROWS[78]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U445 ( .a ({ROUND_KEY_s3[341], ROUND_KEY_s2[341], ROUND_KEY_s1[341], ROUND_KEY_s0[341]}), .b ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, new_AGEMA_signal_2198, CONST_ADDITION[85]}), .c ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, new_AGEMA_signal_2315, n435}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U446 ( .a ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, new_AGEMA_signal_1214, n436}), .b ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, new_AGEMA_signal_2315, n435}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, new_AGEMA_signal_2537, SHIFTROWS[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U454 ( .a ({ROUND_KEY_s3[338], ROUND_KEY_s2[338], ROUND_KEY_s1[338], ROUND_KEY_s0[338]}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, new_AGEMA_signal_2192, CONST_ADDITION[82]}), .c ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, new_AGEMA_signal_2321, n441}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U455 ( .a ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, new_AGEMA_signal_1241, n442}), .b ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, new_AGEMA_signal_2321, n441}), .c ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, new_AGEMA_signal_2540, SHIFTROWS[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U466 ( .a ({ROUND_KEY_s3[334], ROUND_KEY_s2[334], ROUND_KEY_s1[334], ROUND_KEY_s0[334]}), .b ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, CONST_ADDITION[78]}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, n449}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U467 ( .a ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, new_AGEMA_signal_1277, n450}), .b ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, n449}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, new_AGEMA_signal_2543, SHIFTROWS[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U469 ( .a ({ROUND_KEY_s3[333], ROUND_KEY_s2[333], ROUND_KEY_s1[333], ROUND_KEY_s0[333]}), .b ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, CONST_ADDITION[77]}), .c ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, new_AGEMA_signal_2333, n451}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U470 ( .a ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, new_AGEMA_signal_1286, n452}), .b ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, new_AGEMA_signal_2333, n451}), .c ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, new_AGEMA_signal_2546, SHIFTROWS[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U478 ( .a ({ROUND_KEY_s3[330], ROUND_KEY_s2[330], ROUND_KEY_s1[330], ROUND_KEY_s0[330]}), .b ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, CONST_ADDITION[74]}), .c ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, new_AGEMA_signal_2339, n457}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U479 ( .a ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, new_AGEMA_signal_1313, n458}), .b ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, new_AGEMA_signal_2339, n457}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, new_AGEMA_signal_2549, SHIFTROWS[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U490 ( .a ({ROUND_KEY_s3[326], ROUND_KEY_s2[326], ROUND_KEY_s1[326], ROUND_KEY_s0[326]}), .b ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, CONST_ADDITION[70]}), .c ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, new_AGEMA_signal_2345, n465}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U491 ( .a ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, new_AGEMA_signal_1349, n466}), .b ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, new_AGEMA_signal_2345, n465}), .c ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, new_AGEMA_signal_2552, SHIFTROWS[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U493 ( .a ({ROUND_KEY_s3[325], ROUND_KEY_s2[325], ROUND_KEY_s1[325], ROUND_KEY_s0[325]}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, new_AGEMA_signal_2168, CONST_ADDITION[69]}), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, new_AGEMA_signal_2351, n467}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U494 ( .a ({new_AGEMA_signal_1360, new_AGEMA_signal_1359, new_AGEMA_signal_1358, n468}), .b ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, new_AGEMA_signal_2351, n467}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, new_AGEMA_signal_2555, SHIFTROWS[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U502 ( .a ({ROUND_KEY_s3[322], ROUND_KEY_s2[322], ROUND_KEY_s1[322], ROUND_KEY_s0[322]}), .b ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, CONST_ADDITION[66]}), .c ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, new_AGEMA_signal_2357, n473}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U503 ( .a ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, new_AGEMA_signal_1385, n474}), .b ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, new_AGEMA_signal_2357, n473}), .c ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, SHIFTROWS[90]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U514 ( .a ({ROUND_KEY_s3[382], ROUND_KEY_s2[382], ROUND_KEY_s1[382], ROUND_KEY_s0[382]}), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, CONST_ADDITION[126]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, new_AGEMA_signal_2363, n481}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U515 ( .a ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, new_AGEMA_signal_1421, n482}), .b ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, new_AGEMA_signal_2363, n481}), .c ({ROUND_OUT_s3[94], ROUND_OUT_s2[94], ROUND_OUT_s1[94], ROUND_OUT_s0[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U517 ( .a ({ROUND_KEY_s3[381], ROUND_KEY_s2[381], ROUND_KEY_s1[381], ROUND_KEY_s0[381]}), .b ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, new_AGEMA_signal_2273, CONST_ADDITION[125]}), .c ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, new_AGEMA_signal_2369, n483}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U518 ( .a ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, new_AGEMA_signal_1430, n484}), .b ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, new_AGEMA_signal_2369, n483}), .c ({ROUND_OUT_s3[93], ROUND_OUT_s2[93], ROUND_OUT_s1[93], ROUND_OUT_s0[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U527 ( .a ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, new_AGEMA_signal_2267, SUBSTITUTION[122]}), .b ({ROUND_KEY_s3[378], ROUND_KEY_s2[378], ROUND_KEY_s1[378], ROUND_KEY_s0[378]}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, new_AGEMA_signal_2375, n490}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U528 ( .a ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, new_AGEMA_signal_1457, n491}), .b ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, new_AGEMA_signal_2375, n490}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, n492}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U529 ( .a ({1'b0, 1'b0, 1'b0, CONST_IN[2]}), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, new_AGEMA_signal_2567, n492}), .c ({ROUND_OUT_s3[90], ROUND_OUT_s2[90], ROUND_OUT_s1[90], ROUND_OUT_s0[90]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U542 ( .a ({ROUND_KEY_s3[374], ROUND_KEY_s2[374], ROUND_KEY_s1[374], ROUND_KEY_s0[374]}), .b ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, new_AGEMA_signal_2264, CONST_ADDITION[118]}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, n501}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U543 ( .a ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, new_AGEMA_signal_1493, n502}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, n501}), .c ({ROUND_OUT_s3[86], ROUND_OUT_s2[86], ROUND_OUT_s1[86], ROUND_OUT_s0[86]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U545 ( .a ({ROUND_KEY_s3[373], ROUND_KEY_s2[373], ROUND_KEY_s1[373], ROUND_KEY_s0[373]}), .b ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, CONST_ADDITION[117]}), .c ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, new_AGEMA_signal_2387, n503}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U546 ( .a ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, new_AGEMA_signal_1502, n504}), .b ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, new_AGEMA_signal_2387, n503}), .c ({ROUND_OUT_s3[85], ROUND_OUT_s2[85], ROUND_OUT_s1[85], ROUND_OUT_s0[85]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U554 ( .a ({ROUND_KEY_s3[370], ROUND_KEY_s2[370], ROUND_KEY_s1[370], ROUND_KEY_s0[370]}), .b ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, new_AGEMA_signal_2252, CONST_ADDITION[114]}), .c ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, new_AGEMA_signal_2393, n509}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U555 ( .a ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, new_AGEMA_signal_1529, n510}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, new_AGEMA_signal_2393, n509}), .c ({ROUND_OUT_s3[82], ROUND_OUT_s2[82], ROUND_OUT_s1[82], ROUND_OUT_s0[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U566 ( .a ({ROUND_KEY_s3[366], ROUND_KEY_s2[366], ROUND_KEY_s1[366], ROUND_KEY_s0[366]}), .b ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, new_AGEMA_signal_2249, CONST_ADDITION[110]}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, n517}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U567 ( .a ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, new_AGEMA_signal_1565, n518}), .b ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, n517}), .c ({ROUND_OUT_s3[78], ROUND_OUT_s2[78], ROUND_OUT_s1[78], ROUND_OUT_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U569 ( .a ({ROUND_KEY_s3[365], ROUND_KEY_s2[365], ROUND_KEY_s1[365], ROUND_KEY_s0[365]}), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, CONST_ADDITION[109]}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, new_AGEMA_signal_2405, n519}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U570 ( .a ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1574, n520}), .b ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, new_AGEMA_signal_2405, n519}), .c ({ROUND_OUT_s3[77], ROUND_OUT_s2[77], ROUND_OUT_s1[77], ROUND_OUT_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U578 ( .a ({ROUND_KEY_s3[362], ROUND_KEY_s2[362], ROUND_KEY_s1[362], ROUND_KEY_s0[362]}), .b ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, new_AGEMA_signal_2237, CONST_ADDITION[106]}), .c ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, new_AGEMA_signal_2411, n525}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U579 ( .a ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, new_AGEMA_signal_1601, n526}), .b ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, new_AGEMA_signal_2411, n525}), .c ({ROUND_OUT_s3[74], ROUND_OUT_s2[74], ROUND_OUT_s1[74], ROUND_OUT_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U590 ( .a ({ROUND_KEY_s3[358], ROUND_KEY_s2[358], ROUND_KEY_s1[358], ROUND_KEY_s0[358]}), .b ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, CONST_ADDITION[102]}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, new_AGEMA_signal_2417, n533}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U591 ( .a ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, new_AGEMA_signal_1637, n534}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, new_AGEMA_signal_2417, n533}), .c ({ROUND_OUT_s3[70], ROUND_OUT_s2[70], ROUND_OUT_s1[70], ROUND_OUT_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U593 ( .a ({ROUND_KEY_s3[357], ROUND_KEY_s2[357], ROUND_KEY_s1[357], ROUND_KEY_s0[357]}), .b ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, new_AGEMA_signal_2228, CONST_ADDITION[101]}), .c ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, new_AGEMA_signal_2423, n535}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U594 ( .a ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1646, n536}), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, new_AGEMA_signal_2423, n535}), .c ({ROUND_OUT_s3[69], ROUND_OUT_s2[69], ROUND_OUT_s1[69], ROUND_OUT_s0[69]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_0_U6 ( .a ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, S_0_R1[1]}), .b ({ROUND_IN_s3[6], ROUND_IN_s2[6], ROUND_IN_s1[6], ROUND_IN_s0[6]}), .c ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, SHIFTROWS[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_0_U3 ( .a ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, new_AGEMA_signal_1673, S_0_R2[0]}), .b ({ROUND_IN_s3[0], ROUND_IN_s2[0], ROUND_IN_s1[0], ROUND_IN_s0[0]}), .c ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, SHIFTROWS[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_0_U2 ( .a ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, new_AGEMA_signal_1664, S_0_R1[0]}), .b ({ROUND_IN_s3[4], ROUND_IN_s2[4], ROUND_IN_s1[4], ROUND_IN_s0[4]}), .c ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, SHIFTROWS[14]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_0_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[6], ROUND_IN_s2[6], ROUND_IN_s1[6], ROUND_IN_s0[6]}), .b ({ROUND_IN_s3[7], ROUND_IN_s2[7], ROUND_IN_s1[7], ROUND_IN_s0[7]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, new_AGEMA_signal_1664, S_0_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_0_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[2], ROUND_IN_s2[2], ROUND_IN_s1[2], ROUND_IN_s0[2]}), .b ({ROUND_IN_s3[3], ROUND_IN_s2[3], ROUND_IN_s1[3], ROUND_IN_s0[3]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, new_AGEMA_signal_1673, S_0_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_0_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[1], ROUND_IN_s2[1], ROUND_IN_s1[1], ROUND_IN_s0[1]}), .b ({ROUND_IN_s3[2], ROUND_IN_s2[2], ROUND_IN_s1[2], ROUND_IN_s0[2]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, S_0_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_1_U6 ( .a ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1703, S_1_R1[1]}), .b ({ROUND_IN_s3[14], ROUND_IN_s2[14], ROUND_IN_s1[14], ROUND_IN_s0[14]}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, new_AGEMA_signal_2057, SHIFTROWS[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_1_U3 ( .a ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, new_AGEMA_signal_1697, S_1_R2[0]}), .b ({ROUND_IN_s3[8], ROUND_IN_s2[8], ROUND_IN_s1[8], ROUND_IN_s0[8]}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, SHIFTROWS[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_1_U2 ( .a ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, new_AGEMA_signal_1688, S_1_R1[0]}), .b ({ROUND_IN_s3[12], ROUND_IN_s2[12], ROUND_IN_s1[12], ROUND_IN_s0[12]}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, SHIFTROWS[22]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_1_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[14], ROUND_IN_s2[14], ROUND_IN_s1[14], ROUND_IN_s0[14]}), .b ({ROUND_IN_s3[15], ROUND_IN_s2[15], ROUND_IN_s1[15], ROUND_IN_s0[15]}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, new_AGEMA_signal_1688, S_1_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_1_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[10], ROUND_IN_s2[10], ROUND_IN_s1[10], ROUND_IN_s0[10]}), .b ({ROUND_IN_s3[11], ROUND_IN_s2[11], ROUND_IN_s1[11], ROUND_IN_s0[11]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, new_AGEMA_signal_1697, S_1_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_1_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[9], ROUND_IN_s2[9], ROUND_IN_s1[9], ROUND_IN_s0[9]}), .b ({ROUND_IN_s3[10], ROUND_IN_s2[10], ROUND_IN_s1[10], ROUND_IN_s0[10]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1703, S_1_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_2_U6 ( .a ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, new_AGEMA_signal_1727, S_2_R1[1]}), .b ({ROUND_IN_s3[22], ROUND_IN_s2[22], ROUND_IN_s1[22], ROUND_IN_s0[22]}), .c ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, SHIFTROWS[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_2_U3 ( .a ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, new_AGEMA_signal_1721, S_2_R2[0]}), .b ({ROUND_IN_s3[16], ROUND_IN_s2[16], ROUND_IN_s1[16], ROUND_IN_s0[16]}), .c ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, SHIFTROWS[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_2_U2 ( .a ({new_AGEMA_signal_1714, new_AGEMA_signal_1713, new_AGEMA_signal_1712, S_2_R1[0]}), .b ({ROUND_IN_s3[20], ROUND_IN_s2[20], ROUND_IN_s1[20], ROUND_IN_s0[20]}), .c ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, SHIFTROWS[30]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_2_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[22], ROUND_IN_s2[22], ROUND_IN_s1[22], ROUND_IN_s0[22]}), .b ({ROUND_IN_s3[23], ROUND_IN_s2[23], ROUND_IN_s1[23], ROUND_IN_s0[23]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1714, new_AGEMA_signal_1713, new_AGEMA_signal_1712, S_2_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_2_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[18], ROUND_IN_s2[18], ROUND_IN_s1[18], ROUND_IN_s0[18]}), .b ({ROUND_IN_s3[19], ROUND_IN_s2[19], ROUND_IN_s1[19], ROUND_IN_s0[19]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, new_AGEMA_signal_1721, S_2_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_2_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[17], ROUND_IN_s2[17], ROUND_IN_s1[17], ROUND_IN_s0[17]}), .b ({ROUND_IN_s3[18], ROUND_IN_s2[18], ROUND_IN_s1[18], ROUND_IN_s0[18]}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, new_AGEMA_signal_1727, S_2_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_3_U6 ( .a ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, S_3_R1[1]}), .b ({ROUND_IN_s3[30], ROUND_IN_s2[30], ROUND_IN_s1[30], ROUND_IN_s0[30]}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, SHIFTROWS[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_3_U3 ( .a ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, new_AGEMA_signal_1745, S_3_R2[0]}), .b ({ROUND_IN_s3[24], ROUND_IN_s2[24], ROUND_IN_s1[24], ROUND_IN_s0[24]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, SHIFTROWS[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_3_U2 ( .a ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, new_AGEMA_signal_1736, S_3_R1[0]}), .b ({ROUND_IN_s3[28], ROUND_IN_s2[28], ROUND_IN_s1[28], ROUND_IN_s0[28]}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, SHIFTROWS[6]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_3_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[30], ROUND_IN_s2[30], ROUND_IN_s1[30], ROUND_IN_s0[30]}), .b ({ROUND_IN_s3[31], ROUND_IN_s2[31], ROUND_IN_s1[31], ROUND_IN_s0[31]}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, new_AGEMA_signal_1736, S_3_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_3_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[26], ROUND_IN_s2[26], ROUND_IN_s1[26], ROUND_IN_s0[26]}), .b ({ROUND_IN_s3[27], ROUND_IN_s2[27], ROUND_IN_s1[27], ROUND_IN_s0[27]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, new_AGEMA_signal_1745, S_3_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_3_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[25], ROUND_IN_s2[25], ROUND_IN_s1[25], ROUND_IN_s0[25]}), .b ({ROUND_IN_s3[26], ROUND_IN_s2[26], ROUND_IN_s1[26], ROUND_IN_s0[26]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, S_3_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_4_U6 ( .a ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, new_AGEMA_signal_1775, S_4_R1[1]}), .b ({ROUND_IN_s3[38], ROUND_IN_s2[38], ROUND_IN_s1[38], ROUND_IN_s0[38]}), .c ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, SHIFTROWS[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_4_U3 ( .a ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, new_AGEMA_signal_1769, S_4_R2[0]}), .b ({ROUND_IN_s3[32], ROUND_IN_s2[32], ROUND_IN_s1[32], ROUND_IN_s0[32]}), .c ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, SHIFTROWS[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_4_U2 ( .a ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, new_AGEMA_signal_1760, S_4_R1[0]}), .b ({ROUND_IN_s3[36], ROUND_IN_s2[36], ROUND_IN_s1[36], ROUND_IN_s0[36]}), .c ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, new_AGEMA_signal_2114, SHIFTROWS[54]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_4_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[38], ROUND_IN_s2[38], ROUND_IN_s1[38], ROUND_IN_s0[38]}), .b ({ROUND_IN_s3[39], ROUND_IN_s2[39], ROUND_IN_s1[39], ROUND_IN_s0[39]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, new_AGEMA_signal_1760, S_4_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_4_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[34], ROUND_IN_s2[34], ROUND_IN_s1[34], ROUND_IN_s0[34]}), .b ({ROUND_IN_s3[35], ROUND_IN_s2[35], ROUND_IN_s1[35], ROUND_IN_s0[35]}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, new_AGEMA_signal_1769, S_4_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_4_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[33], ROUND_IN_s2[33], ROUND_IN_s1[33], ROUND_IN_s0[33]}), .b ({ROUND_IN_s3[34], ROUND_IN_s2[34], ROUND_IN_s1[34], ROUND_IN_s0[34]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, new_AGEMA_signal_1775, S_4_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_5_U6 ( .a ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, new_AGEMA_signal_1799, S_5_R1[1]}), .b ({ROUND_IN_s3[46], ROUND_IN_s2[46], ROUND_IN_s1[46], ROUND_IN_s0[46]}), .c ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, new_AGEMA_signal_2117, SHIFTROWS[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_5_U3 ( .a ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, new_AGEMA_signal_1793, S_5_R2[0]}), .b ({ROUND_IN_s3[40], ROUND_IN_s2[40], ROUND_IN_s1[40], ROUND_IN_s0[40]}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, new_AGEMA_signal_2123, SHIFTROWS[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_5_U2 ( .a ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, new_AGEMA_signal_1784, S_5_R1[0]}), .b ({ROUND_IN_s3[44], ROUND_IN_s2[44], ROUND_IN_s1[44], ROUND_IN_s0[44]}), .c ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, new_AGEMA_signal_2129, SHIFTROWS[62]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_5_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[46], ROUND_IN_s2[46], ROUND_IN_s1[46], ROUND_IN_s0[46]}), .b ({ROUND_IN_s3[47], ROUND_IN_s2[47], ROUND_IN_s1[47], ROUND_IN_s0[47]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, new_AGEMA_signal_1784, S_5_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_5_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[42], ROUND_IN_s2[42], ROUND_IN_s1[42], ROUND_IN_s0[42]}), .b ({ROUND_IN_s3[43], ROUND_IN_s2[43], ROUND_IN_s1[43], ROUND_IN_s0[43]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, new_AGEMA_signal_1793, S_5_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_5_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[41], ROUND_IN_s2[41], ROUND_IN_s1[41], ROUND_IN_s0[41]}), .b ({ROUND_IN_s3[42], ROUND_IN_s2[42], ROUND_IN_s1[42], ROUND_IN_s0[42]}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, new_AGEMA_signal_1799, S_5_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_6_U6 ( .a ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, new_AGEMA_signal_1823, S_6_R1[1]}), .b ({ROUND_IN_s3[54], ROUND_IN_s2[54], ROUND_IN_s1[54], ROUND_IN_s0[54]}), .c ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, new_AGEMA_signal_2132, SHIFTROWS[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_6_U3 ( .a ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, new_AGEMA_signal_1817, S_6_R2[0]}), .b ({ROUND_IN_s3[48], ROUND_IN_s2[48], ROUND_IN_s1[48], ROUND_IN_s0[48]}), .c ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, new_AGEMA_signal_2138, SHIFTROWS[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_6_U2 ( .a ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, new_AGEMA_signal_1808, S_6_R1[0]}), .b ({ROUND_IN_s3[52], ROUND_IN_s2[52], ROUND_IN_s1[52], ROUND_IN_s0[52]}), .c ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, SHIFTROWS[38]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_6_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[54], ROUND_IN_s2[54], ROUND_IN_s1[54], ROUND_IN_s0[54]}), .b ({ROUND_IN_s3[55], ROUND_IN_s2[55], ROUND_IN_s1[55], ROUND_IN_s0[55]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, new_AGEMA_signal_1808, S_6_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_6_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[50], ROUND_IN_s2[50], ROUND_IN_s1[50], ROUND_IN_s0[50]}), .b ({ROUND_IN_s3[51], ROUND_IN_s2[51], ROUND_IN_s1[51], ROUND_IN_s0[51]}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, new_AGEMA_signal_1817, S_6_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_6_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[49], ROUND_IN_s2[49], ROUND_IN_s1[49], ROUND_IN_s0[49]}), .b ({ROUND_IN_s3[50], ROUND_IN_s2[50], ROUND_IN_s1[50], ROUND_IN_s0[50]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, new_AGEMA_signal_1823, S_6_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_7_U6 ( .a ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1847, S_7_R1[1]}), .b ({ROUND_IN_s3[62], ROUND_IN_s2[62], ROUND_IN_s1[62], ROUND_IN_s0[62]}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, new_AGEMA_signal_2147, SHIFTROWS[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_7_U3 ( .a ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, new_AGEMA_signal_1841, S_7_R2[0]}), .b ({ROUND_IN_s3[56], ROUND_IN_s2[56], ROUND_IN_s1[56], ROUND_IN_s0[56]}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, SHIFTROWS[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_7_U2 ( .a ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, new_AGEMA_signal_1832, S_7_R1[0]}), .b ({ROUND_IN_s3[60], ROUND_IN_s2[60], ROUND_IN_s1[60], ROUND_IN_s0[60]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, new_AGEMA_signal_2159, SHIFTROWS[46]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_7_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[62], ROUND_IN_s2[62], ROUND_IN_s1[62], ROUND_IN_s0[62]}), .b ({ROUND_IN_s3[63], ROUND_IN_s2[63], ROUND_IN_s1[63], ROUND_IN_s0[63]}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, new_AGEMA_signal_1832, S_7_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_7_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[58], ROUND_IN_s2[58], ROUND_IN_s1[58], ROUND_IN_s0[58]}), .b ({ROUND_IN_s3[59], ROUND_IN_s2[59], ROUND_IN_s1[59], ROUND_IN_s0[59]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, new_AGEMA_signal_1841, S_7_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_7_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[57], ROUND_IN_s2[57], ROUND_IN_s1[57], ROUND_IN_s0[57]}), .b ({ROUND_IN_s3[58], ROUND_IN_s2[58], ROUND_IN_s1[58], ROUND_IN_s0[58]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1847, S_7_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_8_U6 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, new_AGEMA_signal_1871, S_8_R1[1]}), .b ({ROUND_IN_s3[70], ROUND_IN_s2[70], ROUND_IN_s1[70], ROUND_IN_s0[70]}), .c ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, CONST_ADDITION[66]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_8_U3 ( .a ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, new_AGEMA_signal_1865, S_8_R2[0]}), .b ({ROUND_IN_s3[64], ROUND_IN_s2[64], ROUND_IN_s1[64], ROUND_IN_s0[64]}), .c ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, new_AGEMA_signal_2168, CONST_ADDITION[69]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_8_U2 ( .a ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, new_AGEMA_signal_1856, S_8_R1[0]}), .b ({ROUND_IN_s3[68], ROUND_IN_s2[68], ROUND_IN_s1[68], ROUND_IN_s0[68]}), .c ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, CONST_ADDITION[70]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_8_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[70], ROUND_IN_s2[70], ROUND_IN_s1[70], ROUND_IN_s0[70]}), .b ({ROUND_IN_s3[71], ROUND_IN_s2[71], ROUND_IN_s1[71], ROUND_IN_s0[71]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, new_AGEMA_signal_1856, S_8_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_8_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[66], ROUND_IN_s2[66], ROUND_IN_s1[66], ROUND_IN_s0[66]}), .b ({ROUND_IN_s3[67], ROUND_IN_s2[67], ROUND_IN_s1[67], ROUND_IN_s0[67]}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, new_AGEMA_signal_1865, S_8_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_8_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[65], ROUND_IN_s2[65], ROUND_IN_s1[65], ROUND_IN_s0[65]}), .b ({ROUND_IN_s3[66], ROUND_IN_s2[66], ROUND_IN_s1[66], ROUND_IN_s0[66]}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, new_AGEMA_signal_1871, S_8_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_9_U6 ( .a ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, new_AGEMA_signal_1895, S_9_R1[1]}), .b ({ROUND_IN_s3[78], ROUND_IN_s2[78], ROUND_IN_s1[78], ROUND_IN_s0[78]}), .c ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, CONST_ADDITION[74]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_9_U3 ( .a ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, new_AGEMA_signal_1889, S_9_R2[0]}), .b ({ROUND_IN_s3[72], ROUND_IN_s2[72], ROUND_IN_s1[72], ROUND_IN_s0[72]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, CONST_ADDITION[77]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_9_U2 ( .a ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, new_AGEMA_signal_1880, S_9_R1[0]}), .b ({ROUND_IN_s3[76], ROUND_IN_s2[76], ROUND_IN_s1[76], ROUND_IN_s0[76]}), .c ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, CONST_ADDITION[78]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_9_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[78], ROUND_IN_s2[78], ROUND_IN_s1[78], ROUND_IN_s0[78]}), .b ({ROUND_IN_s3[79], ROUND_IN_s2[79], ROUND_IN_s1[79], ROUND_IN_s0[79]}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, new_AGEMA_signal_1880, S_9_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_9_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[74], ROUND_IN_s2[74], ROUND_IN_s1[74], ROUND_IN_s0[74]}), .b ({ROUND_IN_s3[75], ROUND_IN_s2[75], ROUND_IN_s1[75], ROUND_IN_s0[75]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, new_AGEMA_signal_1889, S_9_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_9_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[73], ROUND_IN_s2[73], ROUND_IN_s1[73], ROUND_IN_s0[73]}), .b ({ROUND_IN_s3[74], ROUND_IN_s2[74], ROUND_IN_s1[74], ROUND_IN_s0[74]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, new_AGEMA_signal_1895, S_9_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_10_U6 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, new_AGEMA_signal_1919, S_10_R1[1]}), .b ({ROUND_IN_s3[86], ROUND_IN_s2[86], ROUND_IN_s1[86], ROUND_IN_s0[86]}), .c ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, new_AGEMA_signal_2192, CONST_ADDITION[82]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_10_U3 ( .a ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, new_AGEMA_signal_1913, S_10_R2[0]}), .b ({ROUND_IN_s3[80], ROUND_IN_s2[80], ROUND_IN_s1[80], ROUND_IN_s0[80]}), .c ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, new_AGEMA_signal_2198, CONST_ADDITION[85]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_10_U2 ( .a ({new_AGEMA_signal_1906, new_AGEMA_signal_1905, new_AGEMA_signal_1904, S_10_R1[0]}), .b ({ROUND_IN_s3[84], ROUND_IN_s2[84], ROUND_IN_s1[84], ROUND_IN_s0[84]}), .c ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, new_AGEMA_signal_2204, CONST_ADDITION[86]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_10_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[86], ROUND_IN_s2[86], ROUND_IN_s1[86], ROUND_IN_s0[86]}), .b ({ROUND_IN_s3[87], ROUND_IN_s2[87], ROUND_IN_s1[87], ROUND_IN_s0[87]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1906, new_AGEMA_signal_1905, new_AGEMA_signal_1904, S_10_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_10_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[82], ROUND_IN_s2[82], ROUND_IN_s1[82], ROUND_IN_s0[82]}), .b ({ROUND_IN_s3[83], ROUND_IN_s2[83], ROUND_IN_s1[83], ROUND_IN_s0[83]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, new_AGEMA_signal_1913, S_10_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_10_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[81], ROUND_IN_s2[81], ROUND_IN_s1[81], ROUND_IN_s0[81]}), .b ({ROUND_IN_s3[82], ROUND_IN_s2[82], ROUND_IN_s1[82], ROUND_IN_s0[82]}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, new_AGEMA_signal_1919, S_10_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_11_U6 ( .a ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, new_AGEMA_signal_1943, S_11_R1[1]}), .b ({ROUND_IN_s3[94], ROUND_IN_s2[94], ROUND_IN_s1[94], ROUND_IN_s0[94]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, new_AGEMA_signal_2207, CONST_ADDITION[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_11_U3 ( .a ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, new_AGEMA_signal_1937, S_11_R2[0]}), .b ({ROUND_IN_s3[88], ROUND_IN_s2[88], ROUND_IN_s1[88], ROUND_IN_s0[88]}), .c ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, new_AGEMA_signal_2213, CONST_ADDITION[93]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_11_U2 ( .a ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, new_AGEMA_signal_1928, S_11_R1[0]}), .b ({ROUND_IN_s3[92], ROUND_IN_s2[92], ROUND_IN_s1[92], ROUND_IN_s0[92]}), .c ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, new_AGEMA_signal_2219, CONST_ADDITION[94]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_11_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[94], ROUND_IN_s2[94], ROUND_IN_s1[94], ROUND_IN_s0[94]}), .b ({ROUND_IN_s3[95], ROUND_IN_s2[95], ROUND_IN_s1[95], ROUND_IN_s0[95]}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, new_AGEMA_signal_1928, S_11_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_11_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[90], ROUND_IN_s2[90], ROUND_IN_s1[90], ROUND_IN_s0[90]}), .b ({ROUND_IN_s3[91], ROUND_IN_s2[91], ROUND_IN_s1[91], ROUND_IN_s0[91]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, new_AGEMA_signal_1937, S_11_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_11_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[89], ROUND_IN_s2[89], ROUND_IN_s1[89], ROUND_IN_s0[89]}), .b ({ROUND_IN_s3[90], ROUND_IN_s2[90], ROUND_IN_s1[90], ROUND_IN_s0[90]}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, new_AGEMA_signal_1943, S_11_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_12_U6 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, new_AGEMA_signal_1967, S_12_R1[1]}), .b ({ROUND_IN_s3[102], ROUND_IN_s2[102], ROUND_IN_s1[102], ROUND_IN_s0[102]}), .c ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, CONST_ADDITION[98]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_12_U3 ( .a ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, new_AGEMA_signal_1961, S_12_R2[0]}), .b ({ROUND_IN_s3[96], ROUND_IN_s2[96], ROUND_IN_s1[96], ROUND_IN_s0[96]}), .c ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, new_AGEMA_signal_2228, CONST_ADDITION[101]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_12_U2 ( .a ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, new_AGEMA_signal_1952, S_12_R1[0]}), .b ({ROUND_IN_s3[100], ROUND_IN_s2[100], ROUND_IN_s1[100], ROUND_IN_s0[100]}), .c ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, CONST_ADDITION[102]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_12_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[102], ROUND_IN_s2[102], ROUND_IN_s1[102], ROUND_IN_s0[102]}), .b ({ROUND_IN_s3[103], ROUND_IN_s2[103], ROUND_IN_s1[103], ROUND_IN_s0[103]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, new_AGEMA_signal_1952, S_12_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_12_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[98], ROUND_IN_s2[98], ROUND_IN_s1[98], ROUND_IN_s0[98]}), .b ({ROUND_IN_s3[99], ROUND_IN_s2[99], ROUND_IN_s1[99], ROUND_IN_s0[99]}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, new_AGEMA_signal_1961, S_12_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_12_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[97], ROUND_IN_s2[97], ROUND_IN_s1[97], ROUND_IN_s0[97]}), .b ({ROUND_IN_s3[98], ROUND_IN_s2[98], ROUND_IN_s1[98], ROUND_IN_s0[98]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, new_AGEMA_signal_1967, S_12_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_13_U6 ( .a ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1991, S_13_R1[1]}), .b ({ROUND_IN_s3[110], ROUND_IN_s2[110], ROUND_IN_s1[110], ROUND_IN_s0[110]}), .c ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, new_AGEMA_signal_2237, CONST_ADDITION[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_13_U3 ( .a ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, S_13_R2[0]}), .b ({ROUND_IN_s3[104], ROUND_IN_s2[104], ROUND_IN_s1[104], ROUND_IN_s0[104]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, CONST_ADDITION[109]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_13_U2 ( .a ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, new_AGEMA_signal_1976, S_13_R1[0]}), .b ({ROUND_IN_s3[108], ROUND_IN_s2[108], ROUND_IN_s1[108], ROUND_IN_s0[108]}), .c ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, new_AGEMA_signal_2249, CONST_ADDITION[110]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_13_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[110], ROUND_IN_s2[110], ROUND_IN_s1[110], ROUND_IN_s0[110]}), .b ({ROUND_IN_s3[111], ROUND_IN_s2[111], ROUND_IN_s1[111], ROUND_IN_s0[111]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, new_AGEMA_signal_1976, S_13_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_13_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[106], ROUND_IN_s2[106], ROUND_IN_s1[106], ROUND_IN_s0[106]}), .b ({ROUND_IN_s3[107], ROUND_IN_s2[107], ROUND_IN_s1[107], ROUND_IN_s0[107]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, new_AGEMA_signal_1985, S_13_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_13_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[105], ROUND_IN_s2[105], ROUND_IN_s1[105], ROUND_IN_s0[105]}), .b ({ROUND_IN_s3[106], ROUND_IN_s2[106], ROUND_IN_s1[106], ROUND_IN_s0[106]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1991, S_13_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_14_U6 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2015, S_14_R1[1]}), .b ({ROUND_IN_s3[118], ROUND_IN_s2[118], ROUND_IN_s1[118], ROUND_IN_s0[118]}), .c ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, new_AGEMA_signal_2252, CONST_ADDITION[114]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_14_U3 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, new_AGEMA_signal_2009, S_14_R2[0]}), .b ({ROUND_IN_s3[112], ROUND_IN_s2[112], ROUND_IN_s1[112], ROUND_IN_s0[112]}), .c ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, CONST_ADDITION[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_14_U2 ( .a ({new_AGEMA_signal_2002, new_AGEMA_signal_2001, new_AGEMA_signal_2000, S_14_R1[0]}), .b ({ROUND_IN_s3[116], ROUND_IN_s2[116], ROUND_IN_s1[116], ROUND_IN_s0[116]}), .c ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, new_AGEMA_signal_2264, CONST_ADDITION[118]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_14_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[118], ROUND_IN_s2[118], ROUND_IN_s1[118], ROUND_IN_s0[118]}), .b ({ROUND_IN_s3[119], ROUND_IN_s2[119], ROUND_IN_s1[119], ROUND_IN_s0[119]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_2002, new_AGEMA_signal_2001, new_AGEMA_signal_2000, S_14_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_14_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[114], ROUND_IN_s2[114], ROUND_IN_s1[114], ROUND_IN_s0[114]}), .b ({ROUND_IN_s3[115], ROUND_IN_s2[115], ROUND_IN_s1[115], ROUND_IN_s0[115]}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, new_AGEMA_signal_2009, S_14_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_14_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[113], ROUND_IN_s2[113], ROUND_IN_s1[113], ROUND_IN_s0[113]}), .b ({ROUND_IN_s3[114], ROUND_IN_s2[114], ROUND_IN_s1[114], ROUND_IN_s0[114]}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2015, S_14_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_15_U6 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, S_15_R1[1]}), .b ({ROUND_IN_s3[126], ROUND_IN_s2[126], ROUND_IN_s1[126], ROUND_IN_s0[126]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, new_AGEMA_signal_2267, SUBSTITUTION[122]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_15_U3 ( .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, S_15_R2[0]}), .b ({ROUND_IN_s3[120], ROUND_IN_s2[120], ROUND_IN_s1[120], ROUND_IN_s0[120]}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, new_AGEMA_signal_2273, CONST_ADDITION[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_15_U2 ( .a ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2024, S_15_R1[0]}), .b ({ROUND_IN_s3[124], ROUND_IN_s2[124], ROUND_IN_s1[124], ROUND_IN_s0[124]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, CONST_ADDITION[126]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_15_NOR1Inst_0_U1 ( .a ({ROUND_IN_s3[126], ROUND_IN_s2[126], ROUND_IN_s1[126], ROUND_IN_s0[126]}), .b ({ROUND_IN_s3[127], ROUND_IN_s2[127], ROUND_IN_s1[127], ROUND_IN_s0[127]}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2024, S_15_R1[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_15_NOR2Inst_0_U1 ( .a ({ROUND_IN_s3[122], ROUND_IN_s2[122], ROUND_IN_s1[122], ROUND_IN_s0[122]}), .b ({ROUND_IN_s3[123], ROUND_IN_s2[123], ROUND_IN_s1[123], ROUND_IN_s0[123]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, S_15_R2[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_15_NOR1Inst_1_U1 ( .a ({ROUND_IN_s3[121], ROUND_IN_s2[121], ROUND_IN_s1[121], ROUND_IN_s0[121]}), .b ({ROUND_IN_s3[122], ROUND_IN_s2[122], ROUND_IN_s1[122], ROUND_IN_s0[122]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, S_15_R1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U92 ( .a ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, SHIFTROWS[30]}), .b ({ROUND_OUT_s3[30], ROUND_OUT_s2[30], ROUND_OUT_s1[30], ROUND_OUT_s0[30]}), .c ({ROUND_OUT_s3[126], ROUND_OUT_s2[126], ROUND_OUT_s1[126], ROUND_OUT_s0[126]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U91 ( .a ({ROUND_OUT_s3[94], ROUND_OUT_s2[94], ROUND_OUT_s1[94], ROUND_OUT_s0[94]}), .b ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, new_AGEMA_signal_2129, SHIFTROWS[62]}), .c ({ROUND_OUT_s3[30], ROUND_OUT_s2[30], ROUND_OUT_s1[30], ROUND_OUT_s0[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U80 ( .a ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, SHIFTROWS[14]}), .b ({ROUND_OUT_s3[14], ROUND_OUT_s2[14], ROUND_OUT_s1[14], ROUND_OUT_s0[14]}), .c ({ROUND_OUT_s3[110], ROUND_OUT_s2[110], ROUND_OUT_s1[110], ROUND_OUT_s0[110]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U79 ( .a ({ROUND_OUT_s3[78], ROUND_OUT_s2[78], ROUND_OUT_s1[78], ROUND_OUT_s0[78]}), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, new_AGEMA_signal_2159, SHIFTROWS[46]}), .c ({ROUND_OUT_s3[14], ROUND_OUT_s2[14], ROUND_OUT_s1[14], ROUND_OUT_s0[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U78 ( .a ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, SHIFTROWS[13]}), .b ({ROUND_OUT_s3[13], ROUND_OUT_s2[13], ROUND_OUT_s1[13], ROUND_OUT_s0[13]}), .c ({ROUND_OUT_s3[109], ROUND_OUT_s2[109], ROUND_OUT_s1[109], ROUND_OUT_s0[109]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U77 ( .a ({ROUND_OUT_s3[77], ROUND_OUT_s2[77], ROUND_OUT_s1[77], ROUND_OUT_s0[77]}), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, SHIFTROWS[45]}), .c ({ROUND_OUT_s3[13], ROUND_OUT_s2[13], ROUND_OUT_s1[13], ROUND_OUT_s0[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U74 ( .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, SHIFTROWS[22]}), .b ({ROUND_OUT_s3[22], ROUND_OUT_s2[22], ROUND_OUT_s1[22], ROUND_OUT_s0[22]}), .c ({ROUND_OUT_s3[118], ROUND_OUT_s2[118], ROUND_OUT_s1[118], ROUND_OUT_s0[118]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U73 ( .a ({ROUND_OUT_s3[86], ROUND_OUT_s2[86], ROUND_OUT_s1[86], ROUND_OUT_s0[86]}), .b ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, new_AGEMA_signal_2114, SHIFTROWS[54]}), .c ({ROUND_OUT_s3[22], ROUND_OUT_s2[22], ROUND_OUT_s1[22], ROUND_OUT_s0[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U68 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, SHIFTROWS[21]}), .b ({ROUND_OUT_s3[21], ROUND_OUT_s2[21], ROUND_OUT_s1[21], ROUND_OUT_s0[21]}), .c ({ROUND_OUT_s3[117], ROUND_OUT_s2[117], ROUND_OUT_s1[117], ROUND_OUT_s0[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U67 ( .a ({ROUND_OUT_s3[85], ROUND_OUT_s2[85], ROUND_OUT_s1[85], ROUND_OUT_s0[85]}), .b ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, SHIFTROWS[53]}), .c ({ROUND_OUT_s3[21], ROUND_OUT_s2[21], ROUND_OUT_s1[21], ROUND_OUT_s0[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U66 ( .a ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, SHIFTROWS[10]}), .b ({ROUND_OUT_s3[10], ROUND_OUT_s2[10], ROUND_OUT_s1[10], ROUND_OUT_s0[10]}), .c ({ROUND_OUT_s3[106], ROUND_OUT_s2[106], ROUND_OUT_s1[106], ROUND_OUT_s0[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U65 ( .a ({ROUND_OUT_s3[74], ROUND_OUT_s2[74], ROUND_OUT_s1[74], ROUND_OUT_s0[74]}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, new_AGEMA_signal_2147, SHIFTROWS[42]}), .c ({ROUND_OUT_s3[10], ROUND_OUT_s2[10], ROUND_OUT_s1[10], ROUND_OUT_s0[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U62 ( .a ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, SHIFTROWS[29]}), .b ({ROUND_OUT_s3[29], ROUND_OUT_s2[29], ROUND_OUT_s1[29], ROUND_OUT_s0[29]}), .c ({ROUND_OUT_s3[125], ROUND_OUT_s2[125], ROUND_OUT_s1[125], ROUND_OUT_s0[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U61 ( .a ({ROUND_OUT_s3[93], ROUND_OUT_s2[93], ROUND_OUT_s1[93], ROUND_OUT_s0[93]}), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, new_AGEMA_signal_2123, SHIFTROWS[61]}), .c ({ROUND_OUT_s3[29], ROUND_OUT_s2[29], ROUND_OUT_s1[29], ROUND_OUT_s0[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U60 ( .a ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, SHIFTROWS[26]}), .b ({ROUND_OUT_s3[26], ROUND_OUT_s2[26], ROUND_OUT_s1[26], ROUND_OUT_s0[26]}), .c ({ROUND_OUT_s3[122], ROUND_OUT_s2[122], ROUND_OUT_s1[122], ROUND_OUT_s0[122]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U59 ( .a ({ROUND_OUT_s3[90], ROUND_OUT_s2[90], ROUND_OUT_s1[90], ROUND_OUT_s0[90]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, new_AGEMA_signal_2117, SHIFTROWS[58]}), .c ({ROUND_OUT_s3[26], ROUND_OUT_s2[26], ROUND_OUT_s1[26], ROUND_OUT_s0[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U50 ( .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, SHIFTROWS[6]}), .b ({ROUND_OUT_s3[6], ROUND_OUT_s2[6], ROUND_OUT_s1[6], ROUND_OUT_s0[6]}), .c ({ROUND_OUT_s3[102], ROUND_OUT_s2[102], ROUND_OUT_s1[102], ROUND_OUT_s0[102]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U49 ( .a ({ROUND_OUT_s3[70], ROUND_OUT_s2[70], ROUND_OUT_s1[70], ROUND_OUT_s0[70]}), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, SHIFTROWS[38]}), .c ({ROUND_OUT_s3[6], ROUND_OUT_s2[6], ROUND_OUT_s1[6], ROUND_OUT_s0[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U48 ( .a ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, SHIFTROWS[5]}), .b ({ROUND_OUT_s3[5], ROUND_OUT_s2[5], ROUND_OUT_s1[5], ROUND_OUT_s0[5]}), .c ({ROUND_OUT_s3[101], ROUND_OUT_s2[101], ROUND_OUT_s1[101], ROUND_OUT_s0[101]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U47 ( .a ({ROUND_OUT_s3[69], ROUND_OUT_s2[69], ROUND_OUT_s1[69], ROUND_OUT_s0[69]}), .b ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, new_AGEMA_signal_2138, SHIFTROWS[37]}), .c ({ROUND_OUT_s3[5], ROUND_OUT_s2[5], ROUND_OUT_s1[5], ROUND_OUT_s0[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U44 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, new_AGEMA_signal_2057, SHIFTROWS[18]}), .b ({ROUND_OUT_s3[18], ROUND_OUT_s2[18], ROUND_OUT_s1[18], ROUND_OUT_s0[18]}), .c ({ROUND_OUT_s3[114], ROUND_OUT_s2[114], ROUND_OUT_s1[114], ROUND_OUT_s0[114]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U43 ( .a ({ROUND_OUT_s3[82], ROUND_OUT_s2[82], ROUND_OUT_s1[82], ROUND_OUT_s0[82]}), .b ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, SHIFTROWS[50]}), .c ({ROUND_OUT_s3[18], ROUND_OUT_s2[18], ROUND_OUT_s1[18], ROUND_OUT_s0[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U36 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, SHIFTROWS[2]}), .b ({ROUND_OUT_s3[2], ROUND_OUT_s2[2], ROUND_OUT_s1[2], ROUND_OUT_s0[2]}), .c ({ROUND_OUT_s3[98], ROUND_OUT_s2[98], ROUND_OUT_s1[98], ROUND_OUT_s0[98]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U35 ( .a ({ROUND_OUT_s3[66], ROUND_OUT_s2[66], ROUND_OUT_s1[66], ROUND_OUT_s0[66]}), .b ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, new_AGEMA_signal_2132, SHIFTROWS[34]}), .c ({ROUND_OUT_s3[2], ROUND_OUT_s2[2], ROUND_OUT_s1[2], ROUND_OUT_s0[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U30 ( .a ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, new_AGEMA_signal_2132, SHIFTROWS[34]}), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, new_AGEMA_signal_2549, SHIFTROWS[66]}), .c ({ROUND_OUT_s3[34], ROUND_OUT_s2[34], ROUND_OUT_s1[34], ROUND_OUT_s0[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U27 ( .a ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, new_AGEMA_signal_2138, SHIFTROWS[37]}), .b ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, new_AGEMA_signal_2546, SHIFTROWS[69]}), .c ({ROUND_OUT_s3[37], ROUND_OUT_s2[37], ROUND_OUT_s1[37], ROUND_OUT_s0[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U26 ( .a ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, SHIFTROWS[38]}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, new_AGEMA_signal_2543, SHIFTROWS[70]}), .c ({ROUND_OUT_s3[38], ROUND_OUT_s2[38], ROUND_OUT_s1[38], ROUND_OUT_s0[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U22 ( .a ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, new_AGEMA_signal_2147, SHIFTROWS[42]}), .b ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, new_AGEMA_signal_2540, SHIFTROWS[74]}), .c ({ROUND_OUT_s3[42], ROUND_OUT_s2[42], ROUND_OUT_s1[42], ROUND_OUT_s0[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U19 ( .a ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, SHIFTROWS[45]}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, new_AGEMA_signal_2537, SHIFTROWS[77]}), .c ({ROUND_OUT_s3[45], ROUND_OUT_s2[45], ROUND_OUT_s1[45], ROUND_OUT_s0[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U18 ( .a ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, new_AGEMA_signal_2159, SHIFTROWS[46]}), .b ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, new_AGEMA_signal_2534, SHIFTROWS[78]}), .c ({ROUND_OUT_s3[46], ROUND_OUT_s2[46], ROUND_OUT_s1[46], ROUND_OUT_s0[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U14 ( .a ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, SHIFTROWS[50]}), .b ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, new_AGEMA_signal_2531, SHIFTROWS[82]}), .c ({ROUND_OUT_s3[50], ROUND_OUT_s2[50], ROUND_OUT_s1[50], ROUND_OUT_s0[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U11 ( .a ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, SHIFTROWS[53]}), .b ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, new_AGEMA_signal_2528, SHIFTROWS[85]}), .c ({ROUND_OUT_s3[53], ROUND_OUT_s2[53], ROUND_OUT_s1[53], ROUND_OUT_s0[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U10 ( .a ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, new_AGEMA_signal_2114, SHIFTROWS[54]}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, new_AGEMA_signal_2525, SHIFTROWS[86]}), .c ({ROUND_OUT_s3[54], ROUND_OUT_s2[54], ROUND_OUT_s1[54], ROUND_OUT_s0[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U6 ( .a ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, new_AGEMA_signal_2117, SHIFTROWS[58]}), .b ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, new_AGEMA_signal_2558, SHIFTROWS[90]}), .c ({ROUND_OUT_s3[58], ROUND_OUT_s2[58], ROUND_OUT_s1[58], ROUND_OUT_s0[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U3 ( .a ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, new_AGEMA_signal_2123, SHIFTROWS[61]}), .b ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, new_AGEMA_signal_2555, SHIFTROWS[93]}), .c ({ROUND_OUT_s3[61], ROUND_OUT_s2[61], ROUND_OUT_s1[61], ROUND_OUT_s0[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U2 ( .a ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, new_AGEMA_signal_2129, SHIFTROWS[62]}), .b ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, new_AGEMA_signal_2552, SHIFTROWS[94]}), .c ({ROUND_OUT_s3[62], ROUND_OUT_s2[62], ROUND_OUT_s1[62], ROUND_OUT_s0[62]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U401 ( .a ({ROUND_KEY_s3[355], ROUND_KEY_s2[355], ROUND_KEY_s1[355], ROUND_KEY_s0[355]}), .b ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, CONST_ADDITION[99]}), .c ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, new_AGEMA_signal_2741, n405}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U402 ( .a ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, new_AGEMA_signal_1088, n406}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, new_AGEMA_signal_2741, n405}), .c ({ROUND_OUT_s3[67], ROUND_OUT_s2[67], ROUND_OUT_s1[67], ROUND_OUT_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U413 ( .a ({ROUND_KEY_s3[351], ROUND_KEY_s2[351], ROUND_KEY_s1[351], ROUND_KEY_s0[351]}), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, CONST_ADDITION[95]}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, new_AGEMA_signal_2747, n413}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U414 ( .a ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, new_AGEMA_signal_1124, n414}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, new_AGEMA_signal_2747, n413}), .c ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, new_AGEMA_signal_3005, SHIFTROWS[87]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U425 ( .a ({ROUND_KEY_s3[347], ROUND_KEY_s2[347], ROUND_KEY_s1[347], ROUND_KEY_s0[347]}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, CONST_ADDITION[91]}), .c ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, new_AGEMA_signal_2753, n421}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U426 ( .a ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, new_AGEMA_signal_1160, n422}), .b ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, new_AGEMA_signal_2753, n421}), .c ({new_AGEMA_signal_3010, new_AGEMA_signal_3009, new_AGEMA_signal_3008, SHIFTROWS[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U439 ( .a ({ROUND_KEY_s3[343], ROUND_KEY_s2[343], ROUND_KEY_s1[343], ROUND_KEY_s0[343]}), .b ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, CONST_ADDITION[87]}), .c ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, new_AGEMA_signal_2759, n431}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U440 ( .a ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, new_AGEMA_signal_1196, n432}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, new_AGEMA_signal_2759, n431}), .c ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, new_AGEMA_signal_3011, SHIFTROWS[79]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U451 ( .a ({ROUND_KEY_s3[339], ROUND_KEY_s2[339], ROUND_KEY_s1[339], ROUND_KEY_s0[339]}), .b ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, CONST_ADDITION[83]}), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, new_AGEMA_signal_2765, n439}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U452 ( .a ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, new_AGEMA_signal_1232, n440}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, new_AGEMA_signal_2765, n439}), .c ({new_AGEMA_signal_3016, new_AGEMA_signal_3015, new_AGEMA_signal_3014, SHIFTROWS[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U463 ( .a ({ROUND_KEY_s3[335], ROUND_KEY_s2[335], ROUND_KEY_s1[335], ROUND_KEY_s0[335]}), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, new_AGEMA_signal_2681, CONST_ADDITION[79]}), .c ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2771, n447}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U464 ( .a ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, new_AGEMA_signal_1268, n448}), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2771, n447}), .c ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, new_AGEMA_signal_3017, SHIFTROWS[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U475 ( .a ({ROUND_KEY_s3[331], ROUND_KEY_s2[331], ROUND_KEY_s1[331], ROUND_KEY_s0[331]}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, CONST_ADDITION[75]}), .c ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, new_AGEMA_signal_2777, n455}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U476 ( .a ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, new_AGEMA_signal_1304, n456}), .b ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, new_AGEMA_signal_2777, n455}), .c ({new_AGEMA_signal_3022, new_AGEMA_signal_3021, new_AGEMA_signal_3020, SHIFTROWS[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U487 ( .a ({ROUND_KEY_s3[327], ROUND_KEY_s2[327], ROUND_KEY_s1[327], ROUND_KEY_s0[327]}), .b ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, new_AGEMA_signal_2672, CONST_ADDITION[71]}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, new_AGEMA_signal_2783, n463}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U488 ( .a ({new_AGEMA_signal_1342, new_AGEMA_signal_1341, new_AGEMA_signal_1340, n464}), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, new_AGEMA_signal_2783, n463}), .c ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, new_AGEMA_signal_3023, SHIFTROWS[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U499 ( .a ({ROUND_KEY_s3[323], ROUND_KEY_s2[323], ROUND_KEY_s1[323], ROUND_KEY_s0[323]}), .b ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, new_AGEMA_signal_2666, CONST_ADDITION[67]}), .c ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, new_AGEMA_signal_2789, n471}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U500 ( .a ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, new_AGEMA_signal_1376, n472}), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, new_AGEMA_signal_2789, n471}), .c ({new_AGEMA_signal_3028, new_AGEMA_signal_3027, new_AGEMA_signal_3026, SHIFTROWS[91]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U511 ( .a ({ROUND_KEY_s3[383], ROUND_KEY_s2[383], ROUND_KEY_s1[383], ROUND_KEY_s0[383]}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, new_AGEMA_signal_2735, CONST_ADDITION[127]}), .c ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, new_AGEMA_signal_2795, n479}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U512 ( .a ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, new_AGEMA_signal_1412, n480}), .b ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, new_AGEMA_signal_2795, n479}), .c ({ROUND_OUT_s3[95], ROUND_OUT_s2[95], ROUND_OUT_s1[95], ROUND_OUT_s0[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U523 ( .a ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, new_AGEMA_signal_2729, SUBSTITUTION[123]}), .b ({ROUND_KEY_s3[379], ROUND_KEY_s2[379], ROUND_KEY_s1[379], ROUND_KEY_s0[379]}), .c ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, new_AGEMA_signal_2801, n487}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U524 ( .a ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, new_AGEMA_signal_1448, n488}), .b ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, new_AGEMA_signal_2801, n487}), .c ({new_AGEMA_signal_3034, new_AGEMA_signal_3033, new_AGEMA_signal_3032, n489}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U525 ( .a ({1'b0, 1'b0, 1'b0, CONST_IN[3]}), .b ({new_AGEMA_signal_3034, new_AGEMA_signal_3033, new_AGEMA_signal_3032, n489}), .c ({ROUND_OUT_s3[91], ROUND_OUT_s2[91], ROUND_OUT_s1[91], ROUND_OUT_s0[91]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U539 ( .a ({ROUND_KEY_s3[375], ROUND_KEY_s2[375], ROUND_KEY_s1[375], ROUND_KEY_s0[375]}), .b ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, CONST_ADDITION[119]}), .c ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810, n499}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U540 ( .a ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, new_AGEMA_signal_1484, n500}), .b ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810, n499}), .c ({ROUND_OUT_s3[87], ROUND_OUT_s2[87], ROUND_OUT_s1[87], ROUND_OUT_s0[87]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U551 ( .a ({ROUND_KEY_s3[371], ROUND_KEY_s2[371], ROUND_KEY_s1[371], ROUND_KEY_s0[371]}), .b ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, CONST_ADDITION[115]}), .c ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, new_AGEMA_signal_2816, n507}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U552 ( .a ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, new_AGEMA_signal_1520, n508}), .b ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, new_AGEMA_signal_2816, n507}), .c ({ROUND_OUT_s3[83], ROUND_OUT_s2[83], ROUND_OUT_s1[83], ROUND_OUT_s0[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U563 ( .a ({ROUND_KEY_s3[367], ROUND_KEY_s2[367], ROUND_KEY_s1[367], ROUND_KEY_s0[367]}), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, new_AGEMA_signal_2717, CONST_ADDITION[111]}), .c ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, new_AGEMA_signal_2822, n515}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U564 ( .a ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, new_AGEMA_signal_1556, n516}), .b ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, new_AGEMA_signal_2822, n515}), .c ({ROUND_OUT_s3[79], ROUND_OUT_s2[79], ROUND_OUT_s1[79], ROUND_OUT_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U575 ( .a ({ROUND_KEY_s3[363], ROUND_KEY_s2[363], ROUND_KEY_s1[363], ROUND_KEY_s0[363]}), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, CONST_ADDITION[107]}), .c ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, new_AGEMA_signal_2828, n523}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U576 ( .a ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, new_AGEMA_signal_1592, n524}), .b ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, new_AGEMA_signal_2828, n523}), .c ({ROUND_OUT_s3[75], ROUND_OUT_s2[75], ROUND_OUT_s1[75], ROUND_OUT_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U587 ( .a ({ROUND_KEY_s3[359], ROUND_KEY_s2[359], ROUND_KEY_s1[359], ROUND_KEY_s0[359]}), .b ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, CONST_ADDITION[103]}), .c ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, new_AGEMA_signal_2834, n531}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U588 ( .a ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, new_AGEMA_signal_1628, n532}), .b ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, new_AGEMA_signal_2834, n531}), .c ({ROUND_OUT_s3[71], ROUND_OUT_s2[71], ROUND_OUT_s1[71], ROUND_OUT_s0[71]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_0_U5 ( .a ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, new_AGEMA_signal_2429, S_0_R1[2]}), .b ({ROUND_IN_s3[1], ROUND_IN_s2[1], ROUND_IN_s1[1], ROUND_IN_s0[1]}), .c ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, new_AGEMA_signal_2594, SHIFTROWS[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_0_U1 ( .a ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, S_0_R2[1]}), .b ({ROUND_IN_s3[5], ROUND_IN_s2[5], ROUND_IN_s1[5], ROUND_IN_s0[5]}), .c ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, new_AGEMA_signal_2600, SHIFTROWS[15]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_0_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, SHIFTROWS[13]}), .b ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, SHIFTROWS[14]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, S_0_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_0_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[3], ROUND_IN_s2[3], ROUND_IN_s1[3], ROUND_IN_s0[3]}), .b ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, SHIFTROWS[13]}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, new_AGEMA_signal_2429, S_0_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_1_U5 ( .a ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, new_AGEMA_signal_2435, S_1_R1[2]}), .b ({ROUND_IN_s3[9], ROUND_IN_s2[9], ROUND_IN_s1[9], ROUND_IN_s0[9]}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, new_AGEMA_signal_2603, SHIFTROWS[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_1_U1 ( .a ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, new_AGEMA_signal_2432, S_1_R2[1]}), .b ({ROUND_IN_s3[13], ROUND_IN_s2[13], ROUND_IN_s1[13], ROUND_IN_s0[13]}), .c ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, new_AGEMA_signal_2609, SHIFTROWS[23]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_1_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, SHIFTROWS[21]}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, SHIFTROWS[22]}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, new_AGEMA_signal_2432, S_1_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_1_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[11], ROUND_IN_s2[11], ROUND_IN_s1[11], ROUND_IN_s0[11]}), .b ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, SHIFTROWS[21]}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, new_AGEMA_signal_2435, S_1_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_2_U5 ( .a ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, new_AGEMA_signal_2441, S_2_R1[2]}), .b ({ROUND_IN_s3[17], ROUND_IN_s2[17], ROUND_IN_s1[17], ROUND_IN_s0[17]}), .c ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, new_AGEMA_signal_2612, SHIFTROWS[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_2_U1 ( .a ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, new_AGEMA_signal_2438, S_2_R2[1]}), .b ({ROUND_IN_s3[21], ROUND_IN_s2[21], ROUND_IN_s1[21], ROUND_IN_s0[21]}), .c ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, new_AGEMA_signal_2618, SHIFTROWS[31]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_2_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, SHIFTROWS[29]}), .b ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, SHIFTROWS[30]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, new_AGEMA_signal_2438, S_2_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_2_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[19], ROUND_IN_s2[19], ROUND_IN_s1[19], ROUND_IN_s0[19]}), .b ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, SHIFTROWS[29]}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, new_AGEMA_signal_2441, S_2_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_3_U5 ( .a ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, new_AGEMA_signal_2447, S_3_R1[2]}), .b ({ROUND_IN_s3[25], ROUND_IN_s2[25], ROUND_IN_s1[25], ROUND_IN_s0[25]}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, new_AGEMA_signal_2621, SHIFTROWS[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_3_U1 ( .a ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, new_AGEMA_signal_2444, S_3_R2[1]}), .b ({ROUND_IN_s3[29], ROUND_IN_s2[29], ROUND_IN_s1[29], ROUND_IN_s0[29]}), .c ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, new_AGEMA_signal_2627, SHIFTROWS[7]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_3_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, SHIFTROWS[5]}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, SHIFTROWS[6]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, new_AGEMA_signal_2444, S_3_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_3_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[27], ROUND_IN_s2[27], ROUND_IN_s1[27], ROUND_IN_s0[27]}), .b ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, SHIFTROWS[5]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, new_AGEMA_signal_2447, S_3_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_4_U5 ( .a ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, new_AGEMA_signal_2453, S_4_R1[2]}), .b ({ROUND_IN_s3[33], ROUND_IN_s2[33], ROUND_IN_s1[33], ROUND_IN_s0[33]}), .c ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, new_AGEMA_signal_2630, SHIFTROWS[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_4_U1 ( .a ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, new_AGEMA_signal_2450, S_4_R2[1]}), .b ({ROUND_IN_s3[37], ROUND_IN_s2[37], ROUND_IN_s1[37], ROUND_IN_s0[37]}), .c ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, new_AGEMA_signal_2636, SHIFTROWS[55]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_4_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, SHIFTROWS[53]}), .b ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, new_AGEMA_signal_2114, SHIFTROWS[54]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, new_AGEMA_signal_2450, S_4_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_4_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[35], ROUND_IN_s2[35], ROUND_IN_s1[35], ROUND_IN_s0[35]}), .b ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, SHIFTROWS[53]}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, new_AGEMA_signal_2453, S_4_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_5_U5 ( .a ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, new_AGEMA_signal_2459, S_5_R1[2]}), .b ({ROUND_IN_s3[41], ROUND_IN_s2[41], ROUND_IN_s1[41], ROUND_IN_s0[41]}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, SHIFTROWS[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_5_U1 ( .a ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, new_AGEMA_signal_2456, S_5_R2[1]}), .b ({ROUND_IN_s3[45], ROUND_IN_s2[45], ROUND_IN_s1[45], ROUND_IN_s0[45]}), .c ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, new_AGEMA_signal_2645, SHIFTROWS[63]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_5_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, new_AGEMA_signal_2123, SHIFTROWS[61]}), .b ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, new_AGEMA_signal_2129, SHIFTROWS[62]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, new_AGEMA_signal_2456, S_5_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_5_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[43], ROUND_IN_s2[43], ROUND_IN_s1[43], ROUND_IN_s0[43]}), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, new_AGEMA_signal_2123, SHIFTROWS[61]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, new_AGEMA_signal_2459, S_5_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_6_U5 ( .a ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, new_AGEMA_signal_2465, S_6_R1[2]}), .b ({ROUND_IN_s3[49], ROUND_IN_s2[49], ROUND_IN_s1[49], ROUND_IN_s0[49]}), .c ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, new_AGEMA_signal_2648, SHIFTROWS[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_6_U1 ( .a ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, new_AGEMA_signal_2462, S_6_R2[1]}), .b ({ROUND_IN_s3[53], ROUND_IN_s2[53], ROUND_IN_s1[53], ROUND_IN_s0[53]}), .c ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, new_AGEMA_signal_2654, SHIFTROWS[39]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_6_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, new_AGEMA_signal_2138, SHIFTROWS[37]}), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, SHIFTROWS[38]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, new_AGEMA_signal_2462, S_6_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_6_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[51], ROUND_IN_s2[51], ROUND_IN_s1[51], ROUND_IN_s0[51]}), .b ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, new_AGEMA_signal_2138, SHIFTROWS[37]}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, new_AGEMA_signal_2465, S_6_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_7_U5 ( .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, S_7_R1[2]}), .b ({ROUND_IN_s3[57], ROUND_IN_s2[57], ROUND_IN_s1[57], ROUND_IN_s0[57]}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, new_AGEMA_signal_2657, SHIFTROWS[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_7_U1 ( .a ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, new_AGEMA_signal_2468, S_7_R2[1]}), .b ({ROUND_IN_s3[61], ROUND_IN_s2[61], ROUND_IN_s1[61], ROUND_IN_s0[61]}), .c ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, new_AGEMA_signal_2663, SHIFTROWS[47]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_7_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, SHIFTROWS[45]}), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, new_AGEMA_signal_2159, SHIFTROWS[46]}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, new_AGEMA_signal_2468, S_7_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_7_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[59], ROUND_IN_s2[59], ROUND_IN_s1[59], ROUND_IN_s0[59]}), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, SHIFTROWS[45]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, S_7_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_8_U5 ( .a ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, new_AGEMA_signal_2477, S_8_R1[2]}), .b ({ROUND_IN_s3[65], ROUND_IN_s2[65], ROUND_IN_s1[65], ROUND_IN_s0[65]}), .c ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, new_AGEMA_signal_2666, CONST_ADDITION[67]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_8_U1 ( .a ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, new_AGEMA_signal_2474, S_8_R2[1]}), .b ({ROUND_IN_s3[69], ROUND_IN_s2[69], ROUND_IN_s1[69], ROUND_IN_s0[69]}), .c ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, new_AGEMA_signal_2672, CONST_ADDITION[71]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_8_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, new_AGEMA_signal_2168, CONST_ADDITION[69]}), .b ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, CONST_ADDITION[70]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, new_AGEMA_signal_2474, S_8_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_8_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[67], ROUND_IN_s2[67], ROUND_IN_s1[67], ROUND_IN_s0[67]}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, new_AGEMA_signal_2168, CONST_ADDITION[69]}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, new_AGEMA_signal_2477, S_8_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_9_U5 ( .a ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, new_AGEMA_signal_2483, S_9_R1[2]}), .b ({ROUND_IN_s3[73], ROUND_IN_s2[73], ROUND_IN_s1[73], ROUND_IN_s0[73]}), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, CONST_ADDITION[75]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_9_U1 ( .a ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, new_AGEMA_signal_2480, S_9_R2[1]}), .b ({ROUND_IN_s3[77], ROUND_IN_s2[77], ROUND_IN_s1[77], ROUND_IN_s0[77]}), .c ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, new_AGEMA_signal_2681, CONST_ADDITION[79]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_9_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, CONST_ADDITION[77]}), .b ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, CONST_ADDITION[78]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, new_AGEMA_signal_2480, S_9_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_9_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[75], ROUND_IN_s2[75], ROUND_IN_s1[75], ROUND_IN_s0[75]}), .b ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, CONST_ADDITION[77]}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, new_AGEMA_signal_2483, S_9_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_10_U5 ( .a ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, new_AGEMA_signal_2489, S_10_R1[2]}), .b ({ROUND_IN_s3[81], ROUND_IN_s2[81], ROUND_IN_s1[81], ROUND_IN_s0[81]}), .c ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, CONST_ADDITION[83]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_10_U1 ( .a ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, new_AGEMA_signal_2486, S_10_R2[1]}), .b ({ROUND_IN_s3[85], ROUND_IN_s2[85], ROUND_IN_s1[85], ROUND_IN_s0[85]}), .c ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, CONST_ADDITION[87]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_10_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, new_AGEMA_signal_2198, CONST_ADDITION[85]}), .b ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, new_AGEMA_signal_2204, CONST_ADDITION[86]}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, new_AGEMA_signal_2486, S_10_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_10_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[83], ROUND_IN_s2[83], ROUND_IN_s1[83], ROUND_IN_s0[83]}), .b ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, new_AGEMA_signal_2198, CONST_ADDITION[85]}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, new_AGEMA_signal_2489, S_10_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_11_U5 ( .a ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, new_AGEMA_signal_2495, S_11_R1[2]}), .b ({ROUND_IN_s3[89], ROUND_IN_s2[89], ROUND_IN_s1[89], ROUND_IN_s0[89]}), .c ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, CONST_ADDITION[91]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_11_U1 ( .a ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, new_AGEMA_signal_2492, S_11_R2[1]}), .b ({ROUND_IN_s3[93], ROUND_IN_s2[93], ROUND_IN_s1[93], ROUND_IN_s0[93]}), .c ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, CONST_ADDITION[95]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_11_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, new_AGEMA_signal_2213, CONST_ADDITION[93]}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, new_AGEMA_signal_2219, CONST_ADDITION[94]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, new_AGEMA_signal_2492, S_11_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_11_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[91], ROUND_IN_s2[91], ROUND_IN_s1[91], ROUND_IN_s0[91]}), .b ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, new_AGEMA_signal_2213, CONST_ADDITION[93]}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, new_AGEMA_signal_2495, S_11_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_12_U5 ( .a ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, new_AGEMA_signal_2501, S_12_R1[2]}), .b ({ROUND_IN_s3[97], ROUND_IN_s2[97], ROUND_IN_s1[97], ROUND_IN_s0[97]}), .c ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, CONST_ADDITION[99]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_12_U1 ( .a ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, new_AGEMA_signal_2498, S_12_R2[1]}), .b ({ROUND_IN_s3[101], ROUND_IN_s2[101], ROUND_IN_s1[101], ROUND_IN_s0[101]}), .c ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, CONST_ADDITION[103]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_12_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, new_AGEMA_signal_2228, CONST_ADDITION[101]}), .b ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, CONST_ADDITION[102]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, new_AGEMA_signal_2498, S_12_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_12_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[99], ROUND_IN_s2[99], ROUND_IN_s1[99], ROUND_IN_s0[99]}), .b ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, new_AGEMA_signal_2228, CONST_ADDITION[101]}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, new_AGEMA_signal_2501, S_12_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_13_U5 ( .a ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, new_AGEMA_signal_2507, S_13_R1[2]}), .b ({ROUND_IN_s3[105], ROUND_IN_s2[105], ROUND_IN_s1[105], ROUND_IN_s0[105]}), .c ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, CONST_ADDITION[107]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_13_U1 ( .a ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, new_AGEMA_signal_2504, S_13_R2[1]}), .b ({ROUND_IN_s3[109], ROUND_IN_s2[109], ROUND_IN_s1[109], ROUND_IN_s0[109]}), .c ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, new_AGEMA_signal_2717, CONST_ADDITION[111]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_13_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, CONST_ADDITION[109]}), .b ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, new_AGEMA_signal_2249, CONST_ADDITION[110]}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, new_AGEMA_signal_2504, S_13_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_13_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[107], ROUND_IN_s2[107], ROUND_IN_s1[107], ROUND_IN_s0[107]}), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, CONST_ADDITION[109]}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, new_AGEMA_signal_2507, S_13_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_14_U5 ( .a ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, new_AGEMA_signal_2513, S_14_R1[2]}), .b ({ROUND_IN_s3[113], ROUND_IN_s2[113], ROUND_IN_s1[113], ROUND_IN_s0[113]}), .c ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, CONST_ADDITION[115]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_14_U1 ( .a ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, new_AGEMA_signal_2510, S_14_R2[1]}), .b ({ROUND_IN_s3[117], ROUND_IN_s2[117], ROUND_IN_s1[117], ROUND_IN_s0[117]}), .c ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, CONST_ADDITION[119]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_14_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, CONST_ADDITION[117]}), .b ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, new_AGEMA_signal_2264, CONST_ADDITION[118]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, new_AGEMA_signal_2510, S_14_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_14_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[115], ROUND_IN_s2[115], ROUND_IN_s1[115], ROUND_IN_s0[115]}), .b ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, CONST_ADDITION[117]}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, new_AGEMA_signal_2513, S_14_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_15_U5 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, new_AGEMA_signal_2519, S_15_R1[2]}), .b ({ROUND_IN_s3[121], ROUND_IN_s2[121], ROUND_IN_s1[121], ROUND_IN_s0[121]}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, new_AGEMA_signal_2729, SUBSTITUTION[123]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_15_U1 ( .a ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, new_AGEMA_signal_2516, S_15_R2[1]}), .b ({ROUND_IN_s3[125], ROUND_IN_s2[125], ROUND_IN_s1[125], ROUND_IN_s0[125]}), .c ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, new_AGEMA_signal_2735, CONST_ADDITION[127]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_15_NOR2Inst_1_U1 ( .a ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, new_AGEMA_signal_2273, CONST_ADDITION[125]}), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, CONST_ADDITION[126]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, new_AGEMA_signal_2516, S_15_R2[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_15_NOR1Inst_2_U1 ( .a ({ROUND_IN_s3[123], ROUND_IN_s2[123], ROUND_IN_s1[123], ROUND_IN_s0[123]}), .b ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, new_AGEMA_signal_2273, CONST_ADDITION[125]}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, new_AGEMA_signal_2519, S_15_R1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U96 ( .a ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, new_AGEMA_signal_2618, SHIFTROWS[31]}), .b ({ROUND_OUT_s3[31], ROUND_OUT_s2[31], ROUND_OUT_s1[31], ROUND_OUT_s0[31]}), .c ({ROUND_OUT_s3[127], ROUND_OUT_s2[127], ROUND_OUT_s1[127], ROUND_OUT_s0[127]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U95 ( .a ({ROUND_OUT_s3[95], ROUND_OUT_s2[95], ROUND_OUT_s1[95], ROUND_OUT_s0[95]}), .b ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, new_AGEMA_signal_2645, SHIFTROWS[63]}), .c ({ROUND_OUT_s3[31], ROUND_OUT_s2[31], ROUND_OUT_s1[31], ROUND_OUT_s0[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U84 ( .a ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, new_AGEMA_signal_2600, SHIFTROWS[15]}), .b ({ROUND_OUT_s3[15], ROUND_OUT_s2[15], ROUND_OUT_s1[15], ROUND_OUT_s0[15]}), .c ({ROUND_OUT_s3[111], ROUND_OUT_s2[111], ROUND_OUT_s1[111], ROUND_OUT_s0[111]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U83 ( .a ({ROUND_OUT_s3[79], ROUND_OUT_s2[79], ROUND_OUT_s1[79], ROUND_OUT_s0[79]}), .b ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, new_AGEMA_signal_2663, SHIFTROWS[47]}), .c ({ROUND_OUT_s3[15], ROUND_OUT_s2[15], ROUND_OUT_s1[15], ROUND_OUT_s0[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U82 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, new_AGEMA_signal_2609, SHIFTROWS[23]}), .b ({ROUND_OUT_s3[23], ROUND_OUT_s2[23], ROUND_OUT_s1[23], ROUND_OUT_s0[23]}), .c ({ROUND_OUT_s3[119], ROUND_OUT_s2[119], ROUND_OUT_s1[119], ROUND_OUT_s0[119]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U81 ( .a ({ROUND_OUT_s3[87], ROUND_OUT_s2[87], ROUND_OUT_s1[87], ROUND_OUT_s0[87]}), .b ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, new_AGEMA_signal_2636, SHIFTROWS[55]}), .c ({ROUND_OUT_s3[23], ROUND_OUT_s2[23], ROUND_OUT_s1[23], ROUND_OUT_s0[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U76 ( .a ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, new_AGEMA_signal_2612, SHIFTROWS[27]}), .b ({ROUND_OUT_s3[27], ROUND_OUT_s2[27], ROUND_OUT_s1[27], ROUND_OUT_s0[27]}), .c ({ROUND_OUT_s3[123], ROUND_OUT_s2[123], ROUND_OUT_s1[123], ROUND_OUT_s0[123]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U75 ( .a ({ROUND_OUT_s3[91], ROUND_OUT_s2[91], ROUND_OUT_s1[91], ROUND_OUT_s0[91]}), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, SHIFTROWS[59]}), .c ({ROUND_OUT_s3[27], ROUND_OUT_s2[27], ROUND_OUT_s1[27], ROUND_OUT_s0[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U70 ( .a ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, new_AGEMA_signal_2594, SHIFTROWS[11]}), .b ({ROUND_OUT_s3[11], ROUND_OUT_s2[11], ROUND_OUT_s1[11], ROUND_OUT_s0[11]}), .c ({ROUND_OUT_s3[107], ROUND_OUT_s2[107], ROUND_OUT_s1[107], ROUND_OUT_s0[107]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U69 ( .a ({ROUND_OUT_s3[75], ROUND_OUT_s2[75], ROUND_OUT_s1[75], ROUND_OUT_s0[75]}), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, new_AGEMA_signal_2657, SHIFTROWS[43]}), .c ({ROUND_OUT_s3[11], ROUND_OUT_s2[11], ROUND_OUT_s1[11], ROUND_OUT_s0[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U54 ( .a ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, new_AGEMA_signal_2627, SHIFTROWS[7]}), .b ({ROUND_OUT_s3[7], ROUND_OUT_s2[7], ROUND_OUT_s1[7], ROUND_OUT_s0[7]}), .c ({ROUND_OUT_s3[103], ROUND_OUT_s2[103], ROUND_OUT_s1[103], ROUND_OUT_s0[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U53 ( .a ({ROUND_OUT_s3[71], ROUND_OUT_s2[71], ROUND_OUT_s1[71], ROUND_OUT_s0[71]}), .b ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, new_AGEMA_signal_2654, SHIFTROWS[39]}), .c ({ROUND_OUT_s3[7], ROUND_OUT_s2[7], ROUND_OUT_s1[7], ROUND_OUT_s0[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U52 ( .a ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, new_AGEMA_signal_2603, SHIFTROWS[19]}), .b ({ROUND_OUT_s3[19], ROUND_OUT_s2[19], ROUND_OUT_s1[19], ROUND_OUT_s0[19]}), .c ({ROUND_OUT_s3[115], ROUND_OUT_s2[115], ROUND_OUT_s1[115], ROUND_OUT_s0[115]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U51 ( .a ({ROUND_OUT_s3[83], ROUND_OUT_s2[83], ROUND_OUT_s1[83], ROUND_OUT_s0[83]}), .b ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, new_AGEMA_signal_2630, SHIFTROWS[51]}), .c ({ROUND_OUT_s3[19], ROUND_OUT_s2[19], ROUND_OUT_s1[19], ROUND_OUT_s0[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U40 ( .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, new_AGEMA_signal_2621, SHIFTROWS[3]}), .b ({ROUND_OUT_s3[3], ROUND_OUT_s2[3], ROUND_OUT_s1[3], ROUND_OUT_s0[3]}), .c ({ROUND_OUT_s3[99], ROUND_OUT_s2[99], ROUND_OUT_s1[99], ROUND_OUT_s0[99]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U39 ( .a ({ROUND_OUT_s3[67], ROUND_OUT_s2[67], ROUND_OUT_s1[67], ROUND_OUT_s0[67]}), .b ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, new_AGEMA_signal_2648, SHIFTROWS[35]}), .c ({ROUND_OUT_s3[3], ROUND_OUT_s2[3], ROUND_OUT_s1[3], ROUND_OUT_s0[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U29 ( .a ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, new_AGEMA_signal_2648, SHIFTROWS[35]}), .b ({new_AGEMA_signal_3022, new_AGEMA_signal_3021, new_AGEMA_signal_3020, SHIFTROWS[67]}), .c ({ROUND_OUT_s3[35], ROUND_OUT_s2[35], ROUND_OUT_s1[35], ROUND_OUT_s0[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U25 ( .a ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, new_AGEMA_signal_2654, SHIFTROWS[39]}), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, new_AGEMA_signal_3017, SHIFTROWS[71]}), .c ({ROUND_OUT_s3[39], ROUND_OUT_s2[39], ROUND_OUT_s1[39], ROUND_OUT_s0[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U21 ( .a ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, new_AGEMA_signal_2657, SHIFTROWS[43]}), .b ({new_AGEMA_signal_3016, new_AGEMA_signal_3015, new_AGEMA_signal_3014, SHIFTROWS[75]}), .c ({ROUND_OUT_s3[43], ROUND_OUT_s2[43], ROUND_OUT_s1[43], ROUND_OUT_s0[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U17 ( .a ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, new_AGEMA_signal_2663, SHIFTROWS[47]}), .b ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, new_AGEMA_signal_3011, SHIFTROWS[79]}), .c ({ROUND_OUT_s3[47], ROUND_OUT_s2[47], ROUND_OUT_s1[47], ROUND_OUT_s0[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U13 ( .a ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, new_AGEMA_signal_2630, SHIFTROWS[51]}), .b ({new_AGEMA_signal_3010, new_AGEMA_signal_3009, new_AGEMA_signal_3008, SHIFTROWS[83]}), .c ({ROUND_OUT_s3[51], ROUND_OUT_s2[51], ROUND_OUT_s1[51], ROUND_OUT_s0[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U9 ( .a ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, new_AGEMA_signal_2636, SHIFTROWS[55]}), .b ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, new_AGEMA_signal_3005, SHIFTROWS[87]}), .c ({ROUND_OUT_s3[55], ROUND_OUT_s2[55], ROUND_OUT_s1[55], ROUND_OUT_s0[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U5 ( .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, SHIFTROWS[59]}), .b ({new_AGEMA_signal_3028, new_AGEMA_signal_3027, new_AGEMA_signal_3026, SHIFTROWS[91]}), .c ({ROUND_OUT_s3[59], ROUND_OUT_s2[59], ROUND_OUT_s1[59], ROUND_OUT_s0[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U1 ( .a ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, new_AGEMA_signal_2645, SHIFTROWS[63]}), .b ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, new_AGEMA_signal_3023, SHIFTROWS[95]}), .c ({ROUND_OUT_s3[63], ROUND_OUT_s2[63], ROUND_OUT_s1[63], ROUND_OUT_s0[63]}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    not_masked #(.security_order(3), .pipeline(0)) U399 ( .a ({new_AGEMA_signal_3094, new_AGEMA_signal_3093, new_AGEMA_signal_3092, SUBSTITUTION_57}), .b ({new_AGEMA_signal_3184, new_AGEMA_signal_3183, new_AGEMA_signal_3182, SHIFTROWS[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U407 ( .a ({ROUND_KEY_s3[353], ROUND_KEY_s2[353], ROUND_KEY_s1[353], ROUND_KEY_s0[353]}), .b ({new_AGEMA_signal_3124, new_AGEMA_signal_3123, new_AGEMA_signal_3122, CONST_ADDITION[97]}), .c ({new_AGEMA_signal_3190, new_AGEMA_signal_3189, new_AGEMA_signal_3188, n409}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U408 ( .a ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, n410}), .b ({new_AGEMA_signal_3190, new_AGEMA_signal_3189, new_AGEMA_signal_3188, n409}), .c ({ROUND_OUT_s3[65], ROUND_OUT_s2[65], ROUND_OUT_s1[65], ROUND_OUT_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U422 ( .a ({ROUND_KEY_s3[348], ROUND_KEY_s2[348], ROUND_KEY_s1[348], ROUND_KEY_s0[348]}), .b ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, new_AGEMA_signal_3119, CONST_ADDITION[92]}), .c ({new_AGEMA_signal_3196, new_AGEMA_signal_3195, new_AGEMA_signal_3194, n419}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U423 ( .a ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, n420}), .b ({new_AGEMA_signal_3196, new_AGEMA_signal_3195, new_AGEMA_signal_3194, n419}), .c ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, new_AGEMA_signal_3383, SHIFTROWS[84]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U431 ( .a ({new_AGEMA_signal_3118, new_AGEMA_signal_3117, new_AGEMA_signal_3116, SUBSTITUTION_89}), .b ({ROUND_KEY_s3[345], ROUND_KEY_s2[345], ROUND_KEY_s1[345], ROUND_KEY_s0[345]}), .c ({new_AGEMA_signal_3202, new_AGEMA_signal_3201, new_AGEMA_signal_3200, n425}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U432 ( .a ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, n426}), .b ({new_AGEMA_signal_3202, new_AGEMA_signal_3201, new_AGEMA_signal_3200, n425}), .c ({new_AGEMA_signal_3388, new_AGEMA_signal_3387, new_AGEMA_signal_3386, n427}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U433 ( .a ({1'b0, 1'b0, 1'b0, CONST_IN[5]}), .b ({new_AGEMA_signal_3388, new_AGEMA_signal_3387, new_AGEMA_signal_3386, n427}), .c ({new_AGEMA_signal_3508, new_AGEMA_signal_3507, new_AGEMA_signal_3506, SHIFTROWS[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U448 ( .a ({ROUND_KEY_s3[340], ROUND_KEY_s2[340], ROUND_KEY_s1[340], ROUND_KEY_s0[340]}), .b ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, new_AGEMA_signal_3113, CONST_ADDITION[84]}), .c ({new_AGEMA_signal_3208, new_AGEMA_signal_3207, new_AGEMA_signal_3206, n437}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U449 ( .a ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, n438}), .b ({new_AGEMA_signal_3208, new_AGEMA_signal_3207, new_AGEMA_signal_3206, n437}), .c ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, new_AGEMA_signal_3389, SHIFTROWS[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U457 ( .a ({ROUND_KEY_s3[337], ROUND_KEY_s2[337], ROUND_KEY_s1[337], ROUND_KEY_s0[337]}), .b ({new_AGEMA_signal_3112, new_AGEMA_signal_3111, new_AGEMA_signal_3110, CONST_ADDITION[81]}), .c ({new_AGEMA_signal_3214, new_AGEMA_signal_3213, new_AGEMA_signal_3212, n443}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U458 ( .a ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, new_AGEMA_signal_1250, n444}), .b ({new_AGEMA_signal_3214, new_AGEMA_signal_3213, new_AGEMA_signal_3212, n443}), .c ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, new_AGEMA_signal_3392, SHIFTROWS[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U472 ( .a ({ROUND_KEY_s3[332], ROUND_KEY_s2[332], ROUND_KEY_s1[332], ROUND_KEY_s0[332]}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3107, CONST_ADDITION[76]}), .c ({new_AGEMA_signal_3220, new_AGEMA_signal_3219, new_AGEMA_signal_3218, n453}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U473 ( .a ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, new_AGEMA_signal_1295, n454}), .b ({new_AGEMA_signal_3220, new_AGEMA_signal_3219, new_AGEMA_signal_3218, n453}), .c ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, new_AGEMA_signal_3395, SHIFTROWS[68]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U481 ( .a ({ROUND_KEY_s3[329], ROUND_KEY_s2[329], ROUND_KEY_s1[329], ROUND_KEY_s0[329]}), .b ({new_AGEMA_signal_3106, new_AGEMA_signal_3105, new_AGEMA_signal_3104, CONST_ADDITION[73]}), .c ({new_AGEMA_signal_3226, new_AGEMA_signal_3225, new_AGEMA_signal_3224, n459}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U482 ( .a ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, n460}), .b ({new_AGEMA_signal_3226, new_AGEMA_signal_3225, new_AGEMA_signal_3224, n459}), .c ({new_AGEMA_signal_3400, new_AGEMA_signal_3399, new_AGEMA_signal_3398, SHIFTROWS[65]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U496 ( .a ({ROUND_KEY_s3[324], ROUND_KEY_s2[324], ROUND_KEY_s1[324], ROUND_KEY_s0[324]}), .b ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, new_AGEMA_signal_3101, CONST_ADDITION[68]}), .c ({new_AGEMA_signal_3232, new_AGEMA_signal_3231, new_AGEMA_signal_3230, n469}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U497 ( .a ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, n470}), .b ({new_AGEMA_signal_3232, new_AGEMA_signal_3231, new_AGEMA_signal_3230, n469}), .c ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, new_AGEMA_signal_3401, SHIFTROWS[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U505 ( .a ({ROUND_KEY_s3[321], ROUND_KEY_s2[321], ROUND_KEY_s1[321], ROUND_KEY_s0[321]}), .b ({new_AGEMA_signal_3100, new_AGEMA_signal_3099, new_AGEMA_signal_3098, CONST_ADDITION[65]}), .c ({new_AGEMA_signal_3238, new_AGEMA_signal_3237, new_AGEMA_signal_3236, n475}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U506 ( .a ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, n476}), .b ({new_AGEMA_signal_3238, new_AGEMA_signal_3237, new_AGEMA_signal_3236, n475}), .c ({new_AGEMA_signal_3406, new_AGEMA_signal_3405, new_AGEMA_signal_3404, SHIFTROWS[89]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U520 ( .a ({ROUND_KEY_s3[380], ROUND_KEY_s2[380], ROUND_KEY_s1[380], ROUND_KEY_s0[380]}), .b ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, new_AGEMA_signal_3143, CONST_ADDITION[124]}), .c ({new_AGEMA_signal_3244, new_AGEMA_signal_3243, new_AGEMA_signal_3242, n485}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U521 ( .a ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, n486}), .b ({new_AGEMA_signal_3244, new_AGEMA_signal_3243, new_AGEMA_signal_3242, n485}), .c ({ROUND_OUT_s3[92], ROUND_OUT_s2[92], ROUND_OUT_s1[92], ROUND_OUT_s0[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U531 ( .a ({new_AGEMA_signal_3142, new_AGEMA_signal_3141, new_AGEMA_signal_3140, SUBSTITUTION[121]}), .b ({ROUND_KEY_s3[377], ROUND_KEY_s2[377], ROUND_KEY_s1[377], ROUND_KEY_s0[377]}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, new_AGEMA_signal_3251, n493}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U532 ( .a ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, new_AGEMA_signal_1466, n494}), .b ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, new_AGEMA_signal_3251, n493}), .c ({new_AGEMA_signal_3412, new_AGEMA_signal_3411, new_AGEMA_signal_3410, n495}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U533 ( .a ({1'b0, 1'b0, 1'b0, CONST_IN[1]}), .b ({new_AGEMA_signal_3412, new_AGEMA_signal_3411, new_AGEMA_signal_3410, n495}), .c ({ROUND_OUT_s3[89], ROUND_OUT_s2[89], ROUND_OUT_s1[89], ROUND_OUT_s0[89]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U548 ( .a ({ROUND_KEY_s3[372], ROUND_KEY_s2[372], ROUND_KEY_s1[372], ROUND_KEY_s0[372]}), .b ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, new_AGEMA_signal_3137, CONST_ADDITION[116]}), .c ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, new_AGEMA_signal_3257, n505}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U549 ( .a ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, new_AGEMA_signal_1511, n506}), .b ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, new_AGEMA_signal_3257, n505}), .c ({ROUND_OUT_s3[84], ROUND_OUT_s2[84], ROUND_OUT_s1[84], ROUND_OUT_s0[84]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U557 ( .a ({ROUND_KEY_s3[369], ROUND_KEY_s2[369], ROUND_KEY_s1[369], ROUND_KEY_s0[369]}), .b ({new_AGEMA_signal_3136, new_AGEMA_signal_3135, new_AGEMA_signal_3134, CONST_ADDITION[113]}), .c ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, new_AGEMA_signal_3263, n511}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U558 ( .a ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, new_AGEMA_signal_1538, n512}), .b ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, new_AGEMA_signal_3263, n511}), .c ({ROUND_OUT_s3[81], ROUND_OUT_s2[81], ROUND_OUT_s1[81], ROUND_OUT_s0[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U572 ( .a ({ROUND_KEY_s3[364], ROUND_KEY_s2[364], ROUND_KEY_s1[364], ROUND_KEY_s0[364]}), .b ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, new_AGEMA_signal_3131, CONST_ADDITION[108]}), .c ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, new_AGEMA_signal_3269, n521}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U573 ( .a ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, new_AGEMA_signal_1583, n522}), .b ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, new_AGEMA_signal_3269, n521}), .c ({ROUND_OUT_s3[76], ROUND_OUT_s2[76], ROUND_OUT_s1[76], ROUND_OUT_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U581 ( .a ({ROUND_KEY_s3[361], ROUND_KEY_s2[361], ROUND_KEY_s1[361], ROUND_KEY_s0[361]}), .b ({new_AGEMA_signal_3130, new_AGEMA_signal_3129, new_AGEMA_signal_3128, CONST_ADDITION[105]}), .c ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, new_AGEMA_signal_3275, n527}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U582 ( .a ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1610, n528}), .b ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, new_AGEMA_signal_3275, n527}), .c ({ROUND_OUT_s3[73], ROUND_OUT_s2[73], ROUND_OUT_s1[73], ROUND_OUT_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U596 ( .a ({ROUND_KEY_s3[356], ROUND_KEY_s2[356], ROUND_KEY_s1[356], ROUND_KEY_s0[356]}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, new_AGEMA_signal_3125, CONST_ADDITION[100]}), .c ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, new_AGEMA_signal_3281, n537}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U597 ( .a ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, new_AGEMA_signal_1655, n538}), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, new_AGEMA_signal_3281, n537}), .c ({ROUND_OUT_s3[68], ROUND_OUT_s2[68], ROUND_OUT_s1[68], ROUND_OUT_s0[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_0_U7 ( .a ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, new_AGEMA_signal_2837, S_0_R2[2]}), .b ({ROUND_IN_s3[7], ROUND_IN_s2[7], ROUND_IN_s1[7], ROUND_IN_s0[7]}), .c ({new_AGEMA_signal_3052, new_AGEMA_signal_3051, new_AGEMA_signal_3050, SHIFTROWS[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_0_U4 ( .a ({new_AGEMA_signal_2842, new_AGEMA_signal_2841, new_AGEMA_signal_2840, S_0_R1[3]}), .b ({ROUND_IN_s3[3], ROUND_IN_s2[3], ROUND_IN_s1[3], ROUND_IN_s0[3]}), .c ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, new_AGEMA_signal_3053, SHIFTROWS[12]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_0_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, new_AGEMA_signal_2600, SHIFTROWS[15]}), .b ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, SHIFTROWS[10]}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, new_AGEMA_signal_2837, S_0_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_0_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, SHIFTROWS[14]}), .b ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, new_AGEMA_signal_2600, SHIFTROWS[15]}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_2842, new_AGEMA_signal_2841, new_AGEMA_signal_2840, S_0_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_1_U7 ( .a ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, new_AGEMA_signal_2843, S_1_R2[2]}), .b ({ROUND_IN_s3[15], ROUND_IN_s2[15], ROUND_IN_s1[15], ROUND_IN_s0[15]}), .c ({new_AGEMA_signal_3058, new_AGEMA_signal_3057, new_AGEMA_signal_3056, SHIFTROWS[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_1_U4 ( .a ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, S_1_R1[3]}), .b ({ROUND_IN_s3[11], ROUND_IN_s2[11], ROUND_IN_s1[11], ROUND_IN_s0[11]}), .c ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, new_AGEMA_signal_3059, SHIFTROWS[20]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_1_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, new_AGEMA_signal_2609, SHIFTROWS[23]}), .b ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, new_AGEMA_signal_2057, SHIFTROWS[18]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, new_AGEMA_signal_2843, S_1_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_1_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, SHIFTROWS[22]}), .b ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, new_AGEMA_signal_2609, SHIFTROWS[23]}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, S_1_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_2_U7 ( .a ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, new_AGEMA_signal_2849, S_2_R2[2]}), .b ({ROUND_IN_s3[23], ROUND_IN_s2[23], ROUND_IN_s1[23], ROUND_IN_s0[23]}), .c ({new_AGEMA_signal_3064, new_AGEMA_signal_3063, new_AGEMA_signal_3062, SHIFTROWS[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_2_U4 ( .a ({new_AGEMA_signal_2854, new_AGEMA_signal_2853, new_AGEMA_signal_2852, S_2_R1[3]}), .b ({ROUND_IN_s3[19], ROUND_IN_s2[19], ROUND_IN_s1[19], ROUND_IN_s0[19]}), .c ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, new_AGEMA_signal_3065, SHIFTROWS[28]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_2_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, new_AGEMA_signal_2618, SHIFTROWS[31]}), .b ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, SHIFTROWS[26]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, new_AGEMA_signal_2849, S_2_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_2_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, SHIFTROWS[30]}), .b ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, new_AGEMA_signal_2618, SHIFTROWS[31]}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_2854, new_AGEMA_signal_2853, new_AGEMA_signal_2852, S_2_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_3_U7 ( .a ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, new_AGEMA_signal_2855, S_3_R2[2]}), .b ({ROUND_IN_s3[31], ROUND_IN_s2[31], ROUND_IN_s1[31], ROUND_IN_s0[31]}), .c ({new_AGEMA_signal_3070, new_AGEMA_signal_3069, new_AGEMA_signal_3068, SHIFTROWS[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_3_U4 ( .a ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, new_AGEMA_signal_2858, S_3_R1[3]}), .b ({ROUND_IN_s3[27], ROUND_IN_s2[27], ROUND_IN_s1[27], ROUND_IN_s0[27]}), .c ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, new_AGEMA_signal_3071, SHIFTROWS[4]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_3_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, new_AGEMA_signal_2627, SHIFTROWS[7]}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, SHIFTROWS[2]}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, new_AGEMA_signal_2855, S_3_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_3_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, SHIFTROWS[6]}), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, new_AGEMA_signal_2627, SHIFTROWS[7]}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, new_AGEMA_signal_2858, S_3_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_4_U7 ( .a ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, new_AGEMA_signal_2861, S_4_R2[2]}), .b ({ROUND_IN_s3[39], ROUND_IN_s2[39], ROUND_IN_s1[39], ROUND_IN_s0[39]}), .c ({new_AGEMA_signal_3076, new_AGEMA_signal_3075, new_AGEMA_signal_3074, SHIFTROWS[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_4_U4 ( .a ({new_AGEMA_signal_2866, new_AGEMA_signal_2865, new_AGEMA_signal_2864, S_4_R1[3]}), .b ({ROUND_IN_s3[35], ROUND_IN_s2[35], ROUND_IN_s1[35], ROUND_IN_s0[35]}), .c ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, new_AGEMA_signal_3077, SHIFTROWS[52]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_4_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, new_AGEMA_signal_2636, SHIFTROWS[55]}), .b ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, SHIFTROWS[50]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, new_AGEMA_signal_2861, S_4_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_4_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, new_AGEMA_signal_2114, SHIFTROWS[54]}), .b ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, new_AGEMA_signal_2636, SHIFTROWS[55]}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_2866, new_AGEMA_signal_2865, new_AGEMA_signal_2864, S_4_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_5_U7 ( .a ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, new_AGEMA_signal_2867, S_5_R2[2]}), .b ({ROUND_IN_s3[47], ROUND_IN_s2[47], ROUND_IN_s1[47], ROUND_IN_s0[47]}), .c ({new_AGEMA_signal_3082, new_AGEMA_signal_3081, new_AGEMA_signal_3080, SHIFTROWS[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_5_U4 ( .a ({new_AGEMA_signal_2872, new_AGEMA_signal_2871, new_AGEMA_signal_2870, S_5_R1[3]}), .b ({ROUND_IN_s3[43], ROUND_IN_s2[43], ROUND_IN_s1[43], ROUND_IN_s0[43]}), .c ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, new_AGEMA_signal_3083, SHIFTROWS[60]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_5_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, new_AGEMA_signal_2645, SHIFTROWS[63]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, new_AGEMA_signal_2117, SHIFTROWS[58]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, new_AGEMA_signal_2867, S_5_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_5_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, new_AGEMA_signal_2129, SHIFTROWS[62]}), .b ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, new_AGEMA_signal_2645, SHIFTROWS[63]}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_2872, new_AGEMA_signal_2871, new_AGEMA_signal_2870, S_5_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_6_U7 ( .a ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, new_AGEMA_signal_2873, S_6_R2[2]}), .b ({ROUND_IN_s3[55], ROUND_IN_s2[55], ROUND_IN_s1[55], ROUND_IN_s0[55]}), .c ({new_AGEMA_signal_3088, new_AGEMA_signal_3087, new_AGEMA_signal_3086, SHIFTROWS[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_6_U4 ( .a ({new_AGEMA_signal_2878, new_AGEMA_signal_2877, new_AGEMA_signal_2876, S_6_R1[3]}), .b ({ROUND_IN_s3[51], ROUND_IN_s2[51], ROUND_IN_s1[51], ROUND_IN_s0[51]}), .c ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, new_AGEMA_signal_3089, SHIFTROWS[36]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_6_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, new_AGEMA_signal_2654, SHIFTROWS[39]}), .b ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, new_AGEMA_signal_2132, SHIFTROWS[34]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, new_AGEMA_signal_2873, S_6_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_6_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, SHIFTROWS[38]}), .b ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, new_AGEMA_signal_2654, SHIFTROWS[39]}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_2878, new_AGEMA_signal_2877, new_AGEMA_signal_2876, S_6_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_7_U7 ( .a ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, new_AGEMA_signal_2879, S_7_R2[2]}), .b ({ROUND_IN_s3[63], ROUND_IN_s2[63], ROUND_IN_s1[63], ROUND_IN_s0[63]}), .c ({new_AGEMA_signal_3094, new_AGEMA_signal_3093, new_AGEMA_signal_3092, SUBSTITUTION_57}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_7_U4 ( .a ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, new_AGEMA_signal_2882, S_7_R1[3]}), .b ({ROUND_IN_s3[59], ROUND_IN_s2[59], ROUND_IN_s1[59], ROUND_IN_s0[59]}), .c ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, new_AGEMA_signal_3095, SHIFTROWS[44]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_7_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, new_AGEMA_signal_2663, SHIFTROWS[47]}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, new_AGEMA_signal_2147, SHIFTROWS[42]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, new_AGEMA_signal_2879, S_7_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_7_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, new_AGEMA_signal_2159, SHIFTROWS[46]}), .b ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, new_AGEMA_signal_2663, SHIFTROWS[47]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, new_AGEMA_signal_2882, S_7_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_8_U7 ( .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, new_AGEMA_signal_2885, S_8_R2[2]}), .b ({ROUND_IN_s3[71], ROUND_IN_s2[71], ROUND_IN_s1[71], ROUND_IN_s0[71]}), .c ({new_AGEMA_signal_3100, new_AGEMA_signal_3099, new_AGEMA_signal_3098, CONST_ADDITION[65]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_8_U4 ( .a ({new_AGEMA_signal_2890, new_AGEMA_signal_2889, new_AGEMA_signal_2888, S_8_R1[3]}), .b ({ROUND_IN_s3[67], ROUND_IN_s2[67], ROUND_IN_s1[67], ROUND_IN_s0[67]}), .c ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, new_AGEMA_signal_3101, CONST_ADDITION[68]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_8_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, new_AGEMA_signal_2672, CONST_ADDITION[71]}), .b ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, CONST_ADDITION[66]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, new_AGEMA_signal_2885, S_8_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_8_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, CONST_ADDITION[70]}), .b ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, new_AGEMA_signal_2672, CONST_ADDITION[71]}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_2890, new_AGEMA_signal_2889, new_AGEMA_signal_2888, S_8_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_9_U7 ( .a ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, new_AGEMA_signal_2891, S_9_R2[2]}), .b ({ROUND_IN_s3[79], ROUND_IN_s2[79], ROUND_IN_s1[79], ROUND_IN_s0[79]}), .c ({new_AGEMA_signal_3106, new_AGEMA_signal_3105, new_AGEMA_signal_3104, CONST_ADDITION[73]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_9_U4 ( .a ({new_AGEMA_signal_2896, new_AGEMA_signal_2895, new_AGEMA_signal_2894, S_9_R1[3]}), .b ({ROUND_IN_s3[75], ROUND_IN_s2[75], ROUND_IN_s1[75], ROUND_IN_s0[75]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3107, CONST_ADDITION[76]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_9_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, new_AGEMA_signal_2681, CONST_ADDITION[79]}), .b ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, CONST_ADDITION[74]}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, new_AGEMA_signal_2891, S_9_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_9_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, CONST_ADDITION[78]}), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, new_AGEMA_signal_2681, CONST_ADDITION[79]}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_2896, new_AGEMA_signal_2895, new_AGEMA_signal_2894, S_9_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_10_U7 ( .a ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, new_AGEMA_signal_2897, S_10_R2[2]}), .b ({ROUND_IN_s3[87], ROUND_IN_s2[87], ROUND_IN_s1[87], ROUND_IN_s0[87]}), .c ({new_AGEMA_signal_3112, new_AGEMA_signal_3111, new_AGEMA_signal_3110, CONST_ADDITION[81]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_10_U4 ( .a ({new_AGEMA_signal_2902, new_AGEMA_signal_2901, new_AGEMA_signal_2900, S_10_R1[3]}), .b ({ROUND_IN_s3[83], ROUND_IN_s2[83], ROUND_IN_s1[83], ROUND_IN_s0[83]}), .c ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, new_AGEMA_signal_3113, CONST_ADDITION[84]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_10_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, CONST_ADDITION[87]}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, new_AGEMA_signal_2192, CONST_ADDITION[82]}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, new_AGEMA_signal_2897, S_10_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_10_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, new_AGEMA_signal_2204, CONST_ADDITION[86]}), .b ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, new_AGEMA_signal_2690, CONST_ADDITION[87]}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_2902, new_AGEMA_signal_2901, new_AGEMA_signal_2900, S_10_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_11_U7 ( .a ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, new_AGEMA_signal_2903, S_11_R2[2]}), .b ({ROUND_IN_s3[95], ROUND_IN_s2[95], ROUND_IN_s1[95], ROUND_IN_s0[95]}), .c ({new_AGEMA_signal_3118, new_AGEMA_signal_3117, new_AGEMA_signal_3116, SUBSTITUTION_89}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_11_U4 ( .a ({new_AGEMA_signal_2908, new_AGEMA_signal_2907, new_AGEMA_signal_2906, S_11_R1[3]}), .b ({ROUND_IN_s3[91], ROUND_IN_s2[91], ROUND_IN_s1[91], ROUND_IN_s0[91]}), .c ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, new_AGEMA_signal_3119, CONST_ADDITION[92]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_11_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, CONST_ADDITION[95]}), .b ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, new_AGEMA_signal_2207, CONST_ADDITION[90]}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, new_AGEMA_signal_2903, S_11_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_11_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, new_AGEMA_signal_2219, CONST_ADDITION[94]}), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_2699, CONST_ADDITION[95]}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_2908, new_AGEMA_signal_2907, new_AGEMA_signal_2906, S_11_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_12_U7 ( .a ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, new_AGEMA_signal_2909, S_12_R2[2]}), .b ({ROUND_IN_s3[103], ROUND_IN_s2[103], ROUND_IN_s1[103], ROUND_IN_s0[103]}), .c ({new_AGEMA_signal_3124, new_AGEMA_signal_3123, new_AGEMA_signal_3122, CONST_ADDITION[97]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_12_U4 ( .a ({new_AGEMA_signal_2914, new_AGEMA_signal_2913, new_AGEMA_signal_2912, S_12_R1[3]}), .b ({ROUND_IN_s3[99], ROUND_IN_s2[99], ROUND_IN_s1[99], ROUND_IN_s0[99]}), .c ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, new_AGEMA_signal_3125, CONST_ADDITION[100]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_12_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, CONST_ADDITION[103]}), .b ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, CONST_ADDITION[98]}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, new_AGEMA_signal_2909, S_12_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_12_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, CONST_ADDITION[102]}), .b ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, CONST_ADDITION[103]}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_2914, new_AGEMA_signal_2913, new_AGEMA_signal_2912, S_12_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_13_U7 ( .a ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, new_AGEMA_signal_2915, S_13_R2[2]}), .b ({ROUND_IN_s3[111], ROUND_IN_s2[111], ROUND_IN_s1[111], ROUND_IN_s0[111]}), .c ({new_AGEMA_signal_3130, new_AGEMA_signal_3129, new_AGEMA_signal_3128, CONST_ADDITION[105]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_13_U4 ( .a ({new_AGEMA_signal_2920, new_AGEMA_signal_2919, new_AGEMA_signal_2918, S_13_R1[3]}), .b ({ROUND_IN_s3[107], ROUND_IN_s2[107], ROUND_IN_s1[107], ROUND_IN_s0[107]}), .c ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, new_AGEMA_signal_3131, CONST_ADDITION[108]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_13_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, new_AGEMA_signal_2717, CONST_ADDITION[111]}), .b ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, new_AGEMA_signal_2237, CONST_ADDITION[106]}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, new_AGEMA_signal_2915, S_13_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_13_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, new_AGEMA_signal_2249, CONST_ADDITION[110]}), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, new_AGEMA_signal_2717, CONST_ADDITION[111]}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_2920, new_AGEMA_signal_2919, new_AGEMA_signal_2918, S_13_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_14_U7 ( .a ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, new_AGEMA_signal_2921, S_14_R2[2]}), .b ({ROUND_IN_s3[119], ROUND_IN_s2[119], ROUND_IN_s1[119], ROUND_IN_s0[119]}), .c ({new_AGEMA_signal_3136, new_AGEMA_signal_3135, new_AGEMA_signal_3134, CONST_ADDITION[113]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_14_U4 ( .a ({new_AGEMA_signal_2926, new_AGEMA_signal_2925, new_AGEMA_signal_2924, S_14_R1[3]}), .b ({ROUND_IN_s3[115], ROUND_IN_s2[115], ROUND_IN_s1[115], ROUND_IN_s0[115]}), .c ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, new_AGEMA_signal_3137, CONST_ADDITION[116]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_14_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, CONST_ADDITION[119]}), .b ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, new_AGEMA_signal_2252, CONST_ADDITION[114]}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, new_AGEMA_signal_2921, S_14_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_14_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, new_AGEMA_signal_2264, CONST_ADDITION[118]}), .b ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, CONST_ADDITION[119]}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_2926, new_AGEMA_signal_2925, new_AGEMA_signal_2924, S_14_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_15_U7 ( .a ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, new_AGEMA_signal_2927, S_15_R2[2]}), .b ({ROUND_IN_s3[127], ROUND_IN_s2[127], ROUND_IN_s1[127], ROUND_IN_s0[127]}), .c ({new_AGEMA_signal_3142, new_AGEMA_signal_3141, new_AGEMA_signal_3140, SUBSTITUTION[121]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_15_U4 ( .a ({new_AGEMA_signal_2932, new_AGEMA_signal_2931, new_AGEMA_signal_2930, S_15_R1[3]}), .b ({ROUND_IN_s3[123], ROUND_IN_s2[123], ROUND_IN_s1[123], ROUND_IN_s0[123]}), .c ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, new_AGEMA_signal_3143, CONST_ADDITION[124]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_15_NOR2Inst_2_U1 ( .a ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, new_AGEMA_signal_2735, CONST_ADDITION[127]}), .b ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, new_AGEMA_signal_2267, SUBSTITUTION[122]}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, new_AGEMA_signal_2927, S_15_R2[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_15_NOR1Inst_3_U1 ( .a ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, new_AGEMA_signal_2279, CONST_ADDITION[126]}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, new_AGEMA_signal_2735, CONST_ADDITION[127]}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_2932, new_AGEMA_signal_2931, new_AGEMA_signal_2930, S_15_R1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U90 ( .a ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, new_AGEMA_signal_3065, SHIFTROWS[28]}), .b ({ROUND_OUT_s3[28], ROUND_OUT_s2[28], ROUND_OUT_s1[28], ROUND_OUT_s0[28]}), .c ({ROUND_OUT_s3[124], ROUND_OUT_s2[124], ROUND_OUT_s1[124], ROUND_OUT_s0[124]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U89 ( .a ({ROUND_OUT_s3[92], ROUND_OUT_s2[92], ROUND_OUT_s1[92], ROUND_OUT_s0[92]}), .b ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, new_AGEMA_signal_3083, SHIFTROWS[60]}), .c ({ROUND_OUT_s3[28], ROUND_OUT_s2[28], ROUND_OUT_s1[28], ROUND_OUT_s0[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U72 ( .a ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, new_AGEMA_signal_3053, SHIFTROWS[12]}), .b ({ROUND_OUT_s3[12], ROUND_OUT_s2[12], ROUND_OUT_s1[12], ROUND_OUT_s0[12]}), .c ({ROUND_OUT_s3[108], ROUND_OUT_s2[108], ROUND_OUT_s1[108], ROUND_OUT_s0[108]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U71 ( .a ({ROUND_OUT_s3[76], ROUND_OUT_s2[76], ROUND_OUT_s1[76], ROUND_OUT_s0[76]}), .b ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, new_AGEMA_signal_3095, SHIFTROWS[44]}), .c ({ROUND_OUT_s3[12], ROUND_OUT_s2[12], ROUND_OUT_s1[12], ROUND_OUT_s0[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U64 ( .a ({new_AGEMA_signal_3052, new_AGEMA_signal_3051, new_AGEMA_signal_3050, SHIFTROWS[9]}), .b ({ROUND_OUT_s3[9], ROUND_OUT_s2[9], ROUND_OUT_s1[9], ROUND_OUT_s0[9]}), .c ({ROUND_OUT_s3[105], ROUND_OUT_s2[105], ROUND_OUT_s1[105], ROUND_OUT_s0[105]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U63 ( .a ({ROUND_OUT_s3[73], ROUND_OUT_s2[73], ROUND_OUT_s1[73], ROUND_OUT_s0[73]}), .b ({new_AGEMA_signal_3184, new_AGEMA_signal_3183, new_AGEMA_signal_3182, SHIFTROWS[41]}), .c ({ROUND_OUT_s3[9], ROUND_OUT_s2[9], ROUND_OUT_s1[9], ROUND_OUT_s0[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U58 ( .a ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, new_AGEMA_signal_3059, SHIFTROWS[20]}), .b ({ROUND_OUT_s3[20], ROUND_OUT_s2[20], ROUND_OUT_s1[20], ROUND_OUT_s0[20]}), .c ({ROUND_OUT_s3[116], ROUND_OUT_s2[116], ROUND_OUT_s1[116], ROUND_OUT_s0[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U57 ( .a ({ROUND_OUT_s3[84], ROUND_OUT_s2[84], ROUND_OUT_s1[84], ROUND_OUT_s0[84]}), .b ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, new_AGEMA_signal_3077, SHIFTROWS[52]}), .c ({ROUND_OUT_s3[20], ROUND_OUT_s2[20], ROUND_OUT_s1[20], ROUND_OUT_s0[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U46 ( .a ({new_AGEMA_signal_3064, new_AGEMA_signal_3063, new_AGEMA_signal_3062, SHIFTROWS[25]}), .b ({ROUND_OUT_s3[25], ROUND_OUT_s2[25], ROUND_OUT_s1[25], ROUND_OUT_s0[25]}), .c ({ROUND_OUT_s3[121], ROUND_OUT_s2[121], ROUND_OUT_s1[121], ROUND_OUT_s0[121]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U45 ( .a ({ROUND_OUT_s3[89], ROUND_OUT_s2[89], ROUND_OUT_s1[89], ROUND_OUT_s0[89]}), .b ({new_AGEMA_signal_3082, new_AGEMA_signal_3081, new_AGEMA_signal_3080, SHIFTROWS[57]}), .c ({ROUND_OUT_s3[25], ROUND_OUT_s2[25], ROUND_OUT_s1[25], ROUND_OUT_s0[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U42 ( .a ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, new_AGEMA_signal_3071, SHIFTROWS[4]}), .b ({ROUND_OUT_s3[4], ROUND_OUT_s2[4], ROUND_OUT_s1[4], ROUND_OUT_s0[4]}), .c ({ROUND_OUT_s3[100], ROUND_OUT_s2[100], ROUND_OUT_s1[100], ROUND_OUT_s0[100]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U41 ( .a ({ROUND_OUT_s3[68], ROUND_OUT_s2[68], ROUND_OUT_s1[68], ROUND_OUT_s0[68]}), .b ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, new_AGEMA_signal_3089, SHIFTROWS[36]}), .c ({ROUND_OUT_s3[4], ROUND_OUT_s2[4], ROUND_OUT_s1[4], ROUND_OUT_s0[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U38 ( .a ({new_AGEMA_signal_3058, new_AGEMA_signal_3057, new_AGEMA_signal_3056, SHIFTROWS[17]}), .b ({ROUND_OUT_s3[17], ROUND_OUT_s2[17], ROUND_OUT_s1[17], ROUND_OUT_s0[17]}), .c ({ROUND_OUT_s3[113], ROUND_OUT_s2[113], ROUND_OUT_s1[113], ROUND_OUT_s0[113]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U37 ( .a ({ROUND_OUT_s3[81], ROUND_OUT_s2[81], ROUND_OUT_s1[81], ROUND_OUT_s0[81]}), .b ({new_AGEMA_signal_3076, new_AGEMA_signal_3075, new_AGEMA_signal_3074, SHIFTROWS[49]}), .c ({ROUND_OUT_s3[17], ROUND_OUT_s2[17], ROUND_OUT_s1[17], ROUND_OUT_s0[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U34 ( .a ({new_AGEMA_signal_3070, new_AGEMA_signal_3069, new_AGEMA_signal_3068, SHIFTROWS[1]}), .b ({ROUND_OUT_s3[1], ROUND_OUT_s2[1], ROUND_OUT_s1[1], ROUND_OUT_s0[1]}), .c ({ROUND_OUT_s3[97], ROUND_OUT_s2[97], ROUND_OUT_s1[97], ROUND_OUT_s0[97]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U33 ( .a ({ROUND_OUT_s3[65], ROUND_OUT_s2[65], ROUND_OUT_s1[65], ROUND_OUT_s0[65]}), .b ({new_AGEMA_signal_3088, new_AGEMA_signal_3087, new_AGEMA_signal_3086, SHIFTROWS[33]}), .c ({ROUND_OUT_s3[1], ROUND_OUT_s2[1], ROUND_OUT_s1[1], ROUND_OUT_s0[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U31 ( .a ({new_AGEMA_signal_3088, new_AGEMA_signal_3087, new_AGEMA_signal_3086, SHIFTROWS[33]}), .b ({new_AGEMA_signal_3400, new_AGEMA_signal_3399, new_AGEMA_signal_3398, SHIFTROWS[65]}), .c ({ROUND_OUT_s3[33], ROUND_OUT_s2[33], ROUND_OUT_s1[33], ROUND_OUT_s0[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U28 ( .a ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, new_AGEMA_signal_3089, SHIFTROWS[36]}), .b ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, new_AGEMA_signal_3395, SHIFTROWS[68]}), .c ({ROUND_OUT_s3[36], ROUND_OUT_s2[36], ROUND_OUT_s1[36], ROUND_OUT_s0[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U23 ( .a ({new_AGEMA_signal_3184, new_AGEMA_signal_3183, new_AGEMA_signal_3182, SHIFTROWS[41]}), .b ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, new_AGEMA_signal_3392, SHIFTROWS[73]}), .c ({ROUND_OUT_s3[41], ROUND_OUT_s2[41], ROUND_OUT_s1[41], ROUND_OUT_s0[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U20 ( .a ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, new_AGEMA_signal_3095, SHIFTROWS[44]}), .b ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, new_AGEMA_signal_3389, SHIFTROWS[76]}), .c ({ROUND_OUT_s3[44], ROUND_OUT_s2[44], ROUND_OUT_s1[44], ROUND_OUT_s0[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U15 ( .a ({new_AGEMA_signal_3076, new_AGEMA_signal_3075, new_AGEMA_signal_3074, SHIFTROWS[49]}), .b ({new_AGEMA_signal_3508, new_AGEMA_signal_3507, new_AGEMA_signal_3506, SHIFTROWS[81]}), .c ({ROUND_OUT_s3[49], ROUND_OUT_s2[49], ROUND_OUT_s1[49], ROUND_OUT_s0[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U12 ( .a ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, new_AGEMA_signal_3077, SHIFTROWS[52]}), .b ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, new_AGEMA_signal_3383, SHIFTROWS[84]}), .c ({ROUND_OUT_s3[52], ROUND_OUT_s2[52], ROUND_OUT_s1[52], ROUND_OUT_s0[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U7 ( .a ({new_AGEMA_signal_3082, new_AGEMA_signal_3081, new_AGEMA_signal_3080, SHIFTROWS[57]}), .b ({new_AGEMA_signal_3406, new_AGEMA_signal_3405, new_AGEMA_signal_3404, SHIFTROWS[89]}), .c ({ROUND_OUT_s3[57], ROUND_OUT_s2[57], ROUND_OUT_s1[57], ROUND_OUT_s0[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U4 ( .a ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, new_AGEMA_signal_3083, SHIFTROWS[60]}), .b ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, new_AGEMA_signal_3401, SHIFTROWS[92]}), .c ({ROUND_OUT_s3[60], ROUND_OUT_s2[60], ROUND_OUT_s1[60], ROUND_OUT_s0[60]}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U410 ( .a ({ROUND_KEY_s3[352], ROUND_KEY_s2[352], ROUND_KEY_s1[352], ROUND_KEY_s0[352]}), .b ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, new_AGEMA_signal_3464, CONST_ADDITION[96]}), .c ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, new_AGEMA_signal_3503, n411}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U411 ( .a ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, new_AGEMA_signal_1115, n412}), .b ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, new_AGEMA_signal_3503, n411}), .c ({ROUND_OUT_s3[64], ROUND_OUT_s2[64], ROUND_OUT_s1[64], ROUND_OUT_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U435 ( .a ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, new_AGEMA_signal_3461, SUBSTITUTION_88}), .b ({ROUND_KEY_s3[344], ROUND_KEY_s2[344], ROUND_KEY_s1[344], ROUND_KEY_s0[344]}), .c ({new_AGEMA_signal_3514, new_AGEMA_signal_3513, new_AGEMA_signal_3512, n428}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U436 ( .a ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, new_AGEMA_signal_1187, n429}), .b ({new_AGEMA_signal_3514, new_AGEMA_signal_3513, new_AGEMA_signal_3512, n428}), .c ({new_AGEMA_signal_3604, new_AGEMA_signal_3603, new_AGEMA_signal_3602, n430}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U437 ( .a ({1'b0, 1'b0, 1'b0, CONST_IN[4]}), .b ({new_AGEMA_signal_3604, new_AGEMA_signal_3603, new_AGEMA_signal_3602, n430}), .c ({new_AGEMA_signal_3652, new_AGEMA_signal_3651, new_AGEMA_signal_3650, SHIFTROWS[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U460 ( .a ({ROUND_KEY_s3[336], ROUND_KEY_s2[336], ROUND_KEY_s1[336], ROUND_KEY_s0[336]}), .b ({new_AGEMA_signal_3460, new_AGEMA_signal_3459, new_AGEMA_signal_3458, CONST_ADDITION[80]}), .c ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_3518, n445}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U461 ( .a ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, new_AGEMA_signal_1259, n446}), .b ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_3518, n445}), .c ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, new_AGEMA_signal_3605, SHIFTROWS[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U484 ( .a ({ROUND_KEY_s3[328], ROUND_KEY_s2[328], ROUND_KEY_s1[328], ROUND_KEY_s0[328]}), .b ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, new_AGEMA_signal_3455, CONST_ADDITION[72]}), .c ({new_AGEMA_signal_3526, new_AGEMA_signal_3525, new_AGEMA_signal_3524, n461}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U485 ( .a ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, new_AGEMA_signal_1331, n462}), .b ({new_AGEMA_signal_3526, new_AGEMA_signal_3525, new_AGEMA_signal_3524, n461}), .c ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, new_AGEMA_signal_3608, SHIFTROWS[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U508 ( .a ({ROUND_KEY_s3[320], ROUND_KEY_s2[320], ROUND_KEY_s1[320], ROUND_KEY_s0[320]}), .b ({new_AGEMA_signal_3454, new_AGEMA_signal_3453, new_AGEMA_signal_3452, CONST_ADDITION[64]}), .c ({new_AGEMA_signal_3532, new_AGEMA_signal_3531, new_AGEMA_signal_3530, n477}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U509 ( .a ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, new_AGEMA_signal_1403, n478}), .b ({new_AGEMA_signal_3532, new_AGEMA_signal_3531, new_AGEMA_signal_3530, n477}), .c ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, new_AGEMA_signal_3611, SHIFTROWS[88]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U535 ( .a ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, new_AGEMA_signal_3473, SUBSTITUTION[120]}), .b ({ROUND_KEY_s3[376], ROUND_KEY_s2[376], ROUND_KEY_s1[376], ROUND_KEY_s0[376]}), .c ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, new_AGEMA_signal_3539, n496}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U536 ( .a ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, new_AGEMA_signal_1475, n497}), .b ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, new_AGEMA_signal_3539, n496}), .c ({new_AGEMA_signal_3616, new_AGEMA_signal_3615, new_AGEMA_signal_3614, n498}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U537 ( .a ({1'b0, 1'b0, 1'b0, CONST_IN[0]}), .b ({new_AGEMA_signal_3616, new_AGEMA_signal_3615, new_AGEMA_signal_3614, n498}), .c ({ROUND_OUT_s3[88], ROUND_OUT_s2[88], ROUND_OUT_s1[88], ROUND_OUT_s0[88]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U560 ( .a ({ROUND_KEY_s3[368], ROUND_KEY_s2[368], ROUND_KEY_s1[368], ROUND_KEY_s0[368]}), .b ({new_AGEMA_signal_3472, new_AGEMA_signal_3471, new_AGEMA_signal_3470, CONST_ADDITION[112]}), .c ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, new_AGEMA_signal_3545, n513}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U561 ( .a ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, new_AGEMA_signal_1547, n514}), .b ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, new_AGEMA_signal_3545, n513}), .c ({ROUND_OUT_s3[80], ROUND_OUT_s2[80], ROUND_OUT_s1[80], ROUND_OUT_s0[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U584 ( .a ({ROUND_KEY_s3[360], ROUND_KEY_s2[360], ROUND_KEY_s1[360], ROUND_KEY_s0[360]}), .b ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, new_AGEMA_signal_3467, CONST_ADDITION[104]}), .c ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, new_AGEMA_signal_3551, n529}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) U585 ( .a ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, new_AGEMA_signal_1619, n530}), .b ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, new_AGEMA_signal_3551, n529}), .c ({ROUND_OUT_s3[72], ROUND_OUT_s2[72], ROUND_OUT_s1[72], ROUND_OUT_s0[72]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_0_U8 ( .a ({new_AGEMA_signal_3286, new_AGEMA_signal_3285, new_AGEMA_signal_3284, S_0_R2[3]}), .b ({ROUND_IN_s3[2], ROUND_IN_s2[2], ROUND_IN_s1[2], ROUND_IN_s0[2]}), .c ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, new_AGEMA_signal_3428, SHIFTROWS[8]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_0_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3052, new_AGEMA_signal_3051, new_AGEMA_signal_3050, SHIFTROWS[9]}), .b ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, new_AGEMA_signal_2594, SHIFTROWS[11]}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_3286, new_AGEMA_signal_3285, new_AGEMA_signal_3284, S_0_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_1_U8 ( .a ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, new_AGEMA_signal_3287, S_1_R2[3]}), .b ({ROUND_IN_s3[10], ROUND_IN_s2[10], ROUND_IN_s1[10], ROUND_IN_s0[10]}), .c ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, new_AGEMA_signal_3431, SHIFTROWS[16]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_1_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3058, new_AGEMA_signal_3057, new_AGEMA_signal_3056, SHIFTROWS[17]}), .b ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, new_AGEMA_signal_2603, SHIFTROWS[19]}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, new_AGEMA_signal_3287, S_1_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_2_U8 ( .a ({new_AGEMA_signal_3292, new_AGEMA_signal_3291, new_AGEMA_signal_3290, S_2_R2[3]}), .b ({ROUND_IN_s3[18], ROUND_IN_s2[18], ROUND_IN_s1[18], ROUND_IN_s0[18]}), .c ({new_AGEMA_signal_3436, new_AGEMA_signal_3435, new_AGEMA_signal_3434, SHIFTROWS[24]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_2_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3064, new_AGEMA_signal_3063, new_AGEMA_signal_3062, SHIFTROWS[25]}), .b ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, new_AGEMA_signal_2612, SHIFTROWS[27]}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_3292, new_AGEMA_signal_3291, new_AGEMA_signal_3290, S_2_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_3_U8 ( .a ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, new_AGEMA_signal_3293, S_3_R2[3]}), .b ({ROUND_IN_s3[26], ROUND_IN_s2[26], ROUND_IN_s1[26], ROUND_IN_s0[26]}), .c ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, new_AGEMA_signal_3437, SHIFTROWS[0]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_3_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3070, new_AGEMA_signal_3069, new_AGEMA_signal_3068, SHIFTROWS[1]}), .b ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, new_AGEMA_signal_2621, SHIFTROWS[3]}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, new_AGEMA_signal_3293, S_3_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_4_U8 ( .a ({new_AGEMA_signal_3298, new_AGEMA_signal_3297, new_AGEMA_signal_3296, S_4_R2[3]}), .b ({ROUND_IN_s3[34], ROUND_IN_s2[34], ROUND_IN_s1[34], ROUND_IN_s0[34]}), .c ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, new_AGEMA_signal_3440, SHIFTROWS[48]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_4_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3076, new_AGEMA_signal_3075, new_AGEMA_signal_3074, SHIFTROWS[49]}), .b ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, new_AGEMA_signal_2630, SHIFTROWS[51]}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_3298, new_AGEMA_signal_3297, new_AGEMA_signal_3296, S_4_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_5_U8 ( .a ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, new_AGEMA_signal_3299, S_5_R2[3]}), .b ({ROUND_IN_s3[42], ROUND_IN_s2[42], ROUND_IN_s1[42], ROUND_IN_s0[42]}), .c ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, new_AGEMA_signal_3443, SHIFTROWS[56]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_5_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3082, new_AGEMA_signal_3081, new_AGEMA_signal_3080, SHIFTROWS[57]}), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, new_AGEMA_signal_2639, SHIFTROWS[59]}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, new_AGEMA_signal_3299, S_5_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_6_U8 ( .a ({new_AGEMA_signal_3304, new_AGEMA_signal_3303, new_AGEMA_signal_3302, S_6_R2[3]}), .b ({ROUND_IN_s3[50], ROUND_IN_s2[50], ROUND_IN_s1[50], ROUND_IN_s0[50]}), .c ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, SHIFTROWS[32]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_6_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3088, new_AGEMA_signal_3087, new_AGEMA_signal_3086, SHIFTROWS[33]}), .b ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, new_AGEMA_signal_2648, SHIFTROWS[35]}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_3304, new_AGEMA_signal_3303, new_AGEMA_signal_3302, S_6_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_7_U8 ( .a ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, new_AGEMA_signal_3305, S_7_R2[3]}), .b ({ROUND_IN_s3[58], ROUND_IN_s2[58], ROUND_IN_s1[58], ROUND_IN_s0[58]}), .c ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, new_AGEMA_signal_3449, SHIFTROWS[40]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_7_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3094, new_AGEMA_signal_3093, new_AGEMA_signal_3092, SUBSTITUTION_57}), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, new_AGEMA_signal_2657, SHIFTROWS[43]}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, new_AGEMA_signal_3305, S_7_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_8_U8 ( .a ({new_AGEMA_signal_3310, new_AGEMA_signal_3309, new_AGEMA_signal_3308, S_8_R2[3]}), .b ({ROUND_IN_s3[66], ROUND_IN_s2[66], ROUND_IN_s1[66], ROUND_IN_s0[66]}), .c ({new_AGEMA_signal_3454, new_AGEMA_signal_3453, new_AGEMA_signal_3452, CONST_ADDITION[64]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_8_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3100, new_AGEMA_signal_3099, new_AGEMA_signal_3098, CONST_ADDITION[65]}), .b ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, new_AGEMA_signal_2666, CONST_ADDITION[67]}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_3310, new_AGEMA_signal_3309, new_AGEMA_signal_3308, S_8_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_9_U8 ( .a ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, new_AGEMA_signal_3311, S_9_R2[3]}), .b ({ROUND_IN_s3[74], ROUND_IN_s2[74], ROUND_IN_s1[74], ROUND_IN_s0[74]}), .c ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, new_AGEMA_signal_3455, CONST_ADDITION[72]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_9_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3106, new_AGEMA_signal_3105, new_AGEMA_signal_3104, CONST_ADDITION[73]}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, new_AGEMA_signal_2675, CONST_ADDITION[75]}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, new_AGEMA_signal_3311, S_9_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_10_U8 ( .a ({new_AGEMA_signal_3316, new_AGEMA_signal_3315, new_AGEMA_signal_3314, S_10_R2[3]}), .b ({ROUND_IN_s3[82], ROUND_IN_s2[82], ROUND_IN_s1[82], ROUND_IN_s0[82]}), .c ({new_AGEMA_signal_3460, new_AGEMA_signal_3459, new_AGEMA_signal_3458, CONST_ADDITION[80]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_10_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3112, new_AGEMA_signal_3111, new_AGEMA_signal_3110, CONST_ADDITION[81]}), .b ({new_AGEMA_signal_2686, new_AGEMA_signal_2685, new_AGEMA_signal_2684, CONST_ADDITION[83]}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_3316, new_AGEMA_signal_3315, new_AGEMA_signal_3314, S_10_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_11_U8 ( .a ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, new_AGEMA_signal_3317, S_11_R2[3]}), .b ({ROUND_IN_s3[90], ROUND_IN_s2[90], ROUND_IN_s1[90], ROUND_IN_s0[90]}), .c ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, new_AGEMA_signal_3461, SUBSTITUTION_88}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_11_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3118, new_AGEMA_signal_3117, new_AGEMA_signal_3116, SUBSTITUTION_89}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, new_AGEMA_signal_2693, CONST_ADDITION[91]}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, new_AGEMA_signal_3317, S_11_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_12_U8 ( .a ({new_AGEMA_signal_3322, new_AGEMA_signal_3321, new_AGEMA_signal_3320, S_12_R2[3]}), .b ({ROUND_IN_s3[98], ROUND_IN_s2[98], ROUND_IN_s1[98], ROUND_IN_s0[98]}), .c ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, new_AGEMA_signal_3464, CONST_ADDITION[96]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_12_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3124, new_AGEMA_signal_3123, new_AGEMA_signal_3122, CONST_ADDITION[97]}), .b ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, CONST_ADDITION[99]}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_3322, new_AGEMA_signal_3321, new_AGEMA_signal_3320, S_12_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_13_U8 ( .a ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, new_AGEMA_signal_3323, S_13_R2[3]}), .b ({ROUND_IN_s3[106], ROUND_IN_s2[106], ROUND_IN_s1[106], ROUND_IN_s0[106]}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, new_AGEMA_signal_3467, CONST_ADDITION[104]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_13_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3130, new_AGEMA_signal_3129, new_AGEMA_signal_3128, CONST_ADDITION[105]}), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, new_AGEMA_signal_2711, CONST_ADDITION[107]}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, new_AGEMA_signal_3323, S_13_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_14_U8 ( .a ({new_AGEMA_signal_3328, new_AGEMA_signal_3327, new_AGEMA_signal_3326, S_14_R2[3]}), .b ({ROUND_IN_s3[114], ROUND_IN_s2[114], ROUND_IN_s1[114], ROUND_IN_s0[114]}), .c ({new_AGEMA_signal_3472, new_AGEMA_signal_3471, new_AGEMA_signal_3470, CONST_ADDITION[112]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_14_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3136, new_AGEMA_signal_3135, new_AGEMA_signal_3134, CONST_ADDITION[113]}), .b ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, CONST_ADDITION[115]}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_3328, new_AGEMA_signal_3327, new_AGEMA_signal_3326, S_14_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) S_15_U8 ( .a ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, new_AGEMA_signal_3329, S_15_R2[3]}), .b ({ROUND_IN_s3[122], ROUND_IN_s2[122], ROUND_IN_s1[122], ROUND_IN_s0[122]}), .c ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, new_AGEMA_signal_3473, SUBSTITUTION[120]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) S_15_NOR2Inst_3_U1 ( .a ({new_AGEMA_signal_3142, new_AGEMA_signal_3141, new_AGEMA_signal_3140, SUBSTITUTION[121]}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, new_AGEMA_signal_2729, SUBSTITUTION[123]}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, new_AGEMA_signal_3329, S_15_R2[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U94 ( .a ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, new_AGEMA_signal_3437, SHIFTROWS[0]}), .b ({ROUND_OUT_s3[0], ROUND_OUT_s2[0], ROUND_OUT_s1[0], ROUND_OUT_s0[0]}), .c ({ROUND_OUT_s3[96], ROUND_OUT_s2[96], ROUND_OUT_s1[96], ROUND_OUT_s0[96]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U93 ( .a ({ROUND_OUT_s3[64], ROUND_OUT_s2[64], ROUND_OUT_s1[64], ROUND_OUT_s0[64]}), .b ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, SHIFTROWS[32]}), .c ({ROUND_OUT_s3[0], ROUND_OUT_s2[0], ROUND_OUT_s1[0], ROUND_OUT_s0[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U88 ( .a ({new_AGEMA_signal_3436, new_AGEMA_signal_3435, new_AGEMA_signal_3434, SHIFTROWS[24]}), .b ({ROUND_OUT_s3[24], ROUND_OUT_s2[24], ROUND_OUT_s1[24], ROUND_OUT_s0[24]}), .c ({ROUND_OUT_s3[120], ROUND_OUT_s2[120], ROUND_OUT_s1[120], ROUND_OUT_s0[120]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U87 ( .a ({ROUND_OUT_s3[88], ROUND_OUT_s2[88], ROUND_OUT_s1[88], ROUND_OUT_s0[88]}), .b ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, new_AGEMA_signal_3443, SHIFTROWS[56]}), .c ({ROUND_OUT_s3[24], ROUND_OUT_s2[24], ROUND_OUT_s1[24], ROUND_OUT_s0[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U86 ( .a ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, new_AGEMA_signal_3431, SHIFTROWS[16]}), .b ({ROUND_OUT_s3[16], ROUND_OUT_s2[16], ROUND_OUT_s1[16], ROUND_OUT_s0[16]}), .c ({ROUND_OUT_s3[112], ROUND_OUT_s2[112], ROUND_OUT_s1[112], ROUND_OUT_s0[112]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U85 ( .a ({ROUND_OUT_s3[80], ROUND_OUT_s2[80], ROUND_OUT_s1[80], ROUND_OUT_s0[80]}), .b ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, new_AGEMA_signal_3440, SHIFTROWS[48]}), .c ({ROUND_OUT_s3[16], ROUND_OUT_s2[16], ROUND_OUT_s1[16], ROUND_OUT_s0[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U56 ( .a ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, new_AGEMA_signal_3428, SHIFTROWS[8]}), .b ({ROUND_OUT_s3[8], ROUND_OUT_s2[8], ROUND_OUT_s1[8], ROUND_OUT_s0[8]}), .c ({ROUND_OUT_s3[104], ROUND_OUT_s2[104], ROUND_OUT_s1[104], ROUND_OUT_s0[104]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U55 ( .a ({ROUND_OUT_s3[72], ROUND_OUT_s2[72], ROUND_OUT_s1[72], ROUND_OUT_s0[72]}), .b ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, new_AGEMA_signal_3449, SHIFTROWS[40]}), .c ({ROUND_OUT_s3[8], ROUND_OUT_s2[8], ROUND_OUT_s1[8], ROUND_OUT_s0[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U32 ( .a ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, SHIFTROWS[32]}), .b ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, new_AGEMA_signal_3608, SHIFTROWS[64]}), .c ({ROUND_OUT_s3[32], ROUND_OUT_s2[32], ROUND_OUT_s1[32], ROUND_OUT_s0[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U24 ( .a ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, new_AGEMA_signal_3449, SHIFTROWS[40]}), .b ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, new_AGEMA_signal_3605, SHIFTROWS[72]}), .c ({ROUND_OUT_s3[40], ROUND_OUT_s2[40], ROUND_OUT_s1[40], ROUND_OUT_s0[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U16 ( .a ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, new_AGEMA_signal_3440, SHIFTROWS[48]}), .b ({new_AGEMA_signal_3652, new_AGEMA_signal_3651, new_AGEMA_signal_3650, SHIFTROWS[80]}), .c ({ROUND_OUT_s3[48], ROUND_OUT_s2[48], ROUND_OUT_s1[48], ROUND_OUT_s0[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MC_U8 ( .a ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, new_AGEMA_signal_3443, SHIFTROWS[56]}), .b ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, new_AGEMA_signal_3611, SHIFTROWS[88]}), .c ({ROUND_OUT_s3[56], ROUND_OUT_s2[56], ROUND_OUT_s1[56], ROUND_OUT_s0[56]}) ) ;

endmodule
