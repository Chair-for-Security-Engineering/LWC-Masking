/* modified netlist. Source: module SubCells in file ./test/SubCells.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module SubCells_HPC2_ClockGating_d1 (SubC_in_s0, clk, SubC_in_s1, Fresh, /*rst,*/ SubC_out_s0, SubC_out_s1/*, Synch*/);
    input [127:0] SubC_in_s0 ;
    input clk ;
    input [127:0] SubC_in_s1 ;
    //input rst ;
    input [191:0] Fresh ;
    output [127:0] SubC_out_s0 ;
    output [127:0] SubC_out_s1 ;
    //output Synch ;
    wire SB_31_n15 ;
    wire SB_31_n14 ;
    wire SB_31_n13 ;
    wire SB_31_n12 ;
    wire SB_31_n11 ;
    wire SB_31_n10 ;
    wire SB_31_n9 ;
    wire SB_31_T5 ;
    wire SB_31_T4 ;
    wire SB_31_T3 ;
    wire SB_31_T2 ;
    wire SB_31_T1 ;
    wire SB_31_T0 ;
    wire SB_30_n15 ;
    wire SB_30_n14 ;
    wire SB_30_n13 ;
    wire SB_30_n12 ;
    wire SB_30_n11 ;
    wire SB_30_n10 ;
    wire SB_30_n9 ;
    wire SB_30_T5 ;
    wire SB_30_T4 ;
    wire SB_30_T3 ;
    wire SB_30_T2 ;
    wire SB_30_T1 ;
    wire SB_30_T0 ;
    wire SB_29_n15 ;
    wire SB_29_n14 ;
    wire SB_29_n13 ;
    wire SB_29_n12 ;
    wire SB_29_n11 ;
    wire SB_29_n10 ;
    wire SB_29_n9 ;
    wire SB_29_T5 ;
    wire SB_29_T4 ;
    wire SB_29_T3 ;
    wire SB_29_T2 ;
    wire SB_29_T1 ;
    wire SB_29_T0 ;
    wire SB_28_n15 ;
    wire SB_28_n14 ;
    wire SB_28_n13 ;
    wire SB_28_n12 ;
    wire SB_28_n11 ;
    wire SB_28_n10 ;
    wire SB_28_n9 ;
    wire SB_28_T5 ;
    wire SB_28_T4 ;
    wire SB_28_T3 ;
    wire SB_28_T2 ;
    wire SB_28_T1 ;
    wire SB_28_T0 ;
    wire SB_27_n15 ;
    wire SB_27_n14 ;
    wire SB_27_n13 ;
    wire SB_27_n12 ;
    wire SB_27_n11 ;
    wire SB_27_n10 ;
    wire SB_27_n9 ;
    wire SB_27_T5 ;
    wire SB_27_T4 ;
    wire SB_27_T3 ;
    wire SB_27_T2 ;
    wire SB_27_T1 ;
    wire SB_27_T0 ;
    wire SB_26_n15 ;
    wire SB_26_n14 ;
    wire SB_26_n13 ;
    wire SB_26_n12 ;
    wire SB_26_n11 ;
    wire SB_26_n10 ;
    wire SB_26_n9 ;
    wire SB_26_T5 ;
    wire SB_26_T4 ;
    wire SB_26_T3 ;
    wire SB_26_T2 ;
    wire SB_26_T1 ;
    wire SB_26_T0 ;
    wire SB_25_n15 ;
    wire SB_25_n14 ;
    wire SB_25_n13 ;
    wire SB_25_n12 ;
    wire SB_25_n11 ;
    wire SB_25_n10 ;
    wire SB_25_n9 ;
    wire SB_25_T5 ;
    wire SB_25_T4 ;
    wire SB_25_T3 ;
    wire SB_25_T2 ;
    wire SB_25_T1 ;
    wire SB_25_T0 ;
    wire SB_24_n15 ;
    wire SB_24_n14 ;
    wire SB_24_n13 ;
    wire SB_24_n12 ;
    wire SB_24_n11 ;
    wire SB_24_n10 ;
    wire SB_24_n9 ;
    wire SB_24_T5 ;
    wire SB_24_T4 ;
    wire SB_24_T3 ;
    wire SB_24_T2 ;
    wire SB_24_T1 ;
    wire SB_24_T0 ;
    wire SB_23_n15 ;
    wire SB_23_n14 ;
    wire SB_23_n13 ;
    wire SB_23_n12 ;
    wire SB_23_n11 ;
    wire SB_23_n10 ;
    wire SB_23_n9 ;
    wire SB_23_T5 ;
    wire SB_23_T4 ;
    wire SB_23_T3 ;
    wire SB_23_T2 ;
    wire SB_23_T1 ;
    wire SB_23_T0 ;
    wire SB_22_n15 ;
    wire SB_22_n14 ;
    wire SB_22_n13 ;
    wire SB_22_n12 ;
    wire SB_22_n11 ;
    wire SB_22_n10 ;
    wire SB_22_n9 ;
    wire SB_22_T5 ;
    wire SB_22_T4 ;
    wire SB_22_T3 ;
    wire SB_22_T2 ;
    wire SB_22_T1 ;
    wire SB_22_T0 ;
    wire SB_21_n15 ;
    wire SB_21_n14 ;
    wire SB_21_n13 ;
    wire SB_21_n12 ;
    wire SB_21_n11 ;
    wire SB_21_n10 ;
    wire SB_21_n9 ;
    wire SB_21_T5 ;
    wire SB_21_T4 ;
    wire SB_21_T3 ;
    wire SB_21_T2 ;
    wire SB_21_T1 ;
    wire SB_21_T0 ;
    wire SB_20_n15 ;
    wire SB_20_n14 ;
    wire SB_20_n13 ;
    wire SB_20_n12 ;
    wire SB_20_n11 ;
    wire SB_20_n10 ;
    wire SB_20_n9 ;
    wire SB_20_T5 ;
    wire SB_20_T4 ;
    wire SB_20_T3 ;
    wire SB_20_T2 ;
    wire SB_20_T1 ;
    wire SB_20_T0 ;
    wire SB_19_n15 ;
    wire SB_19_n14 ;
    wire SB_19_n13 ;
    wire SB_19_n12 ;
    wire SB_19_n11 ;
    wire SB_19_n10 ;
    wire SB_19_n9 ;
    wire SB_19_T5 ;
    wire SB_19_T4 ;
    wire SB_19_T3 ;
    wire SB_19_T2 ;
    wire SB_19_T1 ;
    wire SB_19_T0 ;
    wire SB_18_n15 ;
    wire SB_18_n14 ;
    wire SB_18_n13 ;
    wire SB_18_n12 ;
    wire SB_18_n11 ;
    wire SB_18_n10 ;
    wire SB_18_n9 ;
    wire SB_18_T5 ;
    wire SB_18_T4 ;
    wire SB_18_T3 ;
    wire SB_18_T2 ;
    wire SB_18_T1 ;
    wire SB_18_T0 ;
    wire SB_17_n15 ;
    wire SB_17_n14 ;
    wire SB_17_n13 ;
    wire SB_17_n12 ;
    wire SB_17_n11 ;
    wire SB_17_n10 ;
    wire SB_17_n9 ;
    wire SB_17_T5 ;
    wire SB_17_T4 ;
    wire SB_17_T3 ;
    wire SB_17_T2 ;
    wire SB_17_T1 ;
    wire SB_17_T0 ;
    wire SB_16_n15 ;
    wire SB_16_n14 ;
    wire SB_16_n13 ;
    wire SB_16_n12 ;
    wire SB_16_n11 ;
    wire SB_16_n10 ;
    wire SB_16_n9 ;
    wire SB_16_T5 ;
    wire SB_16_T4 ;
    wire SB_16_T3 ;
    wire SB_16_T2 ;
    wire SB_16_T1 ;
    wire SB_16_T0 ;
    wire SB_15_n15 ;
    wire SB_15_n14 ;
    wire SB_15_n13 ;
    wire SB_15_n12 ;
    wire SB_15_n11 ;
    wire SB_15_n10 ;
    wire SB_15_n9 ;
    wire SB_15_T5 ;
    wire SB_15_T4 ;
    wire SB_15_T3 ;
    wire SB_15_T2 ;
    wire SB_15_T1 ;
    wire SB_15_T0 ;
    wire SB_14_n15 ;
    wire SB_14_n14 ;
    wire SB_14_n13 ;
    wire SB_14_n12 ;
    wire SB_14_n11 ;
    wire SB_14_n10 ;
    wire SB_14_n9 ;
    wire SB_14_T5 ;
    wire SB_14_T4 ;
    wire SB_14_T3 ;
    wire SB_14_T2 ;
    wire SB_14_T1 ;
    wire SB_14_T0 ;
    wire SB_13_n15 ;
    wire SB_13_n14 ;
    wire SB_13_n13 ;
    wire SB_13_n12 ;
    wire SB_13_n11 ;
    wire SB_13_n10 ;
    wire SB_13_n9 ;
    wire SB_13_T5 ;
    wire SB_13_T4 ;
    wire SB_13_T3 ;
    wire SB_13_T2 ;
    wire SB_13_T1 ;
    wire SB_13_T0 ;
    wire SB_12_n15 ;
    wire SB_12_n14 ;
    wire SB_12_n13 ;
    wire SB_12_n12 ;
    wire SB_12_n11 ;
    wire SB_12_n10 ;
    wire SB_12_n9 ;
    wire SB_12_T5 ;
    wire SB_12_T4 ;
    wire SB_12_T3 ;
    wire SB_12_T2 ;
    wire SB_12_T1 ;
    wire SB_12_T0 ;
    wire SB_11_n15 ;
    wire SB_11_n14 ;
    wire SB_11_n13 ;
    wire SB_11_n12 ;
    wire SB_11_n11 ;
    wire SB_11_n10 ;
    wire SB_11_n9 ;
    wire SB_11_T5 ;
    wire SB_11_T4 ;
    wire SB_11_T3 ;
    wire SB_11_T2 ;
    wire SB_11_T1 ;
    wire SB_11_T0 ;
    wire SB_10_n15 ;
    wire SB_10_n14 ;
    wire SB_10_n13 ;
    wire SB_10_n12 ;
    wire SB_10_n11 ;
    wire SB_10_n10 ;
    wire SB_10_n9 ;
    wire SB_10_T5 ;
    wire SB_10_T4 ;
    wire SB_10_T3 ;
    wire SB_10_T2 ;
    wire SB_10_T1 ;
    wire SB_10_T0 ;
    wire SB_9_n15 ;
    wire SB_9_n14 ;
    wire SB_9_n13 ;
    wire SB_9_n12 ;
    wire SB_9_n11 ;
    wire SB_9_n10 ;
    wire SB_9_n9 ;
    wire SB_9_T5 ;
    wire SB_9_T4 ;
    wire SB_9_T3 ;
    wire SB_9_T2 ;
    wire SB_9_T1 ;
    wire SB_9_T0 ;
    wire SB_8_n15 ;
    wire SB_8_n14 ;
    wire SB_8_n13 ;
    wire SB_8_n12 ;
    wire SB_8_n11 ;
    wire SB_8_n10 ;
    wire SB_8_n9 ;
    wire SB_8_T5 ;
    wire SB_8_T4 ;
    wire SB_8_T3 ;
    wire SB_8_T2 ;
    wire SB_8_T1 ;
    wire SB_8_T0 ;
    wire SB_7_n15 ;
    wire SB_7_n14 ;
    wire SB_7_n13 ;
    wire SB_7_n12 ;
    wire SB_7_n11 ;
    wire SB_7_n10 ;
    wire SB_7_n9 ;
    wire SB_7_T5 ;
    wire SB_7_T4 ;
    wire SB_7_T3 ;
    wire SB_7_T2 ;
    wire SB_7_T1 ;
    wire SB_7_T0 ;
    wire SB_6_n15 ;
    wire SB_6_n14 ;
    wire SB_6_n13 ;
    wire SB_6_n12 ;
    wire SB_6_n11 ;
    wire SB_6_n10 ;
    wire SB_6_n9 ;
    wire SB_6_T5 ;
    wire SB_6_T4 ;
    wire SB_6_T3 ;
    wire SB_6_T2 ;
    wire SB_6_T1 ;
    wire SB_6_T0 ;
    wire SB_5_n15 ;
    wire SB_5_n14 ;
    wire SB_5_n13 ;
    wire SB_5_n12 ;
    wire SB_5_n11 ;
    wire SB_5_n10 ;
    wire SB_5_n9 ;
    wire SB_5_T5 ;
    wire SB_5_T4 ;
    wire SB_5_T3 ;
    wire SB_5_T2 ;
    wire SB_5_T1 ;
    wire SB_5_T0 ;
    wire SB_4_n15 ;
    wire SB_4_n14 ;
    wire SB_4_n13 ;
    wire SB_4_n12 ;
    wire SB_4_n11 ;
    wire SB_4_n10 ;
    wire SB_4_n9 ;
    wire SB_4_T5 ;
    wire SB_4_T4 ;
    wire SB_4_T3 ;
    wire SB_4_T2 ;
    wire SB_4_T1 ;
    wire SB_4_T0 ;
    wire SB_3_n15 ;
    wire SB_3_n14 ;
    wire SB_3_n13 ;
    wire SB_3_n12 ;
    wire SB_3_n11 ;
    wire SB_3_n10 ;
    wire SB_3_n9 ;
    wire SB_3_T5 ;
    wire SB_3_T4 ;
    wire SB_3_T3 ;
    wire SB_3_T2 ;
    wire SB_3_T1 ;
    wire SB_3_T0 ;
    wire SB_2_n15 ;
    wire SB_2_n14 ;
    wire SB_2_n13 ;
    wire SB_2_n12 ;
    wire SB_2_n11 ;
    wire SB_2_n10 ;
    wire SB_2_n9 ;
    wire SB_2_T5 ;
    wire SB_2_T4 ;
    wire SB_2_T3 ;
    wire SB_2_T2 ;
    wire SB_2_T1 ;
    wire SB_2_T0 ;
    wire SB_1_n15 ;
    wire SB_1_n14 ;
    wire SB_1_n13 ;
    wire SB_1_n12 ;
    wire SB_1_n11 ;
    wire SB_1_n10 ;
    wire SB_1_n9 ;
    wire SB_1_T5 ;
    wire SB_1_T4 ;
    wire SB_1_T3 ;
    wire SB_1_T2 ;
    wire SB_1_T1 ;
    wire SB_1_T0 ;
    wire SB_0_n15 ;
    wire SB_0_n14 ;
    wire SB_0_n13 ;
    wire SB_0_n12 ;
    wire SB_0_n11 ;
    wire SB_0_n10 ;
    wire SB_0_n9 ;
    wire SB_0_T5 ;
    wire SB_0_T4 ;
    wire SB_0_T3 ;
    wire SB_0_T2 ;
    wire SB_0_T1 ;
    wire SB_0_T0 ;
    wire new_AGEMA_signal_681 ;
    wire new_AGEMA_signal_684 ;
    wire new_AGEMA_signal_685 ;
    wire new_AGEMA_signal_686 ;
    wire new_AGEMA_signal_687 ;
    wire new_AGEMA_signal_688 ;
    wire new_AGEMA_signal_691 ;
    wire new_AGEMA_signal_694 ;
    wire new_AGEMA_signal_695 ;
    wire new_AGEMA_signal_696 ;
    wire new_AGEMA_signal_697 ;
    wire new_AGEMA_signal_698 ;
    wire new_AGEMA_signal_701 ;
    wire new_AGEMA_signal_704 ;
    wire new_AGEMA_signal_705 ;
    wire new_AGEMA_signal_706 ;
    wire new_AGEMA_signal_707 ;
    wire new_AGEMA_signal_708 ;
    wire new_AGEMA_signal_711 ;
    wire new_AGEMA_signal_714 ;
    wire new_AGEMA_signal_715 ;
    wire new_AGEMA_signal_716 ;
    wire new_AGEMA_signal_717 ;
    wire new_AGEMA_signal_718 ;
    wire new_AGEMA_signal_721 ;
    wire new_AGEMA_signal_724 ;
    wire new_AGEMA_signal_725 ;
    wire new_AGEMA_signal_726 ;
    wire new_AGEMA_signal_727 ;
    wire new_AGEMA_signal_728 ;
    wire new_AGEMA_signal_731 ;
    wire new_AGEMA_signal_734 ;
    wire new_AGEMA_signal_735 ;
    wire new_AGEMA_signal_736 ;
    wire new_AGEMA_signal_737 ;
    wire new_AGEMA_signal_738 ;
    wire new_AGEMA_signal_741 ;
    wire new_AGEMA_signal_744 ;
    wire new_AGEMA_signal_745 ;
    wire new_AGEMA_signal_746 ;
    wire new_AGEMA_signal_747 ;
    wire new_AGEMA_signal_748 ;
    wire new_AGEMA_signal_751 ;
    wire new_AGEMA_signal_754 ;
    wire new_AGEMA_signal_755 ;
    wire new_AGEMA_signal_756 ;
    wire new_AGEMA_signal_757 ;
    wire new_AGEMA_signal_758 ;
    wire new_AGEMA_signal_761 ;
    wire new_AGEMA_signal_764 ;
    wire new_AGEMA_signal_765 ;
    wire new_AGEMA_signal_766 ;
    wire new_AGEMA_signal_767 ;
    wire new_AGEMA_signal_768 ;
    wire new_AGEMA_signal_771 ;
    wire new_AGEMA_signal_774 ;
    wire new_AGEMA_signal_775 ;
    wire new_AGEMA_signal_776 ;
    wire new_AGEMA_signal_777 ;
    wire new_AGEMA_signal_778 ;
    wire new_AGEMA_signal_781 ;
    wire new_AGEMA_signal_784 ;
    wire new_AGEMA_signal_785 ;
    wire new_AGEMA_signal_786 ;
    wire new_AGEMA_signal_787 ;
    wire new_AGEMA_signal_788 ;
    wire new_AGEMA_signal_791 ;
    wire new_AGEMA_signal_794 ;
    wire new_AGEMA_signal_795 ;
    wire new_AGEMA_signal_796 ;
    wire new_AGEMA_signal_797 ;
    wire new_AGEMA_signal_798 ;
    wire new_AGEMA_signal_801 ;
    wire new_AGEMA_signal_804 ;
    wire new_AGEMA_signal_805 ;
    wire new_AGEMA_signal_806 ;
    wire new_AGEMA_signal_807 ;
    wire new_AGEMA_signal_808 ;
    wire new_AGEMA_signal_811 ;
    wire new_AGEMA_signal_814 ;
    wire new_AGEMA_signal_815 ;
    wire new_AGEMA_signal_816 ;
    wire new_AGEMA_signal_817 ;
    wire new_AGEMA_signal_818 ;
    wire new_AGEMA_signal_821 ;
    wire new_AGEMA_signal_824 ;
    wire new_AGEMA_signal_825 ;
    wire new_AGEMA_signal_826 ;
    wire new_AGEMA_signal_827 ;
    wire new_AGEMA_signal_828 ;
    wire new_AGEMA_signal_831 ;
    wire new_AGEMA_signal_834 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_836 ;
    wire new_AGEMA_signal_837 ;
    wire new_AGEMA_signal_838 ;
    wire new_AGEMA_signal_841 ;
    wire new_AGEMA_signal_844 ;
    wire new_AGEMA_signal_845 ;
    wire new_AGEMA_signal_846 ;
    wire new_AGEMA_signal_847 ;
    wire new_AGEMA_signal_848 ;
    wire new_AGEMA_signal_851 ;
    wire new_AGEMA_signal_854 ;
    wire new_AGEMA_signal_855 ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_857 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_861 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_868 ;
    wire new_AGEMA_signal_871 ;
    wire new_AGEMA_signal_874 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_878 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_886 ;
    wire new_AGEMA_signal_887 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_896 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_898 ;
    wire new_AGEMA_signal_901 ;
    wire new_AGEMA_signal_904 ;
    wire new_AGEMA_signal_905 ;
    wire new_AGEMA_signal_906 ;
    wire new_AGEMA_signal_907 ;
    wire new_AGEMA_signal_908 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_915 ;
    wire new_AGEMA_signal_916 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_921 ;
    wire new_AGEMA_signal_924 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_928 ;
    wire new_AGEMA_signal_931 ;
    wire new_AGEMA_signal_934 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U8 ( .a ({SubC_in_s1[63], SubC_in_s0[63]}), .b ({SubC_in_s1[95], SubC_in_s0[95]}), .c ({new_AGEMA_signal_681, SB_31_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U3 ( .a ({SubC_in_s1[31], SubC_in_s0[31]}), .b ({SubC_in_s1[127], SubC_in_s0[127]}), .c ({new_AGEMA_signal_684, SB_31_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U8 ( .a ({SubC_in_s1[62], SubC_in_s0[62]}), .b ({SubC_in_s1[94], SubC_in_s0[94]}), .c ({new_AGEMA_signal_691, SB_30_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U3 ( .a ({SubC_in_s1[30], SubC_in_s0[30]}), .b ({SubC_in_s1[126], SubC_in_s0[126]}), .c ({new_AGEMA_signal_694, SB_30_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U8 ( .a ({SubC_in_s1[61], SubC_in_s0[61]}), .b ({SubC_in_s1[93], SubC_in_s0[93]}), .c ({new_AGEMA_signal_701, SB_29_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U3 ( .a ({SubC_in_s1[29], SubC_in_s0[29]}), .b ({SubC_in_s1[125], SubC_in_s0[125]}), .c ({new_AGEMA_signal_704, SB_29_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U8 ( .a ({SubC_in_s1[60], SubC_in_s0[60]}), .b ({SubC_in_s1[92], SubC_in_s0[92]}), .c ({new_AGEMA_signal_711, SB_28_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U3 ( .a ({SubC_in_s1[28], SubC_in_s0[28]}), .b ({SubC_in_s1[124], SubC_in_s0[124]}), .c ({new_AGEMA_signal_714, SB_28_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U8 ( .a ({SubC_in_s1[59], SubC_in_s0[59]}), .b ({SubC_in_s1[91], SubC_in_s0[91]}), .c ({new_AGEMA_signal_721, SB_27_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U3 ( .a ({SubC_in_s1[27], SubC_in_s0[27]}), .b ({SubC_in_s1[123], SubC_in_s0[123]}), .c ({new_AGEMA_signal_724, SB_27_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U8 ( .a ({SubC_in_s1[58], SubC_in_s0[58]}), .b ({SubC_in_s1[90], SubC_in_s0[90]}), .c ({new_AGEMA_signal_731, SB_26_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U3 ( .a ({SubC_in_s1[26], SubC_in_s0[26]}), .b ({SubC_in_s1[122], SubC_in_s0[122]}), .c ({new_AGEMA_signal_734, SB_26_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U8 ( .a ({SubC_in_s1[57], SubC_in_s0[57]}), .b ({SubC_in_s1[89], SubC_in_s0[89]}), .c ({new_AGEMA_signal_741, SB_25_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U3 ( .a ({SubC_in_s1[25], SubC_in_s0[25]}), .b ({SubC_in_s1[121], SubC_in_s0[121]}), .c ({new_AGEMA_signal_744, SB_25_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U8 ( .a ({SubC_in_s1[56], SubC_in_s0[56]}), .b ({SubC_in_s1[88], SubC_in_s0[88]}), .c ({new_AGEMA_signal_751, SB_24_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U3 ( .a ({SubC_in_s1[24], SubC_in_s0[24]}), .b ({SubC_in_s1[120], SubC_in_s0[120]}), .c ({new_AGEMA_signal_754, SB_24_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U8 ( .a ({SubC_in_s1[55], SubC_in_s0[55]}), .b ({SubC_in_s1[87], SubC_in_s0[87]}), .c ({new_AGEMA_signal_761, SB_23_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U3 ( .a ({SubC_in_s1[23], SubC_in_s0[23]}), .b ({SubC_in_s1[119], SubC_in_s0[119]}), .c ({new_AGEMA_signal_764, SB_23_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U8 ( .a ({SubC_in_s1[54], SubC_in_s0[54]}), .b ({SubC_in_s1[86], SubC_in_s0[86]}), .c ({new_AGEMA_signal_771, SB_22_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U3 ( .a ({SubC_in_s1[22], SubC_in_s0[22]}), .b ({SubC_in_s1[118], SubC_in_s0[118]}), .c ({new_AGEMA_signal_774, SB_22_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U8 ( .a ({SubC_in_s1[53], SubC_in_s0[53]}), .b ({SubC_in_s1[85], SubC_in_s0[85]}), .c ({new_AGEMA_signal_781, SB_21_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U3 ( .a ({SubC_in_s1[21], SubC_in_s0[21]}), .b ({SubC_in_s1[117], SubC_in_s0[117]}), .c ({new_AGEMA_signal_784, SB_21_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U8 ( .a ({SubC_in_s1[52], SubC_in_s0[52]}), .b ({SubC_in_s1[84], SubC_in_s0[84]}), .c ({new_AGEMA_signal_791, SB_20_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U3 ( .a ({SubC_in_s1[20], SubC_in_s0[20]}), .b ({SubC_in_s1[116], SubC_in_s0[116]}), .c ({new_AGEMA_signal_794, SB_20_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U8 ( .a ({SubC_in_s1[51], SubC_in_s0[51]}), .b ({SubC_in_s1[83], SubC_in_s0[83]}), .c ({new_AGEMA_signal_801, SB_19_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U3 ( .a ({SubC_in_s1[19], SubC_in_s0[19]}), .b ({SubC_in_s1[115], SubC_in_s0[115]}), .c ({new_AGEMA_signal_804, SB_19_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U8 ( .a ({SubC_in_s1[50], SubC_in_s0[50]}), .b ({SubC_in_s1[82], SubC_in_s0[82]}), .c ({new_AGEMA_signal_811, SB_18_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U3 ( .a ({SubC_in_s1[18], SubC_in_s0[18]}), .b ({SubC_in_s1[114], SubC_in_s0[114]}), .c ({new_AGEMA_signal_814, SB_18_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U8 ( .a ({SubC_in_s1[49], SubC_in_s0[49]}), .b ({SubC_in_s1[81], SubC_in_s0[81]}), .c ({new_AGEMA_signal_821, SB_17_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U3 ( .a ({SubC_in_s1[17], SubC_in_s0[17]}), .b ({SubC_in_s1[113], SubC_in_s0[113]}), .c ({new_AGEMA_signal_824, SB_17_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U8 ( .a ({SubC_in_s1[48], SubC_in_s0[48]}), .b ({SubC_in_s1[80], SubC_in_s0[80]}), .c ({new_AGEMA_signal_831, SB_16_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U3 ( .a ({SubC_in_s1[16], SubC_in_s0[16]}), .b ({SubC_in_s1[112], SubC_in_s0[112]}), .c ({new_AGEMA_signal_834, SB_16_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U8 ( .a ({SubC_in_s1[47], SubC_in_s0[47]}), .b ({SubC_in_s1[79], SubC_in_s0[79]}), .c ({new_AGEMA_signal_841, SB_15_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U3 ( .a ({SubC_in_s1[15], SubC_in_s0[15]}), .b ({SubC_in_s1[111], SubC_in_s0[111]}), .c ({new_AGEMA_signal_844, SB_15_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U8 ( .a ({SubC_in_s1[46], SubC_in_s0[46]}), .b ({SubC_in_s1[78], SubC_in_s0[78]}), .c ({new_AGEMA_signal_851, SB_14_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U3 ( .a ({SubC_in_s1[14], SubC_in_s0[14]}), .b ({SubC_in_s1[110], SubC_in_s0[110]}), .c ({new_AGEMA_signal_854, SB_14_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U8 ( .a ({SubC_in_s1[45], SubC_in_s0[45]}), .b ({SubC_in_s1[77], SubC_in_s0[77]}), .c ({new_AGEMA_signal_861, SB_13_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U3 ( .a ({SubC_in_s1[13], SubC_in_s0[13]}), .b ({SubC_in_s1[109], SubC_in_s0[109]}), .c ({new_AGEMA_signal_864, SB_13_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U8 ( .a ({SubC_in_s1[44], SubC_in_s0[44]}), .b ({SubC_in_s1[76], SubC_in_s0[76]}), .c ({new_AGEMA_signal_871, SB_12_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U3 ( .a ({SubC_in_s1[12], SubC_in_s0[12]}), .b ({SubC_in_s1[108], SubC_in_s0[108]}), .c ({new_AGEMA_signal_874, SB_12_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U8 ( .a ({SubC_in_s1[43], SubC_in_s0[43]}), .b ({SubC_in_s1[75], SubC_in_s0[75]}), .c ({new_AGEMA_signal_881, SB_11_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U3 ( .a ({SubC_in_s1[11], SubC_in_s0[11]}), .b ({SubC_in_s1[107], SubC_in_s0[107]}), .c ({new_AGEMA_signal_884, SB_11_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U8 ( .a ({SubC_in_s1[42], SubC_in_s0[42]}), .b ({SubC_in_s1[74], SubC_in_s0[74]}), .c ({new_AGEMA_signal_891, SB_10_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U3 ( .a ({SubC_in_s1[10], SubC_in_s0[10]}), .b ({SubC_in_s1[106], SubC_in_s0[106]}), .c ({new_AGEMA_signal_894, SB_10_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U8 ( .a ({SubC_in_s1[41], SubC_in_s0[41]}), .b ({SubC_in_s1[73], SubC_in_s0[73]}), .c ({new_AGEMA_signal_901, SB_9_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U3 ( .a ({SubC_in_s1[9], SubC_in_s0[9]}), .b ({SubC_in_s1[105], SubC_in_s0[105]}), .c ({new_AGEMA_signal_904, SB_9_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U8 ( .a ({SubC_in_s1[40], SubC_in_s0[40]}), .b ({SubC_in_s1[72], SubC_in_s0[72]}), .c ({new_AGEMA_signal_911, SB_8_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U3 ( .a ({SubC_in_s1[8], SubC_in_s0[8]}), .b ({SubC_in_s1[104], SubC_in_s0[104]}), .c ({new_AGEMA_signal_914, SB_8_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U8 ( .a ({SubC_in_s1[39], SubC_in_s0[39]}), .b ({SubC_in_s1[71], SubC_in_s0[71]}), .c ({new_AGEMA_signal_921, SB_7_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U3 ( .a ({SubC_in_s1[7], SubC_in_s0[7]}), .b ({SubC_in_s1[103], SubC_in_s0[103]}), .c ({new_AGEMA_signal_924, SB_7_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U8 ( .a ({SubC_in_s1[38], SubC_in_s0[38]}), .b ({SubC_in_s1[70], SubC_in_s0[70]}), .c ({new_AGEMA_signal_931, SB_6_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U3 ( .a ({SubC_in_s1[6], SubC_in_s0[6]}), .b ({SubC_in_s1[102], SubC_in_s0[102]}), .c ({new_AGEMA_signal_934, SB_6_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U8 ( .a ({SubC_in_s1[37], SubC_in_s0[37]}), .b ({SubC_in_s1[69], SubC_in_s0[69]}), .c ({new_AGEMA_signal_941, SB_5_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U3 ( .a ({SubC_in_s1[5], SubC_in_s0[5]}), .b ({SubC_in_s1[101], SubC_in_s0[101]}), .c ({new_AGEMA_signal_944, SB_5_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U8 ( .a ({SubC_in_s1[36], SubC_in_s0[36]}), .b ({SubC_in_s1[68], SubC_in_s0[68]}), .c ({new_AGEMA_signal_951, SB_4_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U3 ( .a ({SubC_in_s1[4], SubC_in_s0[4]}), .b ({SubC_in_s1[100], SubC_in_s0[100]}), .c ({new_AGEMA_signal_954, SB_4_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U8 ( .a ({SubC_in_s1[35], SubC_in_s0[35]}), .b ({SubC_in_s1[67], SubC_in_s0[67]}), .c ({new_AGEMA_signal_961, SB_3_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U3 ( .a ({SubC_in_s1[3], SubC_in_s0[3]}), .b ({SubC_in_s1[99], SubC_in_s0[99]}), .c ({new_AGEMA_signal_964, SB_3_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U8 ( .a ({SubC_in_s1[34], SubC_in_s0[34]}), .b ({SubC_in_s1[66], SubC_in_s0[66]}), .c ({new_AGEMA_signal_971, SB_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U3 ( .a ({SubC_in_s1[2], SubC_in_s0[2]}), .b ({SubC_in_s1[98], SubC_in_s0[98]}), .c ({new_AGEMA_signal_974, SB_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U8 ( .a ({SubC_in_s1[33], SubC_in_s0[33]}), .b ({SubC_in_s1[65], SubC_in_s0[65]}), .c ({new_AGEMA_signal_981, SB_1_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U3 ( .a ({SubC_in_s1[1], SubC_in_s0[1]}), .b ({SubC_in_s1[97], SubC_in_s0[97]}), .c ({new_AGEMA_signal_984, SB_1_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U8 ( .a ({SubC_in_s1[32], SubC_in_s0[32]}), .b ({SubC_in_s1[64], SubC_in_s0[64]}), .c ({new_AGEMA_signal_991, SB_0_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U3 ( .a ({SubC_in_s1[0], SubC_in_s0[0]}), .b ({SubC_in_s1[96], SubC_in_s0[96]}), .c ({new_AGEMA_signal_994, SB_0_n10}) ) ;
    //ClockGatingController #(4) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U11 ( .a ({new_AGEMA_signal_1000, SB_31_n15}), .b ({new_AGEMA_signal_681, SB_31_n14}), .c ({SubC_out_s1[127], SubC_out_s0[127]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U9 ( .a ({new_AGEMA_signal_681, SB_31_n14}), .b ({new_AGEMA_signal_687, SB_31_T2}), .c ({new_AGEMA_signal_999, SB_31_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U6 ( .a ({new_AGEMA_signal_1161, SB_31_n11}), .b ({new_AGEMA_signal_686, SB_31_T1}), .c ({SubC_out_s1[95], SubC_out_s0[95]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U5 ( .a ({new_AGEMA_signal_1000, SB_31_n15}), .b ({SubC_in_s1[63], SubC_in_s0[63]}), .c ({new_AGEMA_signal_1161, SB_31_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U4 ( .a ({new_AGEMA_signal_684, SB_31_n10}), .b ({new_AGEMA_signal_685, SB_31_T0}), .c ({new_AGEMA_signal_1000, SB_31_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U1 ( .a ({SubC_in_s1[127], SubC_in_s0[127]}), .b ({new_AGEMA_signal_688, SB_31_T3}), .c ({new_AGEMA_signal_1001, SB_31_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_31_t0_AND_U1 ( .a ({SubC_in_s1[127], SubC_in_s0[127]}), .b ({SubC_in_s1[95], SubC_in_s0[95]}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_685, SB_31_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_31_t1_AND_U1 ( .a ({SubC_in_s1[127], SubC_in_s0[127]}), .b ({SubC_in_s1[63], SubC_in_s0[63]}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_686, SB_31_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_31_t2_AND_U1 ( .a ({SubC_in_s1[127], SubC_in_s0[127]}), .b ({SubC_in_s1[31], SubC_in_s0[31]}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_687, SB_31_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_31_t3_AND_U1 ( .a ({SubC_in_s1[95], SubC_in_s0[95]}), .b ({SubC_in_s1[31], SubC_in_s0[31]}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_688, SB_31_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U11 ( .a ({new_AGEMA_signal_1005, SB_30_n15}), .b ({new_AGEMA_signal_691, SB_30_n14}), .c ({SubC_out_s1[126], SubC_out_s0[126]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U9 ( .a ({new_AGEMA_signal_691, SB_30_n14}), .b ({new_AGEMA_signal_697, SB_30_T2}), .c ({new_AGEMA_signal_1004, SB_30_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U6 ( .a ({new_AGEMA_signal_1165, SB_30_n11}), .b ({new_AGEMA_signal_696, SB_30_T1}), .c ({SubC_out_s1[94], SubC_out_s0[94]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U5 ( .a ({new_AGEMA_signal_1005, SB_30_n15}), .b ({SubC_in_s1[62], SubC_in_s0[62]}), .c ({new_AGEMA_signal_1165, SB_30_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U4 ( .a ({new_AGEMA_signal_694, SB_30_n10}), .b ({new_AGEMA_signal_695, SB_30_T0}), .c ({new_AGEMA_signal_1005, SB_30_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U1 ( .a ({SubC_in_s1[126], SubC_in_s0[126]}), .b ({new_AGEMA_signal_698, SB_30_T3}), .c ({new_AGEMA_signal_1006, SB_30_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_30_t0_AND_U1 ( .a ({SubC_in_s1[126], SubC_in_s0[126]}), .b ({SubC_in_s1[94], SubC_in_s0[94]}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_695, SB_30_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_30_t1_AND_U1 ( .a ({SubC_in_s1[126], SubC_in_s0[126]}), .b ({SubC_in_s1[62], SubC_in_s0[62]}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_696, SB_30_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_30_t2_AND_U1 ( .a ({SubC_in_s1[126], SubC_in_s0[126]}), .b ({SubC_in_s1[30], SubC_in_s0[30]}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_697, SB_30_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_30_t3_AND_U1 ( .a ({SubC_in_s1[94], SubC_in_s0[94]}), .b ({SubC_in_s1[30], SubC_in_s0[30]}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_698, SB_30_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U11 ( .a ({new_AGEMA_signal_1010, SB_29_n15}), .b ({new_AGEMA_signal_701, SB_29_n14}), .c ({SubC_out_s1[125], SubC_out_s0[125]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U9 ( .a ({new_AGEMA_signal_701, SB_29_n14}), .b ({new_AGEMA_signal_707, SB_29_T2}), .c ({new_AGEMA_signal_1009, SB_29_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U6 ( .a ({new_AGEMA_signal_1169, SB_29_n11}), .b ({new_AGEMA_signal_706, SB_29_T1}), .c ({SubC_out_s1[93], SubC_out_s0[93]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U5 ( .a ({new_AGEMA_signal_1010, SB_29_n15}), .b ({SubC_in_s1[61], SubC_in_s0[61]}), .c ({new_AGEMA_signal_1169, SB_29_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U4 ( .a ({new_AGEMA_signal_704, SB_29_n10}), .b ({new_AGEMA_signal_705, SB_29_T0}), .c ({new_AGEMA_signal_1010, SB_29_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U1 ( .a ({SubC_in_s1[125], SubC_in_s0[125]}), .b ({new_AGEMA_signal_708, SB_29_T3}), .c ({new_AGEMA_signal_1011, SB_29_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_29_t0_AND_U1 ( .a ({SubC_in_s1[125], SubC_in_s0[125]}), .b ({SubC_in_s1[93], SubC_in_s0[93]}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_705, SB_29_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_29_t1_AND_U1 ( .a ({SubC_in_s1[125], SubC_in_s0[125]}), .b ({SubC_in_s1[61], SubC_in_s0[61]}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_706, SB_29_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_29_t2_AND_U1 ( .a ({SubC_in_s1[125], SubC_in_s0[125]}), .b ({SubC_in_s1[29], SubC_in_s0[29]}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_707, SB_29_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_29_t3_AND_U1 ( .a ({SubC_in_s1[93], SubC_in_s0[93]}), .b ({SubC_in_s1[29], SubC_in_s0[29]}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_708, SB_29_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U11 ( .a ({new_AGEMA_signal_1015, SB_28_n15}), .b ({new_AGEMA_signal_711, SB_28_n14}), .c ({SubC_out_s1[124], SubC_out_s0[124]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U9 ( .a ({new_AGEMA_signal_711, SB_28_n14}), .b ({new_AGEMA_signal_717, SB_28_T2}), .c ({new_AGEMA_signal_1014, SB_28_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U6 ( .a ({new_AGEMA_signal_1173, SB_28_n11}), .b ({new_AGEMA_signal_716, SB_28_T1}), .c ({SubC_out_s1[92], SubC_out_s0[92]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U5 ( .a ({new_AGEMA_signal_1015, SB_28_n15}), .b ({SubC_in_s1[60], SubC_in_s0[60]}), .c ({new_AGEMA_signal_1173, SB_28_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U4 ( .a ({new_AGEMA_signal_714, SB_28_n10}), .b ({new_AGEMA_signal_715, SB_28_T0}), .c ({new_AGEMA_signal_1015, SB_28_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U1 ( .a ({SubC_in_s1[124], SubC_in_s0[124]}), .b ({new_AGEMA_signal_718, SB_28_T3}), .c ({new_AGEMA_signal_1016, SB_28_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_28_t0_AND_U1 ( .a ({SubC_in_s1[124], SubC_in_s0[124]}), .b ({SubC_in_s1[92], SubC_in_s0[92]}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_715, SB_28_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_28_t1_AND_U1 ( .a ({SubC_in_s1[124], SubC_in_s0[124]}), .b ({SubC_in_s1[60], SubC_in_s0[60]}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_716, SB_28_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_28_t2_AND_U1 ( .a ({SubC_in_s1[124], SubC_in_s0[124]}), .b ({SubC_in_s1[28], SubC_in_s0[28]}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_717, SB_28_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_28_t3_AND_U1 ( .a ({SubC_in_s1[92], SubC_in_s0[92]}), .b ({SubC_in_s1[28], SubC_in_s0[28]}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_718, SB_28_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U11 ( .a ({new_AGEMA_signal_1020, SB_27_n15}), .b ({new_AGEMA_signal_721, SB_27_n14}), .c ({SubC_out_s1[123], SubC_out_s0[123]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U9 ( .a ({new_AGEMA_signal_721, SB_27_n14}), .b ({new_AGEMA_signal_727, SB_27_T2}), .c ({new_AGEMA_signal_1019, SB_27_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U6 ( .a ({new_AGEMA_signal_1177, SB_27_n11}), .b ({new_AGEMA_signal_726, SB_27_T1}), .c ({SubC_out_s1[91], SubC_out_s0[91]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U5 ( .a ({new_AGEMA_signal_1020, SB_27_n15}), .b ({SubC_in_s1[59], SubC_in_s0[59]}), .c ({new_AGEMA_signal_1177, SB_27_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U4 ( .a ({new_AGEMA_signal_724, SB_27_n10}), .b ({new_AGEMA_signal_725, SB_27_T0}), .c ({new_AGEMA_signal_1020, SB_27_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U1 ( .a ({SubC_in_s1[123], SubC_in_s0[123]}), .b ({new_AGEMA_signal_728, SB_27_T3}), .c ({new_AGEMA_signal_1021, SB_27_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_27_t0_AND_U1 ( .a ({SubC_in_s1[123], SubC_in_s0[123]}), .b ({SubC_in_s1[91], SubC_in_s0[91]}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_725, SB_27_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_27_t1_AND_U1 ( .a ({SubC_in_s1[123], SubC_in_s0[123]}), .b ({SubC_in_s1[59], SubC_in_s0[59]}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_726, SB_27_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_27_t2_AND_U1 ( .a ({SubC_in_s1[123], SubC_in_s0[123]}), .b ({SubC_in_s1[27], SubC_in_s0[27]}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_727, SB_27_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_27_t3_AND_U1 ( .a ({SubC_in_s1[91], SubC_in_s0[91]}), .b ({SubC_in_s1[27], SubC_in_s0[27]}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_728, SB_27_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U11 ( .a ({new_AGEMA_signal_1025, SB_26_n15}), .b ({new_AGEMA_signal_731, SB_26_n14}), .c ({SubC_out_s1[122], SubC_out_s0[122]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U9 ( .a ({new_AGEMA_signal_731, SB_26_n14}), .b ({new_AGEMA_signal_737, SB_26_T2}), .c ({new_AGEMA_signal_1024, SB_26_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U6 ( .a ({new_AGEMA_signal_1181, SB_26_n11}), .b ({new_AGEMA_signal_736, SB_26_T1}), .c ({SubC_out_s1[90], SubC_out_s0[90]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U5 ( .a ({new_AGEMA_signal_1025, SB_26_n15}), .b ({SubC_in_s1[58], SubC_in_s0[58]}), .c ({new_AGEMA_signal_1181, SB_26_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U4 ( .a ({new_AGEMA_signal_734, SB_26_n10}), .b ({new_AGEMA_signal_735, SB_26_T0}), .c ({new_AGEMA_signal_1025, SB_26_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U1 ( .a ({SubC_in_s1[122], SubC_in_s0[122]}), .b ({new_AGEMA_signal_738, SB_26_T3}), .c ({new_AGEMA_signal_1026, SB_26_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_26_t0_AND_U1 ( .a ({SubC_in_s1[122], SubC_in_s0[122]}), .b ({SubC_in_s1[90], SubC_in_s0[90]}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_735, SB_26_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_26_t1_AND_U1 ( .a ({SubC_in_s1[122], SubC_in_s0[122]}), .b ({SubC_in_s1[58], SubC_in_s0[58]}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_736, SB_26_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_26_t2_AND_U1 ( .a ({SubC_in_s1[122], SubC_in_s0[122]}), .b ({SubC_in_s1[26], SubC_in_s0[26]}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_737, SB_26_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_26_t3_AND_U1 ( .a ({SubC_in_s1[90], SubC_in_s0[90]}), .b ({SubC_in_s1[26], SubC_in_s0[26]}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_738, SB_26_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U11 ( .a ({new_AGEMA_signal_1030, SB_25_n15}), .b ({new_AGEMA_signal_741, SB_25_n14}), .c ({SubC_out_s1[121], SubC_out_s0[121]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U9 ( .a ({new_AGEMA_signal_741, SB_25_n14}), .b ({new_AGEMA_signal_747, SB_25_T2}), .c ({new_AGEMA_signal_1029, SB_25_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U6 ( .a ({new_AGEMA_signal_1185, SB_25_n11}), .b ({new_AGEMA_signal_746, SB_25_T1}), .c ({SubC_out_s1[89], SubC_out_s0[89]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U5 ( .a ({new_AGEMA_signal_1030, SB_25_n15}), .b ({SubC_in_s1[57], SubC_in_s0[57]}), .c ({new_AGEMA_signal_1185, SB_25_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U4 ( .a ({new_AGEMA_signal_744, SB_25_n10}), .b ({new_AGEMA_signal_745, SB_25_T0}), .c ({new_AGEMA_signal_1030, SB_25_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U1 ( .a ({SubC_in_s1[121], SubC_in_s0[121]}), .b ({new_AGEMA_signal_748, SB_25_T3}), .c ({new_AGEMA_signal_1031, SB_25_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_25_t0_AND_U1 ( .a ({SubC_in_s1[121], SubC_in_s0[121]}), .b ({SubC_in_s1[89], SubC_in_s0[89]}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_745, SB_25_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_25_t1_AND_U1 ( .a ({SubC_in_s1[121], SubC_in_s0[121]}), .b ({SubC_in_s1[57], SubC_in_s0[57]}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_746, SB_25_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_25_t2_AND_U1 ( .a ({SubC_in_s1[121], SubC_in_s0[121]}), .b ({SubC_in_s1[25], SubC_in_s0[25]}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_747, SB_25_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_25_t3_AND_U1 ( .a ({SubC_in_s1[89], SubC_in_s0[89]}), .b ({SubC_in_s1[25], SubC_in_s0[25]}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_748, SB_25_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U11 ( .a ({new_AGEMA_signal_1035, SB_24_n15}), .b ({new_AGEMA_signal_751, SB_24_n14}), .c ({SubC_out_s1[120], SubC_out_s0[120]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U9 ( .a ({new_AGEMA_signal_751, SB_24_n14}), .b ({new_AGEMA_signal_757, SB_24_T2}), .c ({new_AGEMA_signal_1034, SB_24_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U6 ( .a ({new_AGEMA_signal_1189, SB_24_n11}), .b ({new_AGEMA_signal_756, SB_24_T1}), .c ({SubC_out_s1[88], SubC_out_s0[88]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U5 ( .a ({new_AGEMA_signal_1035, SB_24_n15}), .b ({SubC_in_s1[56], SubC_in_s0[56]}), .c ({new_AGEMA_signal_1189, SB_24_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U4 ( .a ({new_AGEMA_signal_754, SB_24_n10}), .b ({new_AGEMA_signal_755, SB_24_T0}), .c ({new_AGEMA_signal_1035, SB_24_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U1 ( .a ({SubC_in_s1[120], SubC_in_s0[120]}), .b ({new_AGEMA_signal_758, SB_24_T3}), .c ({new_AGEMA_signal_1036, SB_24_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_24_t0_AND_U1 ( .a ({SubC_in_s1[120], SubC_in_s0[120]}), .b ({SubC_in_s1[88], SubC_in_s0[88]}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_755, SB_24_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_24_t1_AND_U1 ( .a ({SubC_in_s1[120], SubC_in_s0[120]}), .b ({SubC_in_s1[56], SubC_in_s0[56]}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_756, SB_24_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_24_t2_AND_U1 ( .a ({SubC_in_s1[120], SubC_in_s0[120]}), .b ({SubC_in_s1[24], SubC_in_s0[24]}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_757, SB_24_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_24_t3_AND_U1 ( .a ({SubC_in_s1[88], SubC_in_s0[88]}), .b ({SubC_in_s1[24], SubC_in_s0[24]}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_758, SB_24_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U11 ( .a ({new_AGEMA_signal_1040, SB_23_n15}), .b ({new_AGEMA_signal_761, SB_23_n14}), .c ({SubC_out_s1[119], SubC_out_s0[119]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U9 ( .a ({new_AGEMA_signal_761, SB_23_n14}), .b ({new_AGEMA_signal_767, SB_23_T2}), .c ({new_AGEMA_signal_1039, SB_23_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U6 ( .a ({new_AGEMA_signal_1193, SB_23_n11}), .b ({new_AGEMA_signal_766, SB_23_T1}), .c ({SubC_out_s1[87], SubC_out_s0[87]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U5 ( .a ({new_AGEMA_signal_1040, SB_23_n15}), .b ({SubC_in_s1[55], SubC_in_s0[55]}), .c ({new_AGEMA_signal_1193, SB_23_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U4 ( .a ({new_AGEMA_signal_764, SB_23_n10}), .b ({new_AGEMA_signal_765, SB_23_T0}), .c ({new_AGEMA_signal_1040, SB_23_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U1 ( .a ({SubC_in_s1[119], SubC_in_s0[119]}), .b ({new_AGEMA_signal_768, SB_23_T3}), .c ({new_AGEMA_signal_1041, SB_23_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_23_t0_AND_U1 ( .a ({SubC_in_s1[119], SubC_in_s0[119]}), .b ({SubC_in_s1[87], SubC_in_s0[87]}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_765, SB_23_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_23_t1_AND_U1 ( .a ({SubC_in_s1[119], SubC_in_s0[119]}), .b ({SubC_in_s1[55], SubC_in_s0[55]}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_766, SB_23_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_23_t2_AND_U1 ( .a ({SubC_in_s1[119], SubC_in_s0[119]}), .b ({SubC_in_s1[23], SubC_in_s0[23]}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_767, SB_23_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_23_t3_AND_U1 ( .a ({SubC_in_s1[87], SubC_in_s0[87]}), .b ({SubC_in_s1[23], SubC_in_s0[23]}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_768, SB_23_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U11 ( .a ({new_AGEMA_signal_1045, SB_22_n15}), .b ({new_AGEMA_signal_771, SB_22_n14}), .c ({SubC_out_s1[118], SubC_out_s0[118]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U9 ( .a ({new_AGEMA_signal_771, SB_22_n14}), .b ({new_AGEMA_signal_777, SB_22_T2}), .c ({new_AGEMA_signal_1044, SB_22_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U6 ( .a ({new_AGEMA_signal_1197, SB_22_n11}), .b ({new_AGEMA_signal_776, SB_22_T1}), .c ({SubC_out_s1[86], SubC_out_s0[86]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U5 ( .a ({new_AGEMA_signal_1045, SB_22_n15}), .b ({SubC_in_s1[54], SubC_in_s0[54]}), .c ({new_AGEMA_signal_1197, SB_22_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U4 ( .a ({new_AGEMA_signal_774, SB_22_n10}), .b ({new_AGEMA_signal_775, SB_22_T0}), .c ({new_AGEMA_signal_1045, SB_22_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U1 ( .a ({SubC_in_s1[118], SubC_in_s0[118]}), .b ({new_AGEMA_signal_778, SB_22_T3}), .c ({new_AGEMA_signal_1046, SB_22_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_22_t0_AND_U1 ( .a ({SubC_in_s1[118], SubC_in_s0[118]}), .b ({SubC_in_s1[86], SubC_in_s0[86]}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_775, SB_22_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_22_t1_AND_U1 ( .a ({SubC_in_s1[118], SubC_in_s0[118]}), .b ({SubC_in_s1[54], SubC_in_s0[54]}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_776, SB_22_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_22_t2_AND_U1 ( .a ({SubC_in_s1[118], SubC_in_s0[118]}), .b ({SubC_in_s1[22], SubC_in_s0[22]}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_777, SB_22_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_22_t3_AND_U1 ( .a ({SubC_in_s1[86], SubC_in_s0[86]}), .b ({SubC_in_s1[22], SubC_in_s0[22]}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_778, SB_22_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U11 ( .a ({new_AGEMA_signal_1050, SB_21_n15}), .b ({new_AGEMA_signal_781, SB_21_n14}), .c ({SubC_out_s1[117], SubC_out_s0[117]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U9 ( .a ({new_AGEMA_signal_781, SB_21_n14}), .b ({new_AGEMA_signal_787, SB_21_T2}), .c ({new_AGEMA_signal_1049, SB_21_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U6 ( .a ({new_AGEMA_signal_1201, SB_21_n11}), .b ({new_AGEMA_signal_786, SB_21_T1}), .c ({SubC_out_s1[85], SubC_out_s0[85]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U5 ( .a ({new_AGEMA_signal_1050, SB_21_n15}), .b ({SubC_in_s1[53], SubC_in_s0[53]}), .c ({new_AGEMA_signal_1201, SB_21_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U4 ( .a ({new_AGEMA_signal_784, SB_21_n10}), .b ({new_AGEMA_signal_785, SB_21_T0}), .c ({new_AGEMA_signal_1050, SB_21_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U1 ( .a ({SubC_in_s1[117], SubC_in_s0[117]}), .b ({new_AGEMA_signal_788, SB_21_T3}), .c ({new_AGEMA_signal_1051, SB_21_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_21_t0_AND_U1 ( .a ({SubC_in_s1[117], SubC_in_s0[117]}), .b ({SubC_in_s1[85], SubC_in_s0[85]}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_785, SB_21_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_21_t1_AND_U1 ( .a ({SubC_in_s1[117], SubC_in_s0[117]}), .b ({SubC_in_s1[53], SubC_in_s0[53]}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_786, SB_21_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_21_t2_AND_U1 ( .a ({SubC_in_s1[117], SubC_in_s0[117]}), .b ({SubC_in_s1[21], SubC_in_s0[21]}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_787, SB_21_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_21_t3_AND_U1 ( .a ({SubC_in_s1[85], SubC_in_s0[85]}), .b ({SubC_in_s1[21], SubC_in_s0[21]}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_788, SB_21_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U11 ( .a ({new_AGEMA_signal_1055, SB_20_n15}), .b ({new_AGEMA_signal_791, SB_20_n14}), .c ({SubC_out_s1[116], SubC_out_s0[116]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U9 ( .a ({new_AGEMA_signal_791, SB_20_n14}), .b ({new_AGEMA_signal_797, SB_20_T2}), .c ({new_AGEMA_signal_1054, SB_20_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U6 ( .a ({new_AGEMA_signal_1205, SB_20_n11}), .b ({new_AGEMA_signal_796, SB_20_T1}), .c ({SubC_out_s1[84], SubC_out_s0[84]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U5 ( .a ({new_AGEMA_signal_1055, SB_20_n15}), .b ({SubC_in_s1[52], SubC_in_s0[52]}), .c ({new_AGEMA_signal_1205, SB_20_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U4 ( .a ({new_AGEMA_signal_794, SB_20_n10}), .b ({new_AGEMA_signal_795, SB_20_T0}), .c ({new_AGEMA_signal_1055, SB_20_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U1 ( .a ({SubC_in_s1[116], SubC_in_s0[116]}), .b ({new_AGEMA_signal_798, SB_20_T3}), .c ({new_AGEMA_signal_1056, SB_20_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_20_t0_AND_U1 ( .a ({SubC_in_s1[116], SubC_in_s0[116]}), .b ({SubC_in_s1[84], SubC_in_s0[84]}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_795, SB_20_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_20_t1_AND_U1 ( .a ({SubC_in_s1[116], SubC_in_s0[116]}), .b ({SubC_in_s1[52], SubC_in_s0[52]}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_796, SB_20_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_20_t2_AND_U1 ( .a ({SubC_in_s1[116], SubC_in_s0[116]}), .b ({SubC_in_s1[20], SubC_in_s0[20]}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_797, SB_20_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_20_t3_AND_U1 ( .a ({SubC_in_s1[84], SubC_in_s0[84]}), .b ({SubC_in_s1[20], SubC_in_s0[20]}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_798, SB_20_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U11 ( .a ({new_AGEMA_signal_1060, SB_19_n15}), .b ({new_AGEMA_signal_801, SB_19_n14}), .c ({SubC_out_s1[115], SubC_out_s0[115]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U9 ( .a ({new_AGEMA_signal_801, SB_19_n14}), .b ({new_AGEMA_signal_807, SB_19_T2}), .c ({new_AGEMA_signal_1059, SB_19_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U6 ( .a ({new_AGEMA_signal_1209, SB_19_n11}), .b ({new_AGEMA_signal_806, SB_19_T1}), .c ({SubC_out_s1[83], SubC_out_s0[83]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U5 ( .a ({new_AGEMA_signal_1060, SB_19_n15}), .b ({SubC_in_s1[51], SubC_in_s0[51]}), .c ({new_AGEMA_signal_1209, SB_19_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U4 ( .a ({new_AGEMA_signal_804, SB_19_n10}), .b ({new_AGEMA_signal_805, SB_19_T0}), .c ({new_AGEMA_signal_1060, SB_19_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U1 ( .a ({SubC_in_s1[115], SubC_in_s0[115]}), .b ({new_AGEMA_signal_808, SB_19_T3}), .c ({new_AGEMA_signal_1061, SB_19_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_19_t0_AND_U1 ( .a ({SubC_in_s1[115], SubC_in_s0[115]}), .b ({SubC_in_s1[83], SubC_in_s0[83]}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_805, SB_19_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_19_t1_AND_U1 ( .a ({SubC_in_s1[115], SubC_in_s0[115]}), .b ({SubC_in_s1[51], SubC_in_s0[51]}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_806, SB_19_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_19_t2_AND_U1 ( .a ({SubC_in_s1[115], SubC_in_s0[115]}), .b ({SubC_in_s1[19], SubC_in_s0[19]}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_807, SB_19_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_19_t3_AND_U1 ( .a ({SubC_in_s1[83], SubC_in_s0[83]}), .b ({SubC_in_s1[19], SubC_in_s0[19]}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_808, SB_19_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U11 ( .a ({new_AGEMA_signal_1065, SB_18_n15}), .b ({new_AGEMA_signal_811, SB_18_n14}), .c ({SubC_out_s1[114], SubC_out_s0[114]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U9 ( .a ({new_AGEMA_signal_811, SB_18_n14}), .b ({new_AGEMA_signal_817, SB_18_T2}), .c ({new_AGEMA_signal_1064, SB_18_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U6 ( .a ({new_AGEMA_signal_1213, SB_18_n11}), .b ({new_AGEMA_signal_816, SB_18_T1}), .c ({SubC_out_s1[82], SubC_out_s0[82]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U5 ( .a ({new_AGEMA_signal_1065, SB_18_n15}), .b ({SubC_in_s1[50], SubC_in_s0[50]}), .c ({new_AGEMA_signal_1213, SB_18_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U4 ( .a ({new_AGEMA_signal_814, SB_18_n10}), .b ({new_AGEMA_signal_815, SB_18_T0}), .c ({new_AGEMA_signal_1065, SB_18_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U1 ( .a ({SubC_in_s1[114], SubC_in_s0[114]}), .b ({new_AGEMA_signal_818, SB_18_T3}), .c ({new_AGEMA_signal_1066, SB_18_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_18_t0_AND_U1 ( .a ({SubC_in_s1[114], SubC_in_s0[114]}), .b ({SubC_in_s1[82], SubC_in_s0[82]}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_815, SB_18_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_18_t1_AND_U1 ( .a ({SubC_in_s1[114], SubC_in_s0[114]}), .b ({SubC_in_s1[50], SubC_in_s0[50]}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_816, SB_18_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_18_t2_AND_U1 ( .a ({SubC_in_s1[114], SubC_in_s0[114]}), .b ({SubC_in_s1[18], SubC_in_s0[18]}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_817, SB_18_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_18_t3_AND_U1 ( .a ({SubC_in_s1[82], SubC_in_s0[82]}), .b ({SubC_in_s1[18], SubC_in_s0[18]}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_818, SB_18_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U11 ( .a ({new_AGEMA_signal_1070, SB_17_n15}), .b ({new_AGEMA_signal_821, SB_17_n14}), .c ({SubC_out_s1[113], SubC_out_s0[113]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U9 ( .a ({new_AGEMA_signal_821, SB_17_n14}), .b ({new_AGEMA_signal_827, SB_17_T2}), .c ({new_AGEMA_signal_1069, SB_17_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U6 ( .a ({new_AGEMA_signal_1217, SB_17_n11}), .b ({new_AGEMA_signal_826, SB_17_T1}), .c ({SubC_out_s1[81], SubC_out_s0[81]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U5 ( .a ({new_AGEMA_signal_1070, SB_17_n15}), .b ({SubC_in_s1[49], SubC_in_s0[49]}), .c ({new_AGEMA_signal_1217, SB_17_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U4 ( .a ({new_AGEMA_signal_824, SB_17_n10}), .b ({new_AGEMA_signal_825, SB_17_T0}), .c ({new_AGEMA_signal_1070, SB_17_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U1 ( .a ({SubC_in_s1[113], SubC_in_s0[113]}), .b ({new_AGEMA_signal_828, SB_17_T3}), .c ({new_AGEMA_signal_1071, SB_17_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_17_t0_AND_U1 ( .a ({SubC_in_s1[113], SubC_in_s0[113]}), .b ({SubC_in_s1[81], SubC_in_s0[81]}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_825, SB_17_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_17_t1_AND_U1 ( .a ({SubC_in_s1[113], SubC_in_s0[113]}), .b ({SubC_in_s1[49], SubC_in_s0[49]}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_826, SB_17_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_17_t2_AND_U1 ( .a ({SubC_in_s1[113], SubC_in_s0[113]}), .b ({SubC_in_s1[17], SubC_in_s0[17]}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_827, SB_17_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_17_t3_AND_U1 ( .a ({SubC_in_s1[81], SubC_in_s0[81]}), .b ({SubC_in_s1[17], SubC_in_s0[17]}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_828, SB_17_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U11 ( .a ({new_AGEMA_signal_1075, SB_16_n15}), .b ({new_AGEMA_signal_831, SB_16_n14}), .c ({SubC_out_s1[112], SubC_out_s0[112]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U9 ( .a ({new_AGEMA_signal_831, SB_16_n14}), .b ({new_AGEMA_signal_837, SB_16_T2}), .c ({new_AGEMA_signal_1074, SB_16_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U6 ( .a ({new_AGEMA_signal_1221, SB_16_n11}), .b ({new_AGEMA_signal_836, SB_16_T1}), .c ({SubC_out_s1[80], SubC_out_s0[80]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U5 ( .a ({new_AGEMA_signal_1075, SB_16_n15}), .b ({SubC_in_s1[48], SubC_in_s0[48]}), .c ({new_AGEMA_signal_1221, SB_16_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U4 ( .a ({new_AGEMA_signal_834, SB_16_n10}), .b ({new_AGEMA_signal_835, SB_16_T0}), .c ({new_AGEMA_signal_1075, SB_16_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U1 ( .a ({SubC_in_s1[112], SubC_in_s0[112]}), .b ({new_AGEMA_signal_838, SB_16_T3}), .c ({new_AGEMA_signal_1076, SB_16_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_16_t0_AND_U1 ( .a ({SubC_in_s1[112], SubC_in_s0[112]}), .b ({SubC_in_s1[80], SubC_in_s0[80]}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_835, SB_16_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_16_t1_AND_U1 ( .a ({SubC_in_s1[112], SubC_in_s0[112]}), .b ({SubC_in_s1[48], SubC_in_s0[48]}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_836, SB_16_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_16_t2_AND_U1 ( .a ({SubC_in_s1[112], SubC_in_s0[112]}), .b ({SubC_in_s1[16], SubC_in_s0[16]}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_837, SB_16_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_16_t3_AND_U1 ( .a ({SubC_in_s1[80], SubC_in_s0[80]}), .b ({SubC_in_s1[16], SubC_in_s0[16]}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_838, SB_16_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U11 ( .a ({new_AGEMA_signal_1080, SB_15_n15}), .b ({new_AGEMA_signal_841, SB_15_n14}), .c ({SubC_out_s1[111], SubC_out_s0[111]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U9 ( .a ({new_AGEMA_signal_841, SB_15_n14}), .b ({new_AGEMA_signal_847, SB_15_T2}), .c ({new_AGEMA_signal_1079, SB_15_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U6 ( .a ({new_AGEMA_signal_1225, SB_15_n11}), .b ({new_AGEMA_signal_846, SB_15_T1}), .c ({SubC_out_s1[79], SubC_out_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U5 ( .a ({new_AGEMA_signal_1080, SB_15_n15}), .b ({SubC_in_s1[47], SubC_in_s0[47]}), .c ({new_AGEMA_signal_1225, SB_15_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U4 ( .a ({new_AGEMA_signal_844, SB_15_n10}), .b ({new_AGEMA_signal_845, SB_15_T0}), .c ({new_AGEMA_signal_1080, SB_15_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U1 ( .a ({SubC_in_s1[111], SubC_in_s0[111]}), .b ({new_AGEMA_signal_848, SB_15_T3}), .c ({new_AGEMA_signal_1081, SB_15_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_15_t0_AND_U1 ( .a ({SubC_in_s1[111], SubC_in_s0[111]}), .b ({SubC_in_s1[79], SubC_in_s0[79]}), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_845, SB_15_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_15_t1_AND_U1 ( .a ({SubC_in_s1[111], SubC_in_s0[111]}), .b ({SubC_in_s1[47], SubC_in_s0[47]}), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_846, SB_15_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_15_t2_AND_U1 ( .a ({SubC_in_s1[111], SubC_in_s0[111]}), .b ({SubC_in_s1[15], SubC_in_s0[15]}), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_847, SB_15_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_15_t3_AND_U1 ( .a ({SubC_in_s1[79], SubC_in_s0[79]}), .b ({SubC_in_s1[15], SubC_in_s0[15]}), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_848, SB_15_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U11 ( .a ({new_AGEMA_signal_1085, SB_14_n15}), .b ({new_AGEMA_signal_851, SB_14_n14}), .c ({SubC_out_s1[110], SubC_out_s0[110]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U9 ( .a ({new_AGEMA_signal_851, SB_14_n14}), .b ({new_AGEMA_signal_857, SB_14_T2}), .c ({new_AGEMA_signal_1084, SB_14_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U6 ( .a ({new_AGEMA_signal_1229, SB_14_n11}), .b ({new_AGEMA_signal_856, SB_14_T1}), .c ({SubC_out_s1[78], SubC_out_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U5 ( .a ({new_AGEMA_signal_1085, SB_14_n15}), .b ({SubC_in_s1[46], SubC_in_s0[46]}), .c ({new_AGEMA_signal_1229, SB_14_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U4 ( .a ({new_AGEMA_signal_854, SB_14_n10}), .b ({new_AGEMA_signal_855, SB_14_T0}), .c ({new_AGEMA_signal_1085, SB_14_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U1 ( .a ({SubC_in_s1[110], SubC_in_s0[110]}), .b ({new_AGEMA_signal_858, SB_14_T3}), .c ({new_AGEMA_signal_1086, SB_14_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_14_t0_AND_U1 ( .a ({SubC_in_s1[110], SubC_in_s0[110]}), .b ({SubC_in_s1[78], SubC_in_s0[78]}), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_855, SB_14_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_14_t1_AND_U1 ( .a ({SubC_in_s1[110], SubC_in_s0[110]}), .b ({SubC_in_s1[46], SubC_in_s0[46]}), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_856, SB_14_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_14_t2_AND_U1 ( .a ({SubC_in_s1[110], SubC_in_s0[110]}), .b ({SubC_in_s1[14], SubC_in_s0[14]}), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_857, SB_14_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_14_t3_AND_U1 ( .a ({SubC_in_s1[78], SubC_in_s0[78]}), .b ({SubC_in_s1[14], SubC_in_s0[14]}), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_858, SB_14_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U11 ( .a ({new_AGEMA_signal_1090, SB_13_n15}), .b ({new_AGEMA_signal_861, SB_13_n14}), .c ({SubC_out_s1[109], SubC_out_s0[109]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U9 ( .a ({new_AGEMA_signal_861, SB_13_n14}), .b ({new_AGEMA_signal_867, SB_13_T2}), .c ({new_AGEMA_signal_1089, SB_13_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U6 ( .a ({new_AGEMA_signal_1233, SB_13_n11}), .b ({new_AGEMA_signal_866, SB_13_T1}), .c ({SubC_out_s1[77], SubC_out_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U5 ( .a ({new_AGEMA_signal_1090, SB_13_n15}), .b ({SubC_in_s1[45], SubC_in_s0[45]}), .c ({new_AGEMA_signal_1233, SB_13_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U4 ( .a ({new_AGEMA_signal_864, SB_13_n10}), .b ({new_AGEMA_signal_865, SB_13_T0}), .c ({new_AGEMA_signal_1090, SB_13_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U1 ( .a ({SubC_in_s1[109], SubC_in_s0[109]}), .b ({new_AGEMA_signal_868, SB_13_T3}), .c ({new_AGEMA_signal_1091, SB_13_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_13_t0_AND_U1 ( .a ({SubC_in_s1[109], SubC_in_s0[109]}), .b ({SubC_in_s1[77], SubC_in_s0[77]}), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_865, SB_13_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_13_t1_AND_U1 ( .a ({SubC_in_s1[109], SubC_in_s0[109]}), .b ({SubC_in_s1[45], SubC_in_s0[45]}), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_866, SB_13_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_13_t2_AND_U1 ( .a ({SubC_in_s1[109], SubC_in_s0[109]}), .b ({SubC_in_s1[13], SubC_in_s0[13]}), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_867, SB_13_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_13_t3_AND_U1 ( .a ({SubC_in_s1[77], SubC_in_s0[77]}), .b ({SubC_in_s1[13], SubC_in_s0[13]}), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_868, SB_13_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U11 ( .a ({new_AGEMA_signal_1095, SB_12_n15}), .b ({new_AGEMA_signal_871, SB_12_n14}), .c ({SubC_out_s1[108], SubC_out_s0[108]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U9 ( .a ({new_AGEMA_signal_871, SB_12_n14}), .b ({new_AGEMA_signal_877, SB_12_T2}), .c ({new_AGEMA_signal_1094, SB_12_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U6 ( .a ({new_AGEMA_signal_1237, SB_12_n11}), .b ({new_AGEMA_signal_876, SB_12_T1}), .c ({SubC_out_s1[76], SubC_out_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U5 ( .a ({new_AGEMA_signal_1095, SB_12_n15}), .b ({SubC_in_s1[44], SubC_in_s0[44]}), .c ({new_AGEMA_signal_1237, SB_12_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U4 ( .a ({new_AGEMA_signal_874, SB_12_n10}), .b ({new_AGEMA_signal_875, SB_12_T0}), .c ({new_AGEMA_signal_1095, SB_12_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U1 ( .a ({SubC_in_s1[108], SubC_in_s0[108]}), .b ({new_AGEMA_signal_878, SB_12_T3}), .c ({new_AGEMA_signal_1096, SB_12_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_12_t0_AND_U1 ( .a ({SubC_in_s1[108], SubC_in_s0[108]}), .b ({SubC_in_s1[76], SubC_in_s0[76]}), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_875, SB_12_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_12_t1_AND_U1 ( .a ({SubC_in_s1[108], SubC_in_s0[108]}), .b ({SubC_in_s1[44], SubC_in_s0[44]}), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_876, SB_12_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_12_t2_AND_U1 ( .a ({SubC_in_s1[108], SubC_in_s0[108]}), .b ({SubC_in_s1[12], SubC_in_s0[12]}), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_877, SB_12_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_12_t3_AND_U1 ( .a ({SubC_in_s1[76], SubC_in_s0[76]}), .b ({SubC_in_s1[12], SubC_in_s0[12]}), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_878, SB_12_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U11 ( .a ({new_AGEMA_signal_1100, SB_11_n15}), .b ({new_AGEMA_signal_881, SB_11_n14}), .c ({SubC_out_s1[107], SubC_out_s0[107]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U9 ( .a ({new_AGEMA_signal_881, SB_11_n14}), .b ({new_AGEMA_signal_887, SB_11_T2}), .c ({new_AGEMA_signal_1099, SB_11_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U6 ( .a ({new_AGEMA_signal_1241, SB_11_n11}), .b ({new_AGEMA_signal_886, SB_11_T1}), .c ({SubC_out_s1[75], SubC_out_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U5 ( .a ({new_AGEMA_signal_1100, SB_11_n15}), .b ({SubC_in_s1[43], SubC_in_s0[43]}), .c ({new_AGEMA_signal_1241, SB_11_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U4 ( .a ({new_AGEMA_signal_884, SB_11_n10}), .b ({new_AGEMA_signal_885, SB_11_T0}), .c ({new_AGEMA_signal_1100, SB_11_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U1 ( .a ({SubC_in_s1[107], SubC_in_s0[107]}), .b ({new_AGEMA_signal_888, SB_11_T3}), .c ({new_AGEMA_signal_1101, SB_11_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_11_t0_AND_U1 ( .a ({SubC_in_s1[107], SubC_in_s0[107]}), .b ({SubC_in_s1[75], SubC_in_s0[75]}), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_885, SB_11_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_11_t1_AND_U1 ( .a ({SubC_in_s1[107], SubC_in_s0[107]}), .b ({SubC_in_s1[43], SubC_in_s0[43]}), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_886, SB_11_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_11_t2_AND_U1 ( .a ({SubC_in_s1[107], SubC_in_s0[107]}), .b ({SubC_in_s1[11], SubC_in_s0[11]}), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_887, SB_11_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_11_t3_AND_U1 ( .a ({SubC_in_s1[75], SubC_in_s0[75]}), .b ({SubC_in_s1[11], SubC_in_s0[11]}), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_888, SB_11_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U11 ( .a ({new_AGEMA_signal_1105, SB_10_n15}), .b ({new_AGEMA_signal_891, SB_10_n14}), .c ({SubC_out_s1[106], SubC_out_s0[106]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U9 ( .a ({new_AGEMA_signal_891, SB_10_n14}), .b ({new_AGEMA_signal_897, SB_10_T2}), .c ({new_AGEMA_signal_1104, SB_10_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U6 ( .a ({new_AGEMA_signal_1245, SB_10_n11}), .b ({new_AGEMA_signal_896, SB_10_T1}), .c ({SubC_out_s1[74], SubC_out_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U5 ( .a ({new_AGEMA_signal_1105, SB_10_n15}), .b ({SubC_in_s1[42], SubC_in_s0[42]}), .c ({new_AGEMA_signal_1245, SB_10_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U4 ( .a ({new_AGEMA_signal_894, SB_10_n10}), .b ({new_AGEMA_signal_895, SB_10_T0}), .c ({new_AGEMA_signal_1105, SB_10_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U1 ( .a ({SubC_in_s1[106], SubC_in_s0[106]}), .b ({new_AGEMA_signal_898, SB_10_T3}), .c ({new_AGEMA_signal_1106, SB_10_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_10_t0_AND_U1 ( .a ({SubC_in_s1[106], SubC_in_s0[106]}), .b ({SubC_in_s1[74], SubC_in_s0[74]}), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_895, SB_10_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_10_t1_AND_U1 ( .a ({SubC_in_s1[106], SubC_in_s0[106]}), .b ({SubC_in_s1[42], SubC_in_s0[42]}), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_896, SB_10_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_10_t2_AND_U1 ( .a ({SubC_in_s1[106], SubC_in_s0[106]}), .b ({SubC_in_s1[10], SubC_in_s0[10]}), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_897, SB_10_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_10_t3_AND_U1 ( .a ({SubC_in_s1[74], SubC_in_s0[74]}), .b ({SubC_in_s1[10], SubC_in_s0[10]}), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_898, SB_10_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U11 ( .a ({new_AGEMA_signal_1110, SB_9_n15}), .b ({new_AGEMA_signal_901, SB_9_n14}), .c ({SubC_out_s1[105], SubC_out_s0[105]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U9 ( .a ({new_AGEMA_signal_901, SB_9_n14}), .b ({new_AGEMA_signal_907, SB_9_T2}), .c ({new_AGEMA_signal_1109, SB_9_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U6 ( .a ({new_AGEMA_signal_1249, SB_9_n11}), .b ({new_AGEMA_signal_906, SB_9_T1}), .c ({SubC_out_s1[73], SubC_out_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U5 ( .a ({new_AGEMA_signal_1110, SB_9_n15}), .b ({SubC_in_s1[41], SubC_in_s0[41]}), .c ({new_AGEMA_signal_1249, SB_9_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U4 ( .a ({new_AGEMA_signal_904, SB_9_n10}), .b ({new_AGEMA_signal_905, SB_9_T0}), .c ({new_AGEMA_signal_1110, SB_9_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U1 ( .a ({SubC_in_s1[105], SubC_in_s0[105]}), .b ({new_AGEMA_signal_908, SB_9_T3}), .c ({new_AGEMA_signal_1111, SB_9_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_9_t0_AND_U1 ( .a ({SubC_in_s1[105], SubC_in_s0[105]}), .b ({SubC_in_s1[73], SubC_in_s0[73]}), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_905, SB_9_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_9_t1_AND_U1 ( .a ({SubC_in_s1[105], SubC_in_s0[105]}), .b ({SubC_in_s1[41], SubC_in_s0[41]}), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_906, SB_9_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_9_t2_AND_U1 ( .a ({SubC_in_s1[105], SubC_in_s0[105]}), .b ({SubC_in_s1[9], SubC_in_s0[9]}), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_907, SB_9_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_9_t3_AND_U1 ( .a ({SubC_in_s1[73], SubC_in_s0[73]}), .b ({SubC_in_s1[9], SubC_in_s0[9]}), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_908, SB_9_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U11 ( .a ({new_AGEMA_signal_1115, SB_8_n15}), .b ({new_AGEMA_signal_911, SB_8_n14}), .c ({SubC_out_s1[104], SubC_out_s0[104]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U9 ( .a ({new_AGEMA_signal_911, SB_8_n14}), .b ({new_AGEMA_signal_917, SB_8_T2}), .c ({new_AGEMA_signal_1114, SB_8_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U6 ( .a ({new_AGEMA_signal_1253, SB_8_n11}), .b ({new_AGEMA_signal_916, SB_8_T1}), .c ({SubC_out_s1[72], SubC_out_s0[72]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U5 ( .a ({new_AGEMA_signal_1115, SB_8_n15}), .b ({SubC_in_s1[40], SubC_in_s0[40]}), .c ({new_AGEMA_signal_1253, SB_8_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U4 ( .a ({new_AGEMA_signal_914, SB_8_n10}), .b ({new_AGEMA_signal_915, SB_8_T0}), .c ({new_AGEMA_signal_1115, SB_8_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U1 ( .a ({SubC_in_s1[104], SubC_in_s0[104]}), .b ({new_AGEMA_signal_918, SB_8_T3}), .c ({new_AGEMA_signal_1116, SB_8_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_8_t0_AND_U1 ( .a ({SubC_in_s1[104], SubC_in_s0[104]}), .b ({SubC_in_s1[72], SubC_in_s0[72]}), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_915, SB_8_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_8_t1_AND_U1 ( .a ({SubC_in_s1[104], SubC_in_s0[104]}), .b ({SubC_in_s1[40], SubC_in_s0[40]}), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_916, SB_8_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_8_t2_AND_U1 ( .a ({SubC_in_s1[104], SubC_in_s0[104]}), .b ({SubC_in_s1[8], SubC_in_s0[8]}), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_917, SB_8_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_8_t3_AND_U1 ( .a ({SubC_in_s1[72], SubC_in_s0[72]}), .b ({SubC_in_s1[8], SubC_in_s0[8]}), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_918, SB_8_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U11 ( .a ({new_AGEMA_signal_1120, SB_7_n15}), .b ({new_AGEMA_signal_921, SB_7_n14}), .c ({SubC_out_s1[103], SubC_out_s0[103]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U9 ( .a ({new_AGEMA_signal_921, SB_7_n14}), .b ({new_AGEMA_signal_927, SB_7_T2}), .c ({new_AGEMA_signal_1119, SB_7_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U6 ( .a ({new_AGEMA_signal_1257, SB_7_n11}), .b ({new_AGEMA_signal_926, SB_7_T1}), .c ({SubC_out_s1[71], SubC_out_s0[71]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U5 ( .a ({new_AGEMA_signal_1120, SB_7_n15}), .b ({SubC_in_s1[39], SubC_in_s0[39]}), .c ({new_AGEMA_signal_1257, SB_7_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U4 ( .a ({new_AGEMA_signal_924, SB_7_n10}), .b ({new_AGEMA_signal_925, SB_7_T0}), .c ({new_AGEMA_signal_1120, SB_7_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U1 ( .a ({SubC_in_s1[103], SubC_in_s0[103]}), .b ({new_AGEMA_signal_928, SB_7_T3}), .c ({new_AGEMA_signal_1121, SB_7_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_7_t0_AND_U1 ( .a ({SubC_in_s1[103], SubC_in_s0[103]}), .b ({SubC_in_s1[71], SubC_in_s0[71]}), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_925, SB_7_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_7_t1_AND_U1 ( .a ({SubC_in_s1[103], SubC_in_s0[103]}), .b ({SubC_in_s1[39], SubC_in_s0[39]}), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_926, SB_7_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_7_t2_AND_U1 ( .a ({SubC_in_s1[103], SubC_in_s0[103]}), .b ({SubC_in_s1[7], SubC_in_s0[7]}), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_927, SB_7_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_7_t3_AND_U1 ( .a ({SubC_in_s1[71], SubC_in_s0[71]}), .b ({SubC_in_s1[7], SubC_in_s0[7]}), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_928, SB_7_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U11 ( .a ({new_AGEMA_signal_1125, SB_6_n15}), .b ({new_AGEMA_signal_931, SB_6_n14}), .c ({SubC_out_s1[102], SubC_out_s0[102]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U9 ( .a ({new_AGEMA_signal_931, SB_6_n14}), .b ({new_AGEMA_signal_937, SB_6_T2}), .c ({new_AGEMA_signal_1124, SB_6_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U6 ( .a ({new_AGEMA_signal_1261, SB_6_n11}), .b ({new_AGEMA_signal_936, SB_6_T1}), .c ({SubC_out_s1[70], SubC_out_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U5 ( .a ({new_AGEMA_signal_1125, SB_6_n15}), .b ({SubC_in_s1[38], SubC_in_s0[38]}), .c ({new_AGEMA_signal_1261, SB_6_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U4 ( .a ({new_AGEMA_signal_934, SB_6_n10}), .b ({new_AGEMA_signal_935, SB_6_T0}), .c ({new_AGEMA_signal_1125, SB_6_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U1 ( .a ({SubC_in_s1[102], SubC_in_s0[102]}), .b ({new_AGEMA_signal_938, SB_6_T3}), .c ({new_AGEMA_signal_1126, SB_6_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_6_t0_AND_U1 ( .a ({SubC_in_s1[102], SubC_in_s0[102]}), .b ({SubC_in_s1[70], SubC_in_s0[70]}), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_935, SB_6_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_6_t1_AND_U1 ( .a ({SubC_in_s1[102], SubC_in_s0[102]}), .b ({SubC_in_s1[38], SubC_in_s0[38]}), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_936, SB_6_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_6_t2_AND_U1 ( .a ({SubC_in_s1[102], SubC_in_s0[102]}), .b ({SubC_in_s1[6], SubC_in_s0[6]}), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_937, SB_6_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_6_t3_AND_U1 ( .a ({SubC_in_s1[70], SubC_in_s0[70]}), .b ({SubC_in_s1[6], SubC_in_s0[6]}), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_938, SB_6_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U11 ( .a ({new_AGEMA_signal_1130, SB_5_n15}), .b ({new_AGEMA_signal_941, SB_5_n14}), .c ({SubC_out_s1[101], SubC_out_s0[101]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U9 ( .a ({new_AGEMA_signal_941, SB_5_n14}), .b ({new_AGEMA_signal_947, SB_5_T2}), .c ({new_AGEMA_signal_1129, SB_5_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U6 ( .a ({new_AGEMA_signal_1265, SB_5_n11}), .b ({new_AGEMA_signal_946, SB_5_T1}), .c ({SubC_out_s1[69], SubC_out_s0[69]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U5 ( .a ({new_AGEMA_signal_1130, SB_5_n15}), .b ({SubC_in_s1[37], SubC_in_s0[37]}), .c ({new_AGEMA_signal_1265, SB_5_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U4 ( .a ({new_AGEMA_signal_944, SB_5_n10}), .b ({new_AGEMA_signal_945, SB_5_T0}), .c ({new_AGEMA_signal_1130, SB_5_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U1 ( .a ({SubC_in_s1[101], SubC_in_s0[101]}), .b ({new_AGEMA_signal_948, SB_5_T3}), .c ({new_AGEMA_signal_1131, SB_5_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_5_t0_AND_U1 ( .a ({SubC_in_s1[101], SubC_in_s0[101]}), .b ({SubC_in_s1[69], SubC_in_s0[69]}), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_945, SB_5_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_5_t1_AND_U1 ( .a ({SubC_in_s1[101], SubC_in_s0[101]}), .b ({SubC_in_s1[37], SubC_in_s0[37]}), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_946, SB_5_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_5_t2_AND_U1 ( .a ({SubC_in_s1[101], SubC_in_s0[101]}), .b ({SubC_in_s1[5], SubC_in_s0[5]}), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_947, SB_5_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_5_t3_AND_U1 ( .a ({SubC_in_s1[69], SubC_in_s0[69]}), .b ({SubC_in_s1[5], SubC_in_s0[5]}), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_948, SB_5_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U11 ( .a ({new_AGEMA_signal_1135, SB_4_n15}), .b ({new_AGEMA_signal_951, SB_4_n14}), .c ({SubC_out_s1[100], SubC_out_s0[100]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U9 ( .a ({new_AGEMA_signal_951, SB_4_n14}), .b ({new_AGEMA_signal_957, SB_4_T2}), .c ({new_AGEMA_signal_1134, SB_4_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U6 ( .a ({new_AGEMA_signal_1269, SB_4_n11}), .b ({new_AGEMA_signal_956, SB_4_T1}), .c ({SubC_out_s1[68], SubC_out_s0[68]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U5 ( .a ({new_AGEMA_signal_1135, SB_4_n15}), .b ({SubC_in_s1[36], SubC_in_s0[36]}), .c ({new_AGEMA_signal_1269, SB_4_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U4 ( .a ({new_AGEMA_signal_954, SB_4_n10}), .b ({new_AGEMA_signal_955, SB_4_T0}), .c ({new_AGEMA_signal_1135, SB_4_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U1 ( .a ({SubC_in_s1[100], SubC_in_s0[100]}), .b ({new_AGEMA_signal_958, SB_4_T3}), .c ({new_AGEMA_signal_1136, SB_4_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_4_t0_AND_U1 ( .a ({SubC_in_s1[100], SubC_in_s0[100]}), .b ({SubC_in_s1[68], SubC_in_s0[68]}), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_955, SB_4_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_4_t1_AND_U1 ( .a ({SubC_in_s1[100], SubC_in_s0[100]}), .b ({SubC_in_s1[36], SubC_in_s0[36]}), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_956, SB_4_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_4_t2_AND_U1 ( .a ({SubC_in_s1[100], SubC_in_s0[100]}), .b ({SubC_in_s1[4], SubC_in_s0[4]}), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_957, SB_4_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_4_t3_AND_U1 ( .a ({SubC_in_s1[68], SubC_in_s0[68]}), .b ({SubC_in_s1[4], SubC_in_s0[4]}), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_958, SB_4_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U11 ( .a ({new_AGEMA_signal_1140, SB_3_n15}), .b ({new_AGEMA_signal_961, SB_3_n14}), .c ({SubC_out_s1[99], SubC_out_s0[99]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U9 ( .a ({new_AGEMA_signal_961, SB_3_n14}), .b ({new_AGEMA_signal_967, SB_3_T2}), .c ({new_AGEMA_signal_1139, SB_3_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U6 ( .a ({new_AGEMA_signal_1273, SB_3_n11}), .b ({new_AGEMA_signal_966, SB_3_T1}), .c ({SubC_out_s1[67], SubC_out_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U5 ( .a ({new_AGEMA_signal_1140, SB_3_n15}), .b ({SubC_in_s1[35], SubC_in_s0[35]}), .c ({new_AGEMA_signal_1273, SB_3_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U4 ( .a ({new_AGEMA_signal_964, SB_3_n10}), .b ({new_AGEMA_signal_965, SB_3_T0}), .c ({new_AGEMA_signal_1140, SB_3_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U1 ( .a ({SubC_in_s1[99], SubC_in_s0[99]}), .b ({new_AGEMA_signal_968, SB_3_T3}), .c ({new_AGEMA_signal_1141, SB_3_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_3_t0_AND_U1 ( .a ({SubC_in_s1[99], SubC_in_s0[99]}), .b ({SubC_in_s1[67], SubC_in_s0[67]}), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_965, SB_3_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_3_t1_AND_U1 ( .a ({SubC_in_s1[99], SubC_in_s0[99]}), .b ({SubC_in_s1[35], SubC_in_s0[35]}), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_966, SB_3_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_3_t2_AND_U1 ( .a ({SubC_in_s1[99], SubC_in_s0[99]}), .b ({SubC_in_s1[3], SubC_in_s0[3]}), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_967, SB_3_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_3_t3_AND_U1 ( .a ({SubC_in_s1[67], SubC_in_s0[67]}), .b ({SubC_in_s1[3], SubC_in_s0[3]}), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_968, SB_3_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U11 ( .a ({new_AGEMA_signal_1145, SB_2_n15}), .b ({new_AGEMA_signal_971, SB_2_n14}), .c ({SubC_out_s1[98], SubC_out_s0[98]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U9 ( .a ({new_AGEMA_signal_971, SB_2_n14}), .b ({new_AGEMA_signal_977, SB_2_T2}), .c ({new_AGEMA_signal_1144, SB_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U6 ( .a ({new_AGEMA_signal_1277, SB_2_n11}), .b ({new_AGEMA_signal_976, SB_2_T1}), .c ({SubC_out_s1[66], SubC_out_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U5 ( .a ({new_AGEMA_signal_1145, SB_2_n15}), .b ({SubC_in_s1[34], SubC_in_s0[34]}), .c ({new_AGEMA_signal_1277, SB_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U4 ( .a ({new_AGEMA_signal_974, SB_2_n10}), .b ({new_AGEMA_signal_975, SB_2_T0}), .c ({new_AGEMA_signal_1145, SB_2_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U1 ( .a ({SubC_in_s1[98], SubC_in_s0[98]}), .b ({new_AGEMA_signal_978, SB_2_T3}), .c ({new_AGEMA_signal_1146, SB_2_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_2_t0_AND_U1 ( .a ({SubC_in_s1[98], SubC_in_s0[98]}), .b ({SubC_in_s1[66], SubC_in_s0[66]}), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_975, SB_2_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_2_t1_AND_U1 ( .a ({SubC_in_s1[98], SubC_in_s0[98]}), .b ({SubC_in_s1[34], SubC_in_s0[34]}), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_976, SB_2_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_2_t2_AND_U1 ( .a ({SubC_in_s1[98], SubC_in_s0[98]}), .b ({SubC_in_s1[2], SubC_in_s0[2]}), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_977, SB_2_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_2_t3_AND_U1 ( .a ({SubC_in_s1[66], SubC_in_s0[66]}), .b ({SubC_in_s1[2], SubC_in_s0[2]}), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_978, SB_2_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U11 ( .a ({new_AGEMA_signal_1150, SB_1_n15}), .b ({new_AGEMA_signal_981, SB_1_n14}), .c ({SubC_out_s1[97], SubC_out_s0[97]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U9 ( .a ({new_AGEMA_signal_981, SB_1_n14}), .b ({new_AGEMA_signal_987, SB_1_T2}), .c ({new_AGEMA_signal_1149, SB_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U6 ( .a ({new_AGEMA_signal_1281, SB_1_n11}), .b ({new_AGEMA_signal_986, SB_1_T1}), .c ({SubC_out_s1[65], SubC_out_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U5 ( .a ({new_AGEMA_signal_1150, SB_1_n15}), .b ({SubC_in_s1[33], SubC_in_s0[33]}), .c ({new_AGEMA_signal_1281, SB_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U4 ( .a ({new_AGEMA_signal_984, SB_1_n10}), .b ({new_AGEMA_signal_985, SB_1_T0}), .c ({new_AGEMA_signal_1150, SB_1_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U1 ( .a ({SubC_in_s1[97], SubC_in_s0[97]}), .b ({new_AGEMA_signal_988, SB_1_T3}), .c ({new_AGEMA_signal_1151, SB_1_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_1_t0_AND_U1 ( .a ({SubC_in_s1[97], SubC_in_s0[97]}), .b ({SubC_in_s1[65], SubC_in_s0[65]}), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_985, SB_1_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_1_t1_AND_U1 ( .a ({SubC_in_s1[97], SubC_in_s0[97]}), .b ({SubC_in_s1[33], SubC_in_s0[33]}), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_986, SB_1_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_1_t2_AND_U1 ( .a ({SubC_in_s1[97], SubC_in_s0[97]}), .b ({SubC_in_s1[1], SubC_in_s0[1]}), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_987, SB_1_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_1_t3_AND_U1 ( .a ({SubC_in_s1[65], SubC_in_s0[65]}), .b ({SubC_in_s1[1], SubC_in_s0[1]}), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_988, SB_1_T3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U11 ( .a ({new_AGEMA_signal_1155, SB_0_n15}), .b ({new_AGEMA_signal_991, SB_0_n14}), .c ({SubC_out_s1[96], SubC_out_s0[96]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U9 ( .a ({new_AGEMA_signal_991, SB_0_n14}), .b ({new_AGEMA_signal_997, SB_0_T2}), .c ({new_AGEMA_signal_1154, SB_0_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U6 ( .a ({new_AGEMA_signal_1285, SB_0_n11}), .b ({new_AGEMA_signal_996, SB_0_T1}), .c ({SubC_out_s1[64], SubC_out_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U5 ( .a ({new_AGEMA_signal_1155, SB_0_n15}), .b ({SubC_in_s1[32], SubC_in_s0[32]}), .c ({new_AGEMA_signal_1285, SB_0_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U4 ( .a ({new_AGEMA_signal_994, SB_0_n10}), .b ({new_AGEMA_signal_995, SB_0_T0}), .c ({new_AGEMA_signal_1155, SB_0_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U1 ( .a ({SubC_in_s1[96], SubC_in_s0[96]}), .b ({new_AGEMA_signal_998, SB_0_T3}), .c ({new_AGEMA_signal_1156, SB_0_n9}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_0_t0_AND_U1 ( .a ({SubC_in_s1[96], SubC_in_s0[96]}), .b ({SubC_in_s1[64], SubC_in_s0[64]}), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_995, SB_0_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_0_t1_AND_U1 ( .a ({SubC_in_s1[96], SubC_in_s0[96]}), .b ({SubC_in_s1[32], SubC_in_s0[32]}), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_996, SB_0_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_0_t2_AND_U1 ( .a ({SubC_in_s1[96], SubC_in_s0[96]}), .b ({SubC_in_s1[0], SubC_in_s0[0]}), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_997, SB_0_T2}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_0_t3_AND_U1 ( .a ({SubC_in_s1[64], SubC_in_s0[64]}), .b ({SubC_in_s1[0], SubC_in_s0[0]}), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_998, SB_0_T3}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U10 ( .a ({new_AGEMA_signal_1160, SB_31_n13}), .b ({new_AGEMA_signal_999, SB_31_n12}), .c ({SubC_out_s1[63], SubC_out_s0[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U7 ( .a ({new_AGEMA_signal_1002, SB_31_T4}), .b ({new_AGEMA_signal_688, SB_31_T3}), .c ({new_AGEMA_signal_1160, SB_31_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_31_U2 ( .a ({new_AGEMA_signal_1001, SB_31_n9}), .b ({new_AGEMA_signal_1003, SB_31_T5}), .c ({SubC_out_s1[31], SubC_out_s0[31]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_31_t4_AND_U1 ( .a ({SubC_in_s1[63], SubC_in_s0[63]}), .b ({new_AGEMA_signal_688, SB_31_T3}), .clk (clk), .r (Fresh[128]), .c ({new_AGEMA_signal_1002, SB_31_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_31_t5_AND_U1 ( .a ({SubC_in_s1[63], SubC_in_s0[63]}), .b ({new_AGEMA_signal_687, SB_31_T2}), .clk (clk), .r (Fresh[129]), .c ({new_AGEMA_signal_1003, SB_31_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U10 ( .a ({new_AGEMA_signal_1164, SB_30_n13}), .b ({new_AGEMA_signal_1004, SB_30_n12}), .c ({SubC_out_s1[62], SubC_out_s0[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U7 ( .a ({new_AGEMA_signal_1007, SB_30_T4}), .b ({new_AGEMA_signal_698, SB_30_T3}), .c ({new_AGEMA_signal_1164, SB_30_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_30_U2 ( .a ({new_AGEMA_signal_1006, SB_30_n9}), .b ({new_AGEMA_signal_1008, SB_30_T5}), .c ({SubC_out_s1[30], SubC_out_s0[30]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_30_t4_AND_U1 ( .a ({SubC_in_s1[62], SubC_in_s0[62]}), .b ({new_AGEMA_signal_698, SB_30_T3}), .clk (clk), .r (Fresh[130]), .c ({new_AGEMA_signal_1007, SB_30_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_30_t5_AND_U1 ( .a ({SubC_in_s1[62], SubC_in_s0[62]}), .b ({new_AGEMA_signal_697, SB_30_T2}), .clk (clk), .r (Fresh[131]), .c ({new_AGEMA_signal_1008, SB_30_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U10 ( .a ({new_AGEMA_signal_1168, SB_29_n13}), .b ({new_AGEMA_signal_1009, SB_29_n12}), .c ({SubC_out_s1[61], SubC_out_s0[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U7 ( .a ({new_AGEMA_signal_1012, SB_29_T4}), .b ({new_AGEMA_signal_708, SB_29_T3}), .c ({new_AGEMA_signal_1168, SB_29_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_29_U2 ( .a ({new_AGEMA_signal_1011, SB_29_n9}), .b ({new_AGEMA_signal_1013, SB_29_T5}), .c ({SubC_out_s1[29], SubC_out_s0[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_29_t4_AND_U1 ( .a ({SubC_in_s1[61], SubC_in_s0[61]}), .b ({new_AGEMA_signal_708, SB_29_T3}), .clk (clk), .r (Fresh[132]), .c ({new_AGEMA_signal_1012, SB_29_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_29_t5_AND_U1 ( .a ({SubC_in_s1[61], SubC_in_s0[61]}), .b ({new_AGEMA_signal_707, SB_29_T2}), .clk (clk), .r (Fresh[133]), .c ({new_AGEMA_signal_1013, SB_29_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U10 ( .a ({new_AGEMA_signal_1172, SB_28_n13}), .b ({new_AGEMA_signal_1014, SB_28_n12}), .c ({SubC_out_s1[60], SubC_out_s0[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U7 ( .a ({new_AGEMA_signal_1017, SB_28_T4}), .b ({new_AGEMA_signal_718, SB_28_T3}), .c ({new_AGEMA_signal_1172, SB_28_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_28_U2 ( .a ({new_AGEMA_signal_1016, SB_28_n9}), .b ({new_AGEMA_signal_1018, SB_28_T5}), .c ({SubC_out_s1[28], SubC_out_s0[28]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_28_t4_AND_U1 ( .a ({SubC_in_s1[60], SubC_in_s0[60]}), .b ({new_AGEMA_signal_718, SB_28_T3}), .clk (clk), .r (Fresh[134]), .c ({new_AGEMA_signal_1017, SB_28_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_28_t5_AND_U1 ( .a ({SubC_in_s1[60], SubC_in_s0[60]}), .b ({new_AGEMA_signal_717, SB_28_T2}), .clk (clk), .r (Fresh[135]), .c ({new_AGEMA_signal_1018, SB_28_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U10 ( .a ({new_AGEMA_signal_1176, SB_27_n13}), .b ({new_AGEMA_signal_1019, SB_27_n12}), .c ({SubC_out_s1[59], SubC_out_s0[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U7 ( .a ({new_AGEMA_signal_1022, SB_27_T4}), .b ({new_AGEMA_signal_728, SB_27_T3}), .c ({new_AGEMA_signal_1176, SB_27_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_27_U2 ( .a ({new_AGEMA_signal_1021, SB_27_n9}), .b ({new_AGEMA_signal_1023, SB_27_T5}), .c ({SubC_out_s1[27], SubC_out_s0[27]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_27_t4_AND_U1 ( .a ({SubC_in_s1[59], SubC_in_s0[59]}), .b ({new_AGEMA_signal_728, SB_27_T3}), .clk (clk), .r (Fresh[136]), .c ({new_AGEMA_signal_1022, SB_27_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_27_t5_AND_U1 ( .a ({SubC_in_s1[59], SubC_in_s0[59]}), .b ({new_AGEMA_signal_727, SB_27_T2}), .clk (clk), .r (Fresh[137]), .c ({new_AGEMA_signal_1023, SB_27_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U10 ( .a ({new_AGEMA_signal_1180, SB_26_n13}), .b ({new_AGEMA_signal_1024, SB_26_n12}), .c ({SubC_out_s1[58], SubC_out_s0[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U7 ( .a ({new_AGEMA_signal_1027, SB_26_T4}), .b ({new_AGEMA_signal_738, SB_26_T3}), .c ({new_AGEMA_signal_1180, SB_26_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_26_U2 ( .a ({new_AGEMA_signal_1026, SB_26_n9}), .b ({new_AGEMA_signal_1028, SB_26_T5}), .c ({SubC_out_s1[26], SubC_out_s0[26]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_26_t4_AND_U1 ( .a ({SubC_in_s1[58], SubC_in_s0[58]}), .b ({new_AGEMA_signal_738, SB_26_T3}), .clk (clk), .r (Fresh[138]), .c ({new_AGEMA_signal_1027, SB_26_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_26_t5_AND_U1 ( .a ({SubC_in_s1[58], SubC_in_s0[58]}), .b ({new_AGEMA_signal_737, SB_26_T2}), .clk (clk), .r (Fresh[139]), .c ({new_AGEMA_signal_1028, SB_26_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U10 ( .a ({new_AGEMA_signal_1184, SB_25_n13}), .b ({new_AGEMA_signal_1029, SB_25_n12}), .c ({SubC_out_s1[57], SubC_out_s0[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U7 ( .a ({new_AGEMA_signal_1032, SB_25_T4}), .b ({new_AGEMA_signal_748, SB_25_T3}), .c ({new_AGEMA_signal_1184, SB_25_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_25_U2 ( .a ({new_AGEMA_signal_1031, SB_25_n9}), .b ({new_AGEMA_signal_1033, SB_25_T5}), .c ({SubC_out_s1[25], SubC_out_s0[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_25_t4_AND_U1 ( .a ({SubC_in_s1[57], SubC_in_s0[57]}), .b ({new_AGEMA_signal_748, SB_25_T3}), .clk (clk), .r (Fresh[140]), .c ({new_AGEMA_signal_1032, SB_25_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_25_t5_AND_U1 ( .a ({SubC_in_s1[57], SubC_in_s0[57]}), .b ({new_AGEMA_signal_747, SB_25_T2}), .clk (clk), .r (Fresh[141]), .c ({new_AGEMA_signal_1033, SB_25_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U10 ( .a ({new_AGEMA_signal_1188, SB_24_n13}), .b ({new_AGEMA_signal_1034, SB_24_n12}), .c ({SubC_out_s1[56], SubC_out_s0[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U7 ( .a ({new_AGEMA_signal_1037, SB_24_T4}), .b ({new_AGEMA_signal_758, SB_24_T3}), .c ({new_AGEMA_signal_1188, SB_24_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_24_U2 ( .a ({new_AGEMA_signal_1036, SB_24_n9}), .b ({new_AGEMA_signal_1038, SB_24_T5}), .c ({SubC_out_s1[24], SubC_out_s0[24]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_24_t4_AND_U1 ( .a ({SubC_in_s1[56], SubC_in_s0[56]}), .b ({new_AGEMA_signal_758, SB_24_T3}), .clk (clk), .r (Fresh[142]), .c ({new_AGEMA_signal_1037, SB_24_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_24_t5_AND_U1 ( .a ({SubC_in_s1[56], SubC_in_s0[56]}), .b ({new_AGEMA_signal_757, SB_24_T2}), .clk (clk), .r (Fresh[143]), .c ({new_AGEMA_signal_1038, SB_24_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U10 ( .a ({new_AGEMA_signal_1192, SB_23_n13}), .b ({new_AGEMA_signal_1039, SB_23_n12}), .c ({SubC_out_s1[55], SubC_out_s0[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U7 ( .a ({new_AGEMA_signal_1042, SB_23_T4}), .b ({new_AGEMA_signal_768, SB_23_T3}), .c ({new_AGEMA_signal_1192, SB_23_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_23_U2 ( .a ({new_AGEMA_signal_1041, SB_23_n9}), .b ({new_AGEMA_signal_1043, SB_23_T5}), .c ({SubC_out_s1[23], SubC_out_s0[23]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_23_t4_AND_U1 ( .a ({SubC_in_s1[55], SubC_in_s0[55]}), .b ({new_AGEMA_signal_768, SB_23_T3}), .clk (clk), .r (Fresh[144]), .c ({new_AGEMA_signal_1042, SB_23_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_23_t5_AND_U1 ( .a ({SubC_in_s1[55], SubC_in_s0[55]}), .b ({new_AGEMA_signal_767, SB_23_T2}), .clk (clk), .r (Fresh[145]), .c ({new_AGEMA_signal_1043, SB_23_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U10 ( .a ({new_AGEMA_signal_1196, SB_22_n13}), .b ({new_AGEMA_signal_1044, SB_22_n12}), .c ({SubC_out_s1[54], SubC_out_s0[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U7 ( .a ({new_AGEMA_signal_1047, SB_22_T4}), .b ({new_AGEMA_signal_778, SB_22_T3}), .c ({new_AGEMA_signal_1196, SB_22_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_22_U2 ( .a ({new_AGEMA_signal_1046, SB_22_n9}), .b ({new_AGEMA_signal_1048, SB_22_T5}), .c ({SubC_out_s1[22], SubC_out_s0[22]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_22_t4_AND_U1 ( .a ({SubC_in_s1[54], SubC_in_s0[54]}), .b ({new_AGEMA_signal_778, SB_22_T3}), .clk (clk), .r (Fresh[146]), .c ({new_AGEMA_signal_1047, SB_22_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_22_t5_AND_U1 ( .a ({SubC_in_s1[54], SubC_in_s0[54]}), .b ({new_AGEMA_signal_777, SB_22_T2}), .clk (clk), .r (Fresh[147]), .c ({new_AGEMA_signal_1048, SB_22_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U10 ( .a ({new_AGEMA_signal_1200, SB_21_n13}), .b ({new_AGEMA_signal_1049, SB_21_n12}), .c ({SubC_out_s1[53], SubC_out_s0[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U7 ( .a ({new_AGEMA_signal_1052, SB_21_T4}), .b ({new_AGEMA_signal_788, SB_21_T3}), .c ({new_AGEMA_signal_1200, SB_21_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_21_U2 ( .a ({new_AGEMA_signal_1051, SB_21_n9}), .b ({new_AGEMA_signal_1053, SB_21_T5}), .c ({SubC_out_s1[21], SubC_out_s0[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_21_t4_AND_U1 ( .a ({SubC_in_s1[53], SubC_in_s0[53]}), .b ({new_AGEMA_signal_788, SB_21_T3}), .clk (clk), .r (Fresh[148]), .c ({new_AGEMA_signal_1052, SB_21_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_21_t5_AND_U1 ( .a ({SubC_in_s1[53], SubC_in_s0[53]}), .b ({new_AGEMA_signal_787, SB_21_T2}), .clk (clk), .r (Fresh[149]), .c ({new_AGEMA_signal_1053, SB_21_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U10 ( .a ({new_AGEMA_signal_1204, SB_20_n13}), .b ({new_AGEMA_signal_1054, SB_20_n12}), .c ({SubC_out_s1[52], SubC_out_s0[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U7 ( .a ({new_AGEMA_signal_1057, SB_20_T4}), .b ({new_AGEMA_signal_798, SB_20_T3}), .c ({new_AGEMA_signal_1204, SB_20_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_20_U2 ( .a ({new_AGEMA_signal_1056, SB_20_n9}), .b ({new_AGEMA_signal_1058, SB_20_T5}), .c ({SubC_out_s1[20], SubC_out_s0[20]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_20_t4_AND_U1 ( .a ({SubC_in_s1[52], SubC_in_s0[52]}), .b ({new_AGEMA_signal_798, SB_20_T3}), .clk (clk), .r (Fresh[150]), .c ({new_AGEMA_signal_1057, SB_20_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_20_t5_AND_U1 ( .a ({SubC_in_s1[52], SubC_in_s0[52]}), .b ({new_AGEMA_signal_797, SB_20_T2}), .clk (clk), .r (Fresh[151]), .c ({new_AGEMA_signal_1058, SB_20_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U10 ( .a ({new_AGEMA_signal_1208, SB_19_n13}), .b ({new_AGEMA_signal_1059, SB_19_n12}), .c ({SubC_out_s1[51], SubC_out_s0[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U7 ( .a ({new_AGEMA_signal_1062, SB_19_T4}), .b ({new_AGEMA_signal_808, SB_19_T3}), .c ({new_AGEMA_signal_1208, SB_19_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_19_U2 ( .a ({new_AGEMA_signal_1061, SB_19_n9}), .b ({new_AGEMA_signal_1063, SB_19_T5}), .c ({SubC_out_s1[19], SubC_out_s0[19]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_19_t4_AND_U1 ( .a ({SubC_in_s1[51], SubC_in_s0[51]}), .b ({new_AGEMA_signal_808, SB_19_T3}), .clk (clk), .r (Fresh[152]), .c ({new_AGEMA_signal_1062, SB_19_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_19_t5_AND_U1 ( .a ({SubC_in_s1[51], SubC_in_s0[51]}), .b ({new_AGEMA_signal_807, SB_19_T2}), .clk (clk), .r (Fresh[153]), .c ({new_AGEMA_signal_1063, SB_19_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U10 ( .a ({new_AGEMA_signal_1212, SB_18_n13}), .b ({new_AGEMA_signal_1064, SB_18_n12}), .c ({SubC_out_s1[50], SubC_out_s0[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U7 ( .a ({new_AGEMA_signal_1067, SB_18_T4}), .b ({new_AGEMA_signal_818, SB_18_T3}), .c ({new_AGEMA_signal_1212, SB_18_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_18_U2 ( .a ({new_AGEMA_signal_1066, SB_18_n9}), .b ({new_AGEMA_signal_1068, SB_18_T5}), .c ({SubC_out_s1[18], SubC_out_s0[18]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_18_t4_AND_U1 ( .a ({SubC_in_s1[50], SubC_in_s0[50]}), .b ({new_AGEMA_signal_818, SB_18_T3}), .clk (clk), .r (Fresh[154]), .c ({new_AGEMA_signal_1067, SB_18_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_18_t5_AND_U1 ( .a ({SubC_in_s1[50], SubC_in_s0[50]}), .b ({new_AGEMA_signal_817, SB_18_T2}), .clk (clk), .r (Fresh[155]), .c ({new_AGEMA_signal_1068, SB_18_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U10 ( .a ({new_AGEMA_signal_1216, SB_17_n13}), .b ({new_AGEMA_signal_1069, SB_17_n12}), .c ({SubC_out_s1[49], SubC_out_s0[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U7 ( .a ({new_AGEMA_signal_1072, SB_17_T4}), .b ({new_AGEMA_signal_828, SB_17_T3}), .c ({new_AGEMA_signal_1216, SB_17_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_17_U2 ( .a ({new_AGEMA_signal_1071, SB_17_n9}), .b ({new_AGEMA_signal_1073, SB_17_T5}), .c ({SubC_out_s1[17], SubC_out_s0[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_17_t4_AND_U1 ( .a ({SubC_in_s1[49], SubC_in_s0[49]}), .b ({new_AGEMA_signal_828, SB_17_T3}), .clk (clk), .r (Fresh[156]), .c ({new_AGEMA_signal_1072, SB_17_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_17_t5_AND_U1 ( .a ({SubC_in_s1[49], SubC_in_s0[49]}), .b ({new_AGEMA_signal_827, SB_17_T2}), .clk (clk), .r (Fresh[157]), .c ({new_AGEMA_signal_1073, SB_17_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U10 ( .a ({new_AGEMA_signal_1220, SB_16_n13}), .b ({new_AGEMA_signal_1074, SB_16_n12}), .c ({SubC_out_s1[48], SubC_out_s0[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U7 ( .a ({new_AGEMA_signal_1077, SB_16_T4}), .b ({new_AGEMA_signal_838, SB_16_T3}), .c ({new_AGEMA_signal_1220, SB_16_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_16_U2 ( .a ({new_AGEMA_signal_1076, SB_16_n9}), .b ({new_AGEMA_signal_1078, SB_16_T5}), .c ({SubC_out_s1[16], SubC_out_s0[16]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_16_t4_AND_U1 ( .a ({SubC_in_s1[48], SubC_in_s0[48]}), .b ({new_AGEMA_signal_838, SB_16_T3}), .clk (clk), .r (Fresh[158]), .c ({new_AGEMA_signal_1077, SB_16_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_16_t5_AND_U1 ( .a ({SubC_in_s1[48], SubC_in_s0[48]}), .b ({new_AGEMA_signal_837, SB_16_T2}), .clk (clk), .r (Fresh[159]), .c ({new_AGEMA_signal_1078, SB_16_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U10 ( .a ({new_AGEMA_signal_1224, SB_15_n13}), .b ({new_AGEMA_signal_1079, SB_15_n12}), .c ({SubC_out_s1[47], SubC_out_s0[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U7 ( .a ({new_AGEMA_signal_1082, SB_15_T4}), .b ({new_AGEMA_signal_848, SB_15_T3}), .c ({new_AGEMA_signal_1224, SB_15_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_15_U2 ( .a ({new_AGEMA_signal_1081, SB_15_n9}), .b ({new_AGEMA_signal_1083, SB_15_T5}), .c ({SubC_out_s1[15], SubC_out_s0[15]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_15_t4_AND_U1 ( .a ({SubC_in_s1[47], SubC_in_s0[47]}), .b ({new_AGEMA_signal_848, SB_15_T3}), .clk (clk), .r (Fresh[160]), .c ({new_AGEMA_signal_1082, SB_15_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_15_t5_AND_U1 ( .a ({SubC_in_s1[47], SubC_in_s0[47]}), .b ({new_AGEMA_signal_847, SB_15_T2}), .clk (clk), .r (Fresh[161]), .c ({new_AGEMA_signal_1083, SB_15_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U10 ( .a ({new_AGEMA_signal_1228, SB_14_n13}), .b ({new_AGEMA_signal_1084, SB_14_n12}), .c ({SubC_out_s1[46], SubC_out_s0[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U7 ( .a ({new_AGEMA_signal_1087, SB_14_T4}), .b ({new_AGEMA_signal_858, SB_14_T3}), .c ({new_AGEMA_signal_1228, SB_14_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_14_U2 ( .a ({new_AGEMA_signal_1086, SB_14_n9}), .b ({new_AGEMA_signal_1088, SB_14_T5}), .c ({SubC_out_s1[14], SubC_out_s0[14]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_14_t4_AND_U1 ( .a ({SubC_in_s1[46], SubC_in_s0[46]}), .b ({new_AGEMA_signal_858, SB_14_T3}), .clk (clk), .r (Fresh[162]), .c ({new_AGEMA_signal_1087, SB_14_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_14_t5_AND_U1 ( .a ({SubC_in_s1[46], SubC_in_s0[46]}), .b ({new_AGEMA_signal_857, SB_14_T2}), .clk (clk), .r (Fresh[163]), .c ({new_AGEMA_signal_1088, SB_14_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U10 ( .a ({new_AGEMA_signal_1232, SB_13_n13}), .b ({new_AGEMA_signal_1089, SB_13_n12}), .c ({SubC_out_s1[45], SubC_out_s0[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U7 ( .a ({new_AGEMA_signal_1092, SB_13_T4}), .b ({new_AGEMA_signal_868, SB_13_T3}), .c ({new_AGEMA_signal_1232, SB_13_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_13_U2 ( .a ({new_AGEMA_signal_1091, SB_13_n9}), .b ({new_AGEMA_signal_1093, SB_13_T5}), .c ({SubC_out_s1[13], SubC_out_s0[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_13_t4_AND_U1 ( .a ({SubC_in_s1[45], SubC_in_s0[45]}), .b ({new_AGEMA_signal_868, SB_13_T3}), .clk (clk), .r (Fresh[164]), .c ({new_AGEMA_signal_1092, SB_13_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_13_t5_AND_U1 ( .a ({SubC_in_s1[45], SubC_in_s0[45]}), .b ({new_AGEMA_signal_867, SB_13_T2}), .clk (clk), .r (Fresh[165]), .c ({new_AGEMA_signal_1093, SB_13_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U10 ( .a ({new_AGEMA_signal_1236, SB_12_n13}), .b ({new_AGEMA_signal_1094, SB_12_n12}), .c ({SubC_out_s1[44], SubC_out_s0[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U7 ( .a ({new_AGEMA_signal_1097, SB_12_T4}), .b ({new_AGEMA_signal_878, SB_12_T3}), .c ({new_AGEMA_signal_1236, SB_12_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_12_U2 ( .a ({new_AGEMA_signal_1096, SB_12_n9}), .b ({new_AGEMA_signal_1098, SB_12_T5}), .c ({SubC_out_s1[12], SubC_out_s0[12]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_12_t4_AND_U1 ( .a ({SubC_in_s1[44], SubC_in_s0[44]}), .b ({new_AGEMA_signal_878, SB_12_T3}), .clk (clk), .r (Fresh[166]), .c ({new_AGEMA_signal_1097, SB_12_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_12_t5_AND_U1 ( .a ({SubC_in_s1[44], SubC_in_s0[44]}), .b ({new_AGEMA_signal_877, SB_12_T2}), .clk (clk), .r (Fresh[167]), .c ({new_AGEMA_signal_1098, SB_12_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U10 ( .a ({new_AGEMA_signal_1240, SB_11_n13}), .b ({new_AGEMA_signal_1099, SB_11_n12}), .c ({SubC_out_s1[43], SubC_out_s0[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U7 ( .a ({new_AGEMA_signal_1102, SB_11_T4}), .b ({new_AGEMA_signal_888, SB_11_T3}), .c ({new_AGEMA_signal_1240, SB_11_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_11_U2 ( .a ({new_AGEMA_signal_1101, SB_11_n9}), .b ({new_AGEMA_signal_1103, SB_11_T5}), .c ({SubC_out_s1[11], SubC_out_s0[11]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_11_t4_AND_U1 ( .a ({SubC_in_s1[43], SubC_in_s0[43]}), .b ({new_AGEMA_signal_888, SB_11_T3}), .clk (clk), .r (Fresh[168]), .c ({new_AGEMA_signal_1102, SB_11_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_11_t5_AND_U1 ( .a ({SubC_in_s1[43], SubC_in_s0[43]}), .b ({new_AGEMA_signal_887, SB_11_T2}), .clk (clk), .r (Fresh[169]), .c ({new_AGEMA_signal_1103, SB_11_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U10 ( .a ({new_AGEMA_signal_1244, SB_10_n13}), .b ({new_AGEMA_signal_1104, SB_10_n12}), .c ({SubC_out_s1[42], SubC_out_s0[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U7 ( .a ({new_AGEMA_signal_1107, SB_10_T4}), .b ({new_AGEMA_signal_898, SB_10_T3}), .c ({new_AGEMA_signal_1244, SB_10_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_10_U2 ( .a ({new_AGEMA_signal_1106, SB_10_n9}), .b ({new_AGEMA_signal_1108, SB_10_T5}), .c ({SubC_out_s1[10], SubC_out_s0[10]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_10_t4_AND_U1 ( .a ({SubC_in_s1[42], SubC_in_s0[42]}), .b ({new_AGEMA_signal_898, SB_10_T3}), .clk (clk), .r (Fresh[170]), .c ({new_AGEMA_signal_1107, SB_10_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_10_t5_AND_U1 ( .a ({SubC_in_s1[42], SubC_in_s0[42]}), .b ({new_AGEMA_signal_897, SB_10_T2}), .clk (clk), .r (Fresh[171]), .c ({new_AGEMA_signal_1108, SB_10_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U10 ( .a ({new_AGEMA_signal_1248, SB_9_n13}), .b ({new_AGEMA_signal_1109, SB_9_n12}), .c ({SubC_out_s1[41], SubC_out_s0[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U7 ( .a ({new_AGEMA_signal_1112, SB_9_T4}), .b ({new_AGEMA_signal_908, SB_9_T3}), .c ({new_AGEMA_signal_1248, SB_9_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_9_U2 ( .a ({new_AGEMA_signal_1111, SB_9_n9}), .b ({new_AGEMA_signal_1113, SB_9_T5}), .c ({SubC_out_s1[9], SubC_out_s0[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_9_t4_AND_U1 ( .a ({SubC_in_s1[41], SubC_in_s0[41]}), .b ({new_AGEMA_signal_908, SB_9_T3}), .clk (clk), .r (Fresh[172]), .c ({new_AGEMA_signal_1112, SB_9_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_9_t5_AND_U1 ( .a ({SubC_in_s1[41], SubC_in_s0[41]}), .b ({new_AGEMA_signal_907, SB_9_T2}), .clk (clk), .r (Fresh[173]), .c ({new_AGEMA_signal_1113, SB_9_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U10 ( .a ({new_AGEMA_signal_1252, SB_8_n13}), .b ({new_AGEMA_signal_1114, SB_8_n12}), .c ({SubC_out_s1[40], SubC_out_s0[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U7 ( .a ({new_AGEMA_signal_1117, SB_8_T4}), .b ({new_AGEMA_signal_918, SB_8_T3}), .c ({new_AGEMA_signal_1252, SB_8_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_8_U2 ( .a ({new_AGEMA_signal_1116, SB_8_n9}), .b ({new_AGEMA_signal_1118, SB_8_T5}), .c ({SubC_out_s1[8], SubC_out_s0[8]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_8_t4_AND_U1 ( .a ({SubC_in_s1[40], SubC_in_s0[40]}), .b ({new_AGEMA_signal_918, SB_8_T3}), .clk (clk), .r (Fresh[174]), .c ({new_AGEMA_signal_1117, SB_8_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_8_t5_AND_U1 ( .a ({SubC_in_s1[40], SubC_in_s0[40]}), .b ({new_AGEMA_signal_917, SB_8_T2}), .clk (clk), .r (Fresh[175]), .c ({new_AGEMA_signal_1118, SB_8_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U10 ( .a ({new_AGEMA_signal_1256, SB_7_n13}), .b ({new_AGEMA_signal_1119, SB_7_n12}), .c ({SubC_out_s1[39], SubC_out_s0[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U7 ( .a ({new_AGEMA_signal_1122, SB_7_T4}), .b ({new_AGEMA_signal_928, SB_7_T3}), .c ({new_AGEMA_signal_1256, SB_7_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_7_U2 ( .a ({new_AGEMA_signal_1121, SB_7_n9}), .b ({new_AGEMA_signal_1123, SB_7_T5}), .c ({SubC_out_s1[7], SubC_out_s0[7]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_7_t4_AND_U1 ( .a ({SubC_in_s1[39], SubC_in_s0[39]}), .b ({new_AGEMA_signal_928, SB_7_T3}), .clk (clk), .r (Fresh[176]), .c ({new_AGEMA_signal_1122, SB_7_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_7_t5_AND_U1 ( .a ({SubC_in_s1[39], SubC_in_s0[39]}), .b ({new_AGEMA_signal_927, SB_7_T2}), .clk (clk), .r (Fresh[177]), .c ({new_AGEMA_signal_1123, SB_7_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U10 ( .a ({new_AGEMA_signal_1260, SB_6_n13}), .b ({new_AGEMA_signal_1124, SB_6_n12}), .c ({SubC_out_s1[38], SubC_out_s0[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U7 ( .a ({new_AGEMA_signal_1127, SB_6_T4}), .b ({new_AGEMA_signal_938, SB_6_T3}), .c ({new_AGEMA_signal_1260, SB_6_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_6_U2 ( .a ({new_AGEMA_signal_1126, SB_6_n9}), .b ({new_AGEMA_signal_1128, SB_6_T5}), .c ({SubC_out_s1[6], SubC_out_s0[6]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_6_t4_AND_U1 ( .a ({SubC_in_s1[38], SubC_in_s0[38]}), .b ({new_AGEMA_signal_938, SB_6_T3}), .clk (clk), .r (Fresh[178]), .c ({new_AGEMA_signal_1127, SB_6_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_6_t5_AND_U1 ( .a ({SubC_in_s1[38], SubC_in_s0[38]}), .b ({new_AGEMA_signal_937, SB_6_T2}), .clk (clk), .r (Fresh[179]), .c ({new_AGEMA_signal_1128, SB_6_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U10 ( .a ({new_AGEMA_signal_1264, SB_5_n13}), .b ({new_AGEMA_signal_1129, SB_5_n12}), .c ({SubC_out_s1[37], SubC_out_s0[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U7 ( .a ({new_AGEMA_signal_1132, SB_5_T4}), .b ({new_AGEMA_signal_948, SB_5_T3}), .c ({new_AGEMA_signal_1264, SB_5_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_5_U2 ( .a ({new_AGEMA_signal_1131, SB_5_n9}), .b ({new_AGEMA_signal_1133, SB_5_T5}), .c ({SubC_out_s1[5], SubC_out_s0[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_5_t4_AND_U1 ( .a ({SubC_in_s1[37], SubC_in_s0[37]}), .b ({new_AGEMA_signal_948, SB_5_T3}), .clk (clk), .r (Fresh[180]), .c ({new_AGEMA_signal_1132, SB_5_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_5_t5_AND_U1 ( .a ({SubC_in_s1[37], SubC_in_s0[37]}), .b ({new_AGEMA_signal_947, SB_5_T2}), .clk (clk), .r (Fresh[181]), .c ({new_AGEMA_signal_1133, SB_5_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U10 ( .a ({new_AGEMA_signal_1268, SB_4_n13}), .b ({new_AGEMA_signal_1134, SB_4_n12}), .c ({SubC_out_s1[36], SubC_out_s0[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U7 ( .a ({new_AGEMA_signal_1137, SB_4_T4}), .b ({new_AGEMA_signal_958, SB_4_T3}), .c ({new_AGEMA_signal_1268, SB_4_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_4_U2 ( .a ({new_AGEMA_signal_1136, SB_4_n9}), .b ({new_AGEMA_signal_1138, SB_4_T5}), .c ({SubC_out_s1[4], SubC_out_s0[4]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_4_t4_AND_U1 ( .a ({SubC_in_s1[36], SubC_in_s0[36]}), .b ({new_AGEMA_signal_958, SB_4_T3}), .clk (clk), .r (Fresh[182]), .c ({new_AGEMA_signal_1137, SB_4_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_4_t5_AND_U1 ( .a ({SubC_in_s1[36], SubC_in_s0[36]}), .b ({new_AGEMA_signal_957, SB_4_T2}), .clk (clk), .r (Fresh[183]), .c ({new_AGEMA_signal_1138, SB_4_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U10 ( .a ({new_AGEMA_signal_1272, SB_3_n13}), .b ({new_AGEMA_signal_1139, SB_3_n12}), .c ({SubC_out_s1[35], SubC_out_s0[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U7 ( .a ({new_AGEMA_signal_1142, SB_3_T4}), .b ({new_AGEMA_signal_968, SB_3_T3}), .c ({new_AGEMA_signal_1272, SB_3_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_3_U2 ( .a ({new_AGEMA_signal_1141, SB_3_n9}), .b ({new_AGEMA_signal_1143, SB_3_T5}), .c ({SubC_out_s1[3], SubC_out_s0[3]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_3_t4_AND_U1 ( .a ({SubC_in_s1[35], SubC_in_s0[35]}), .b ({new_AGEMA_signal_968, SB_3_T3}), .clk (clk), .r (Fresh[184]), .c ({new_AGEMA_signal_1142, SB_3_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_3_t5_AND_U1 ( .a ({SubC_in_s1[35], SubC_in_s0[35]}), .b ({new_AGEMA_signal_967, SB_3_T2}), .clk (clk), .r (Fresh[185]), .c ({new_AGEMA_signal_1143, SB_3_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U10 ( .a ({new_AGEMA_signal_1276, SB_2_n13}), .b ({new_AGEMA_signal_1144, SB_2_n12}), .c ({SubC_out_s1[34], SubC_out_s0[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U7 ( .a ({new_AGEMA_signal_1147, SB_2_T4}), .b ({new_AGEMA_signal_978, SB_2_T3}), .c ({new_AGEMA_signal_1276, SB_2_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_2_U2 ( .a ({new_AGEMA_signal_1146, SB_2_n9}), .b ({new_AGEMA_signal_1148, SB_2_T5}), .c ({SubC_out_s1[2], SubC_out_s0[2]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_2_t4_AND_U1 ( .a ({SubC_in_s1[34], SubC_in_s0[34]}), .b ({new_AGEMA_signal_978, SB_2_T3}), .clk (clk), .r (Fresh[186]), .c ({new_AGEMA_signal_1147, SB_2_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_2_t5_AND_U1 ( .a ({SubC_in_s1[34], SubC_in_s0[34]}), .b ({new_AGEMA_signal_977, SB_2_T2}), .clk (clk), .r (Fresh[187]), .c ({new_AGEMA_signal_1148, SB_2_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U10 ( .a ({new_AGEMA_signal_1280, SB_1_n13}), .b ({new_AGEMA_signal_1149, SB_1_n12}), .c ({SubC_out_s1[33], SubC_out_s0[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U7 ( .a ({new_AGEMA_signal_1152, SB_1_T4}), .b ({new_AGEMA_signal_988, SB_1_T3}), .c ({new_AGEMA_signal_1280, SB_1_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_1_U2 ( .a ({new_AGEMA_signal_1151, SB_1_n9}), .b ({new_AGEMA_signal_1153, SB_1_T5}), .c ({SubC_out_s1[1], SubC_out_s0[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_1_t4_AND_U1 ( .a ({SubC_in_s1[33], SubC_in_s0[33]}), .b ({new_AGEMA_signal_988, SB_1_T3}), .clk (clk), .r (Fresh[188]), .c ({new_AGEMA_signal_1152, SB_1_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_1_t5_AND_U1 ( .a ({SubC_in_s1[33], SubC_in_s0[33]}), .b ({new_AGEMA_signal_987, SB_1_T2}), .clk (clk), .r (Fresh[189]), .c ({new_AGEMA_signal_1153, SB_1_T5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U10 ( .a ({new_AGEMA_signal_1284, SB_0_n13}), .b ({new_AGEMA_signal_1154, SB_0_n12}), .c ({SubC_out_s1[32], SubC_out_s0[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U7 ( .a ({new_AGEMA_signal_1157, SB_0_T4}), .b ({new_AGEMA_signal_998, SB_0_T3}), .c ({new_AGEMA_signal_1284, SB_0_n13}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(0)) SB_0_U2 ( .a ({new_AGEMA_signal_1156, SB_0_n9}), .b ({new_AGEMA_signal_1158, SB_0_T5}), .c ({SubC_out_s1[0], SubC_out_s0[0]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_0_t4_AND_U1 ( .a ({SubC_in_s1[32], SubC_in_s0[32]}), .b ({new_AGEMA_signal_998, SB_0_T3}), .clk (clk), .r (Fresh[190]), .c ({new_AGEMA_signal_1157, SB_0_T4}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) SB_0_t5_AND_U1 ( .a ({SubC_in_s1[32], SubC_in_s0[32]}), .b ({new_AGEMA_signal_997, SB_0_T2}), .clk (clk), .r (Fresh[191]), .c ({new_AGEMA_signal_1158, SB_0_T5}) ) ;

endmodule
