/* modified netlist. Source: module Photon_256 in file ./test/Photon_256.v */
/* clock gating is added to the circuit, the latency increased 6 time(s)  */

module Photon_256_HPC2_ClockGating_d2 (w0_s0, w1_s0, temp_s0, k, p256_sel, clk, w0_s1, w0_s2, w1_s1, w1_s2, temp_s1, temp_s2, Fresh, /*rst,*/ y0_s0, y1_s0, temp_next_s0, temp_next_s1, temp_next_s2, y0_s1, y0_s2, y1_s1, y1_s2/*, Synch*/);
    input [127:0] w0_s0 ;
    input [127:0] w1_s0 ;
    input [127:0] temp_s0 ;
    input [3:0] k ;
    input p256_sel ;
    input clk ;
    input [127:0] w0_s1 ;
    input [127:0] w0_s2 ;
    input [127:0] w1_s1 ;
    input [127:0] w1_s2 ;
    input [127:0] temp_s1 ;
    input [127:0] temp_s2 ;
    //input rst ;
    input [3359:0] Fresh ;
    output [127:0] y0_s0 ;
    output [127:0] y1_s0 ;
    output [127:0] temp_next_s0 ;
    output [127:0] temp_next_s1 ;
    output [127:0] temp_next_s2 ;
    output [127:0] y0_s1 ;
    output [127:0] y0_s2 ;
    output [127:0] y1_s1 ;
    output [127:0] y1_s2 ;
    //output Synch ;
    wire add_sub1_0_n8 ;
    wire add_sub1_0_n7 ;
    wire add_sub1_0_n6 ;
    wire add_sub1_0_n5 ;
    wire add_sub1_0_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_0_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t0 ;
    wire add_sub1_1_n8 ;
    wire add_sub1_1_n7 ;
    wire add_sub1_1_n6 ;
    wire add_sub1_1_n5 ;
    wire add_sub1_1_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_1_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t0 ;
    wire add_sub1_2_n8 ;
    wire add_sub1_2_n7 ;
    wire add_sub1_2_n6 ;
    wire add_sub1_2_n5 ;
    wire add_sub1_2_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_2_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t0 ;
    wire add_sub1_3_n8 ;
    wire add_sub1_3_n7 ;
    wire add_sub1_3_n6 ;
    wire add_sub1_3_n5 ;
    wire add_sub1_3_addc_rom_ic_out_0_ ;
    wire add_sub1_3_addc_rom_ic_out_1_ ;
    wire add_sub1_3_addc_rom_ic_out_2_ ;
    wire add_sub1_3_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_3_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t0 ;
    wire mcs1_mcs_mat1_0_n128 ;
    wire mcs1_mcs_mat1_0_n127 ;
    wire mcs1_mcs_mat1_0_n126 ;
    wire mcs1_mcs_mat1_0_n125 ;
    wire mcs1_mcs_mat1_0_n124 ;
    wire mcs1_mcs_mat1_0_n123 ;
    wire mcs1_mcs_mat1_0_n122 ;
    wire mcs1_mcs_mat1_0_n121 ;
    wire mcs1_mcs_mat1_0_n120 ;
    wire mcs1_mcs_mat1_0_n119 ;
    wire mcs1_mcs_mat1_0_n118 ;
    wire mcs1_mcs_mat1_0_n117 ;
    wire mcs1_mcs_mat1_0_n116 ;
    wire mcs1_mcs_mat1_0_n115 ;
    wire mcs1_mcs_mat1_0_n114 ;
    wire mcs1_mcs_mat1_0_n113 ;
    wire mcs1_mcs_mat1_0_n112 ;
    wire mcs1_mcs_mat1_0_n111 ;
    wire mcs1_mcs_mat1_0_n110 ;
    wire mcs1_mcs_mat1_0_n109 ;
    wire mcs1_mcs_mat1_0_n108 ;
    wire mcs1_mcs_mat1_0_n107 ;
    wire mcs1_mcs_mat1_0_n106 ;
    wire mcs1_mcs_mat1_0_n105 ;
    wire mcs1_mcs_mat1_0_n104 ;
    wire mcs1_mcs_mat1_0_n103 ;
    wire mcs1_mcs_mat1_0_n102 ;
    wire mcs1_mcs_mat1_0_n101 ;
    wire mcs1_mcs_mat1_0_n100 ;
    wire mcs1_mcs_mat1_0_n99 ;
    wire mcs1_mcs_mat1_0_n98 ;
    wire mcs1_mcs_mat1_0_n97 ;
    wire mcs1_mcs_mat1_0_n96 ;
    wire mcs1_mcs_mat1_0_n95 ;
    wire mcs1_mcs_mat1_0_n94 ;
    wire mcs1_mcs_mat1_0_n93 ;
    wire mcs1_mcs_mat1_0_n92 ;
    wire mcs1_mcs_mat1_0_n91 ;
    wire mcs1_mcs_mat1_0_n90 ;
    wire mcs1_mcs_mat1_0_n89 ;
    wire mcs1_mcs_mat1_0_n88 ;
    wire mcs1_mcs_mat1_0_n87 ;
    wire mcs1_mcs_mat1_0_n86 ;
    wire mcs1_mcs_mat1_0_n85 ;
    wire mcs1_mcs_mat1_0_n84 ;
    wire mcs1_mcs_mat1_0_n83 ;
    wire mcs1_mcs_mat1_0_n82 ;
    wire mcs1_mcs_mat1_0_n81 ;
    wire mcs1_mcs_mat1_0_n80 ;
    wire mcs1_mcs_mat1_0_n79 ;
    wire mcs1_mcs_mat1_0_n78 ;
    wire mcs1_mcs_mat1_0_n77 ;
    wire mcs1_mcs_mat1_0_n76 ;
    wire mcs1_mcs_mat1_0_n75 ;
    wire mcs1_mcs_mat1_0_n74 ;
    wire mcs1_mcs_mat1_0_n73 ;
    wire mcs1_mcs_mat1_0_n72 ;
    wire mcs1_mcs_mat1_0_n71 ;
    wire mcs1_mcs_mat1_0_n70 ;
    wire mcs1_mcs_mat1_0_n69 ;
    wire mcs1_mcs_mat1_0_n68 ;
    wire mcs1_mcs_mat1_0_n67 ;
    wire mcs1_mcs_mat1_0_n66 ;
    wire mcs1_mcs_mat1_0_n65 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_1_n128 ;
    wire mcs1_mcs_mat1_1_n127 ;
    wire mcs1_mcs_mat1_1_n126 ;
    wire mcs1_mcs_mat1_1_n125 ;
    wire mcs1_mcs_mat1_1_n124 ;
    wire mcs1_mcs_mat1_1_n123 ;
    wire mcs1_mcs_mat1_1_n122 ;
    wire mcs1_mcs_mat1_1_n121 ;
    wire mcs1_mcs_mat1_1_n120 ;
    wire mcs1_mcs_mat1_1_n119 ;
    wire mcs1_mcs_mat1_1_n118 ;
    wire mcs1_mcs_mat1_1_n117 ;
    wire mcs1_mcs_mat1_1_n116 ;
    wire mcs1_mcs_mat1_1_n115 ;
    wire mcs1_mcs_mat1_1_n114 ;
    wire mcs1_mcs_mat1_1_n113 ;
    wire mcs1_mcs_mat1_1_n112 ;
    wire mcs1_mcs_mat1_1_n111 ;
    wire mcs1_mcs_mat1_1_n110 ;
    wire mcs1_mcs_mat1_1_n109 ;
    wire mcs1_mcs_mat1_1_n108 ;
    wire mcs1_mcs_mat1_1_n107 ;
    wire mcs1_mcs_mat1_1_n106 ;
    wire mcs1_mcs_mat1_1_n105 ;
    wire mcs1_mcs_mat1_1_n104 ;
    wire mcs1_mcs_mat1_1_n103 ;
    wire mcs1_mcs_mat1_1_n102 ;
    wire mcs1_mcs_mat1_1_n101 ;
    wire mcs1_mcs_mat1_1_n100 ;
    wire mcs1_mcs_mat1_1_n99 ;
    wire mcs1_mcs_mat1_1_n98 ;
    wire mcs1_mcs_mat1_1_n97 ;
    wire mcs1_mcs_mat1_1_n96 ;
    wire mcs1_mcs_mat1_1_n95 ;
    wire mcs1_mcs_mat1_1_n94 ;
    wire mcs1_mcs_mat1_1_n93 ;
    wire mcs1_mcs_mat1_1_n92 ;
    wire mcs1_mcs_mat1_1_n91 ;
    wire mcs1_mcs_mat1_1_n90 ;
    wire mcs1_mcs_mat1_1_n89 ;
    wire mcs1_mcs_mat1_1_n88 ;
    wire mcs1_mcs_mat1_1_n87 ;
    wire mcs1_mcs_mat1_1_n86 ;
    wire mcs1_mcs_mat1_1_n85 ;
    wire mcs1_mcs_mat1_1_n84 ;
    wire mcs1_mcs_mat1_1_n83 ;
    wire mcs1_mcs_mat1_1_n82 ;
    wire mcs1_mcs_mat1_1_n81 ;
    wire mcs1_mcs_mat1_1_n80 ;
    wire mcs1_mcs_mat1_1_n79 ;
    wire mcs1_mcs_mat1_1_n78 ;
    wire mcs1_mcs_mat1_1_n77 ;
    wire mcs1_mcs_mat1_1_n76 ;
    wire mcs1_mcs_mat1_1_n75 ;
    wire mcs1_mcs_mat1_1_n74 ;
    wire mcs1_mcs_mat1_1_n73 ;
    wire mcs1_mcs_mat1_1_n72 ;
    wire mcs1_mcs_mat1_1_n71 ;
    wire mcs1_mcs_mat1_1_n70 ;
    wire mcs1_mcs_mat1_1_n69 ;
    wire mcs1_mcs_mat1_1_n68 ;
    wire mcs1_mcs_mat1_1_n67 ;
    wire mcs1_mcs_mat1_1_n66 ;
    wire mcs1_mcs_mat1_1_n65 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_2_n128 ;
    wire mcs1_mcs_mat1_2_n127 ;
    wire mcs1_mcs_mat1_2_n126 ;
    wire mcs1_mcs_mat1_2_n125 ;
    wire mcs1_mcs_mat1_2_n124 ;
    wire mcs1_mcs_mat1_2_n123 ;
    wire mcs1_mcs_mat1_2_n122 ;
    wire mcs1_mcs_mat1_2_n121 ;
    wire mcs1_mcs_mat1_2_n120 ;
    wire mcs1_mcs_mat1_2_n119 ;
    wire mcs1_mcs_mat1_2_n118 ;
    wire mcs1_mcs_mat1_2_n117 ;
    wire mcs1_mcs_mat1_2_n116 ;
    wire mcs1_mcs_mat1_2_n115 ;
    wire mcs1_mcs_mat1_2_n114 ;
    wire mcs1_mcs_mat1_2_n113 ;
    wire mcs1_mcs_mat1_2_n112 ;
    wire mcs1_mcs_mat1_2_n111 ;
    wire mcs1_mcs_mat1_2_n110 ;
    wire mcs1_mcs_mat1_2_n109 ;
    wire mcs1_mcs_mat1_2_n108 ;
    wire mcs1_mcs_mat1_2_n107 ;
    wire mcs1_mcs_mat1_2_n106 ;
    wire mcs1_mcs_mat1_2_n105 ;
    wire mcs1_mcs_mat1_2_n104 ;
    wire mcs1_mcs_mat1_2_n103 ;
    wire mcs1_mcs_mat1_2_n102 ;
    wire mcs1_mcs_mat1_2_n101 ;
    wire mcs1_mcs_mat1_2_n100 ;
    wire mcs1_mcs_mat1_2_n99 ;
    wire mcs1_mcs_mat1_2_n98 ;
    wire mcs1_mcs_mat1_2_n97 ;
    wire mcs1_mcs_mat1_2_n96 ;
    wire mcs1_mcs_mat1_2_n95 ;
    wire mcs1_mcs_mat1_2_n94 ;
    wire mcs1_mcs_mat1_2_n93 ;
    wire mcs1_mcs_mat1_2_n92 ;
    wire mcs1_mcs_mat1_2_n91 ;
    wire mcs1_mcs_mat1_2_n90 ;
    wire mcs1_mcs_mat1_2_n89 ;
    wire mcs1_mcs_mat1_2_n88 ;
    wire mcs1_mcs_mat1_2_n87 ;
    wire mcs1_mcs_mat1_2_n86 ;
    wire mcs1_mcs_mat1_2_n85 ;
    wire mcs1_mcs_mat1_2_n84 ;
    wire mcs1_mcs_mat1_2_n83 ;
    wire mcs1_mcs_mat1_2_n82 ;
    wire mcs1_mcs_mat1_2_n81 ;
    wire mcs1_mcs_mat1_2_n80 ;
    wire mcs1_mcs_mat1_2_n79 ;
    wire mcs1_mcs_mat1_2_n78 ;
    wire mcs1_mcs_mat1_2_n77 ;
    wire mcs1_mcs_mat1_2_n76 ;
    wire mcs1_mcs_mat1_2_n75 ;
    wire mcs1_mcs_mat1_2_n74 ;
    wire mcs1_mcs_mat1_2_n73 ;
    wire mcs1_mcs_mat1_2_n72 ;
    wire mcs1_mcs_mat1_2_n71 ;
    wire mcs1_mcs_mat1_2_n70 ;
    wire mcs1_mcs_mat1_2_n69 ;
    wire mcs1_mcs_mat1_2_n68 ;
    wire mcs1_mcs_mat1_2_n67 ;
    wire mcs1_mcs_mat1_2_n66 ;
    wire mcs1_mcs_mat1_2_n65 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_3_n128 ;
    wire mcs1_mcs_mat1_3_n127 ;
    wire mcs1_mcs_mat1_3_n126 ;
    wire mcs1_mcs_mat1_3_n125 ;
    wire mcs1_mcs_mat1_3_n124 ;
    wire mcs1_mcs_mat1_3_n123 ;
    wire mcs1_mcs_mat1_3_n122 ;
    wire mcs1_mcs_mat1_3_n121 ;
    wire mcs1_mcs_mat1_3_n120 ;
    wire mcs1_mcs_mat1_3_n119 ;
    wire mcs1_mcs_mat1_3_n118 ;
    wire mcs1_mcs_mat1_3_n117 ;
    wire mcs1_mcs_mat1_3_n116 ;
    wire mcs1_mcs_mat1_3_n115 ;
    wire mcs1_mcs_mat1_3_n114 ;
    wire mcs1_mcs_mat1_3_n113 ;
    wire mcs1_mcs_mat1_3_n112 ;
    wire mcs1_mcs_mat1_3_n111 ;
    wire mcs1_mcs_mat1_3_n110 ;
    wire mcs1_mcs_mat1_3_n109 ;
    wire mcs1_mcs_mat1_3_n108 ;
    wire mcs1_mcs_mat1_3_n107 ;
    wire mcs1_mcs_mat1_3_n106 ;
    wire mcs1_mcs_mat1_3_n105 ;
    wire mcs1_mcs_mat1_3_n104 ;
    wire mcs1_mcs_mat1_3_n103 ;
    wire mcs1_mcs_mat1_3_n102 ;
    wire mcs1_mcs_mat1_3_n101 ;
    wire mcs1_mcs_mat1_3_n100 ;
    wire mcs1_mcs_mat1_3_n99 ;
    wire mcs1_mcs_mat1_3_n98 ;
    wire mcs1_mcs_mat1_3_n97 ;
    wire mcs1_mcs_mat1_3_n96 ;
    wire mcs1_mcs_mat1_3_n95 ;
    wire mcs1_mcs_mat1_3_n94 ;
    wire mcs1_mcs_mat1_3_n93 ;
    wire mcs1_mcs_mat1_3_n92 ;
    wire mcs1_mcs_mat1_3_n91 ;
    wire mcs1_mcs_mat1_3_n90 ;
    wire mcs1_mcs_mat1_3_n89 ;
    wire mcs1_mcs_mat1_3_n88 ;
    wire mcs1_mcs_mat1_3_n87 ;
    wire mcs1_mcs_mat1_3_n86 ;
    wire mcs1_mcs_mat1_3_n85 ;
    wire mcs1_mcs_mat1_3_n84 ;
    wire mcs1_mcs_mat1_3_n83 ;
    wire mcs1_mcs_mat1_3_n82 ;
    wire mcs1_mcs_mat1_3_n81 ;
    wire mcs1_mcs_mat1_3_n80 ;
    wire mcs1_mcs_mat1_3_n79 ;
    wire mcs1_mcs_mat1_3_n78 ;
    wire mcs1_mcs_mat1_3_n77 ;
    wire mcs1_mcs_mat1_3_n76 ;
    wire mcs1_mcs_mat1_3_n75 ;
    wire mcs1_mcs_mat1_3_n74 ;
    wire mcs1_mcs_mat1_3_n73 ;
    wire mcs1_mcs_mat1_3_n72 ;
    wire mcs1_mcs_mat1_3_n71 ;
    wire mcs1_mcs_mat1_3_n70 ;
    wire mcs1_mcs_mat1_3_n69 ;
    wire mcs1_mcs_mat1_3_n68 ;
    wire mcs1_mcs_mat1_3_n67 ;
    wire mcs1_mcs_mat1_3_n66 ;
    wire mcs1_mcs_mat1_3_n65 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_4_n128 ;
    wire mcs1_mcs_mat1_4_n127 ;
    wire mcs1_mcs_mat1_4_n126 ;
    wire mcs1_mcs_mat1_4_n125 ;
    wire mcs1_mcs_mat1_4_n124 ;
    wire mcs1_mcs_mat1_4_n123 ;
    wire mcs1_mcs_mat1_4_n122 ;
    wire mcs1_mcs_mat1_4_n121 ;
    wire mcs1_mcs_mat1_4_n120 ;
    wire mcs1_mcs_mat1_4_n119 ;
    wire mcs1_mcs_mat1_4_n118 ;
    wire mcs1_mcs_mat1_4_n117 ;
    wire mcs1_mcs_mat1_4_n116 ;
    wire mcs1_mcs_mat1_4_n115 ;
    wire mcs1_mcs_mat1_4_n114 ;
    wire mcs1_mcs_mat1_4_n113 ;
    wire mcs1_mcs_mat1_4_n112 ;
    wire mcs1_mcs_mat1_4_n111 ;
    wire mcs1_mcs_mat1_4_n110 ;
    wire mcs1_mcs_mat1_4_n109 ;
    wire mcs1_mcs_mat1_4_n108 ;
    wire mcs1_mcs_mat1_4_n107 ;
    wire mcs1_mcs_mat1_4_n106 ;
    wire mcs1_mcs_mat1_4_n105 ;
    wire mcs1_mcs_mat1_4_n104 ;
    wire mcs1_mcs_mat1_4_n103 ;
    wire mcs1_mcs_mat1_4_n102 ;
    wire mcs1_mcs_mat1_4_n101 ;
    wire mcs1_mcs_mat1_4_n100 ;
    wire mcs1_mcs_mat1_4_n99 ;
    wire mcs1_mcs_mat1_4_n98 ;
    wire mcs1_mcs_mat1_4_n97 ;
    wire mcs1_mcs_mat1_4_n96 ;
    wire mcs1_mcs_mat1_4_n95 ;
    wire mcs1_mcs_mat1_4_n94 ;
    wire mcs1_mcs_mat1_4_n93 ;
    wire mcs1_mcs_mat1_4_n92 ;
    wire mcs1_mcs_mat1_4_n91 ;
    wire mcs1_mcs_mat1_4_n90 ;
    wire mcs1_mcs_mat1_4_n89 ;
    wire mcs1_mcs_mat1_4_n88 ;
    wire mcs1_mcs_mat1_4_n87 ;
    wire mcs1_mcs_mat1_4_n86 ;
    wire mcs1_mcs_mat1_4_n85 ;
    wire mcs1_mcs_mat1_4_n84 ;
    wire mcs1_mcs_mat1_4_n83 ;
    wire mcs1_mcs_mat1_4_n82 ;
    wire mcs1_mcs_mat1_4_n81 ;
    wire mcs1_mcs_mat1_4_n80 ;
    wire mcs1_mcs_mat1_4_n79 ;
    wire mcs1_mcs_mat1_4_n78 ;
    wire mcs1_mcs_mat1_4_n77 ;
    wire mcs1_mcs_mat1_4_n76 ;
    wire mcs1_mcs_mat1_4_n75 ;
    wire mcs1_mcs_mat1_4_n74 ;
    wire mcs1_mcs_mat1_4_n73 ;
    wire mcs1_mcs_mat1_4_n72 ;
    wire mcs1_mcs_mat1_4_n71 ;
    wire mcs1_mcs_mat1_4_n70 ;
    wire mcs1_mcs_mat1_4_n69 ;
    wire mcs1_mcs_mat1_4_n68 ;
    wire mcs1_mcs_mat1_4_n67 ;
    wire mcs1_mcs_mat1_4_n66 ;
    wire mcs1_mcs_mat1_4_n65 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_5_n128 ;
    wire mcs1_mcs_mat1_5_n127 ;
    wire mcs1_mcs_mat1_5_n126 ;
    wire mcs1_mcs_mat1_5_n125 ;
    wire mcs1_mcs_mat1_5_n124 ;
    wire mcs1_mcs_mat1_5_n123 ;
    wire mcs1_mcs_mat1_5_n122 ;
    wire mcs1_mcs_mat1_5_n121 ;
    wire mcs1_mcs_mat1_5_n120 ;
    wire mcs1_mcs_mat1_5_n119 ;
    wire mcs1_mcs_mat1_5_n118 ;
    wire mcs1_mcs_mat1_5_n117 ;
    wire mcs1_mcs_mat1_5_n116 ;
    wire mcs1_mcs_mat1_5_n115 ;
    wire mcs1_mcs_mat1_5_n114 ;
    wire mcs1_mcs_mat1_5_n113 ;
    wire mcs1_mcs_mat1_5_n112 ;
    wire mcs1_mcs_mat1_5_n111 ;
    wire mcs1_mcs_mat1_5_n110 ;
    wire mcs1_mcs_mat1_5_n109 ;
    wire mcs1_mcs_mat1_5_n108 ;
    wire mcs1_mcs_mat1_5_n107 ;
    wire mcs1_mcs_mat1_5_n106 ;
    wire mcs1_mcs_mat1_5_n105 ;
    wire mcs1_mcs_mat1_5_n104 ;
    wire mcs1_mcs_mat1_5_n103 ;
    wire mcs1_mcs_mat1_5_n102 ;
    wire mcs1_mcs_mat1_5_n101 ;
    wire mcs1_mcs_mat1_5_n100 ;
    wire mcs1_mcs_mat1_5_n99 ;
    wire mcs1_mcs_mat1_5_n98 ;
    wire mcs1_mcs_mat1_5_n97 ;
    wire mcs1_mcs_mat1_5_n96 ;
    wire mcs1_mcs_mat1_5_n95 ;
    wire mcs1_mcs_mat1_5_n94 ;
    wire mcs1_mcs_mat1_5_n93 ;
    wire mcs1_mcs_mat1_5_n92 ;
    wire mcs1_mcs_mat1_5_n91 ;
    wire mcs1_mcs_mat1_5_n90 ;
    wire mcs1_mcs_mat1_5_n89 ;
    wire mcs1_mcs_mat1_5_n88 ;
    wire mcs1_mcs_mat1_5_n87 ;
    wire mcs1_mcs_mat1_5_n86 ;
    wire mcs1_mcs_mat1_5_n85 ;
    wire mcs1_mcs_mat1_5_n84 ;
    wire mcs1_mcs_mat1_5_n83 ;
    wire mcs1_mcs_mat1_5_n82 ;
    wire mcs1_mcs_mat1_5_n81 ;
    wire mcs1_mcs_mat1_5_n80 ;
    wire mcs1_mcs_mat1_5_n79 ;
    wire mcs1_mcs_mat1_5_n78 ;
    wire mcs1_mcs_mat1_5_n77 ;
    wire mcs1_mcs_mat1_5_n76 ;
    wire mcs1_mcs_mat1_5_n75 ;
    wire mcs1_mcs_mat1_5_n74 ;
    wire mcs1_mcs_mat1_5_n73 ;
    wire mcs1_mcs_mat1_5_n72 ;
    wire mcs1_mcs_mat1_5_n71 ;
    wire mcs1_mcs_mat1_5_n70 ;
    wire mcs1_mcs_mat1_5_n69 ;
    wire mcs1_mcs_mat1_5_n68 ;
    wire mcs1_mcs_mat1_5_n67 ;
    wire mcs1_mcs_mat1_5_n66 ;
    wire mcs1_mcs_mat1_5_n65 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_6_n128 ;
    wire mcs1_mcs_mat1_6_n127 ;
    wire mcs1_mcs_mat1_6_n126 ;
    wire mcs1_mcs_mat1_6_n125 ;
    wire mcs1_mcs_mat1_6_n124 ;
    wire mcs1_mcs_mat1_6_n123 ;
    wire mcs1_mcs_mat1_6_n122 ;
    wire mcs1_mcs_mat1_6_n121 ;
    wire mcs1_mcs_mat1_6_n120 ;
    wire mcs1_mcs_mat1_6_n119 ;
    wire mcs1_mcs_mat1_6_n118 ;
    wire mcs1_mcs_mat1_6_n117 ;
    wire mcs1_mcs_mat1_6_n116 ;
    wire mcs1_mcs_mat1_6_n115 ;
    wire mcs1_mcs_mat1_6_n114 ;
    wire mcs1_mcs_mat1_6_n113 ;
    wire mcs1_mcs_mat1_6_n112 ;
    wire mcs1_mcs_mat1_6_n111 ;
    wire mcs1_mcs_mat1_6_n110 ;
    wire mcs1_mcs_mat1_6_n109 ;
    wire mcs1_mcs_mat1_6_n108 ;
    wire mcs1_mcs_mat1_6_n107 ;
    wire mcs1_mcs_mat1_6_n106 ;
    wire mcs1_mcs_mat1_6_n105 ;
    wire mcs1_mcs_mat1_6_n104 ;
    wire mcs1_mcs_mat1_6_n103 ;
    wire mcs1_mcs_mat1_6_n102 ;
    wire mcs1_mcs_mat1_6_n101 ;
    wire mcs1_mcs_mat1_6_n100 ;
    wire mcs1_mcs_mat1_6_n99 ;
    wire mcs1_mcs_mat1_6_n98 ;
    wire mcs1_mcs_mat1_6_n97 ;
    wire mcs1_mcs_mat1_6_n96 ;
    wire mcs1_mcs_mat1_6_n95 ;
    wire mcs1_mcs_mat1_6_n94 ;
    wire mcs1_mcs_mat1_6_n93 ;
    wire mcs1_mcs_mat1_6_n92 ;
    wire mcs1_mcs_mat1_6_n91 ;
    wire mcs1_mcs_mat1_6_n90 ;
    wire mcs1_mcs_mat1_6_n89 ;
    wire mcs1_mcs_mat1_6_n88 ;
    wire mcs1_mcs_mat1_6_n87 ;
    wire mcs1_mcs_mat1_6_n86 ;
    wire mcs1_mcs_mat1_6_n85 ;
    wire mcs1_mcs_mat1_6_n84 ;
    wire mcs1_mcs_mat1_6_n83 ;
    wire mcs1_mcs_mat1_6_n82 ;
    wire mcs1_mcs_mat1_6_n81 ;
    wire mcs1_mcs_mat1_6_n80 ;
    wire mcs1_mcs_mat1_6_n79 ;
    wire mcs1_mcs_mat1_6_n78 ;
    wire mcs1_mcs_mat1_6_n77 ;
    wire mcs1_mcs_mat1_6_n76 ;
    wire mcs1_mcs_mat1_6_n75 ;
    wire mcs1_mcs_mat1_6_n74 ;
    wire mcs1_mcs_mat1_6_n73 ;
    wire mcs1_mcs_mat1_6_n72 ;
    wire mcs1_mcs_mat1_6_n71 ;
    wire mcs1_mcs_mat1_6_n70 ;
    wire mcs1_mcs_mat1_6_n69 ;
    wire mcs1_mcs_mat1_6_n68 ;
    wire mcs1_mcs_mat1_6_n67 ;
    wire mcs1_mcs_mat1_6_n66 ;
    wire mcs1_mcs_mat1_6_n65 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_7_n128 ;
    wire mcs1_mcs_mat1_7_n127 ;
    wire mcs1_mcs_mat1_7_n126 ;
    wire mcs1_mcs_mat1_7_n125 ;
    wire mcs1_mcs_mat1_7_n124 ;
    wire mcs1_mcs_mat1_7_n123 ;
    wire mcs1_mcs_mat1_7_n122 ;
    wire mcs1_mcs_mat1_7_n121 ;
    wire mcs1_mcs_mat1_7_n120 ;
    wire mcs1_mcs_mat1_7_n119 ;
    wire mcs1_mcs_mat1_7_n118 ;
    wire mcs1_mcs_mat1_7_n117 ;
    wire mcs1_mcs_mat1_7_n116 ;
    wire mcs1_mcs_mat1_7_n115 ;
    wire mcs1_mcs_mat1_7_n114 ;
    wire mcs1_mcs_mat1_7_n113 ;
    wire mcs1_mcs_mat1_7_n112 ;
    wire mcs1_mcs_mat1_7_n111 ;
    wire mcs1_mcs_mat1_7_n110 ;
    wire mcs1_mcs_mat1_7_n109 ;
    wire mcs1_mcs_mat1_7_n108 ;
    wire mcs1_mcs_mat1_7_n107 ;
    wire mcs1_mcs_mat1_7_n106 ;
    wire mcs1_mcs_mat1_7_n105 ;
    wire mcs1_mcs_mat1_7_n104 ;
    wire mcs1_mcs_mat1_7_n103 ;
    wire mcs1_mcs_mat1_7_n102 ;
    wire mcs1_mcs_mat1_7_n101 ;
    wire mcs1_mcs_mat1_7_n100 ;
    wire mcs1_mcs_mat1_7_n99 ;
    wire mcs1_mcs_mat1_7_n98 ;
    wire mcs1_mcs_mat1_7_n97 ;
    wire mcs1_mcs_mat1_7_n96 ;
    wire mcs1_mcs_mat1_7_n95 ;
    wire mcs1_mcs_mat1_7_n94 ;
    wire mcs1_mcs_mat1_7_n93 ;
    wire mcs1_mcs_mat1_7_n92 ;
    wire mcs1_mcs_mat1_7_n91 ;
    wire mcs1_mcs_mat1_7_n90 ;
    wire mcs1_mcs_mat1_7_n89 ;
    wire mcs1_mcs_mat1_7_n88 ;
    wire mcs1_mcs_mat1_7_n87 ;
    wire mcs1_mcs_mat1_7_n86 ;
    wire mcs1_mcs_mat1_7_n85 ;
    wire mcs1_mcs_mat1_7_n84 ;
    wire mcs1_mcs_mat1_7_n83 ;
    wire mcs1_mcs_mat1_7_n82 ;
    wire mcs1_mcs_mat1_7_n81 ;
    wire mcs1_mcs_mat1_7_n80 ;
    wire mcs1_mcs_mat1_7_n79 ;
    wire mcs1_mcs_mat1_7_n78 ;
    wire mcs1_mcs_mat1_7_n77 ;
    wire mcs1_mcs_mat1_7_n76 ;
    wire mcs1_mcs_mat1_7_n75 ;
    wire mcs1_mcs_mat1_7_n74 ;
    wire mcs1_mcs_mat1_7_n73 ;
    wire mcs1_mcs_mat1_7_n72 ;
    wire mcs1_mcs_mat1_7_n71 ;
    wire mcs1_mcs_mat1_7_n70 ;
    wire mcs1_mcs_mat1_7_n69 ;
    wire mcs1_mcs_mat1_7_n68 ;
    wire mcs1_mcs_mat1_7_n67 ;
    wire mcs1_mcs_mat1_7_n66 ;
    wire mcs1_mcs_mat1_7_n65 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x0x4 ;
    wire [127:0] addc_in ;
    wire [127:0] subc_out ;
    wire [124:1] shiftr_out ;
    wire [255:128] mcs_out ;
    wire [127:0] y0_1 ;
    wire [3:0] add_sub1_0_addc_out ;
    wire [2:0] add_sub1_0_addc_rom_ic_out ;
    wire [3:0] add_sub1_0_addc_rom_rc_out ;
    wire [3:0] add_sub1_1_addc_out ;
    wire [2:0] add_sub1_1_addc_rom_ic_out ;
    wire [3:0] add_sub1_1_addc_rom_rc_out ;
    wire [3:0] add_sub1_2_addc_out ;
    wire [2:0] add_sub1_2_addc_rom_ic_out ;
    wire [3:0] add_sub1_2_addc_rom_rc_out ;
    wire [3:0] add_sub1_3_addc_out ;
    wire [3:0] add_sub1_3_addc_rom_rc_out ;
    wire [127:0] mcs1_mcs_mat1_0_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_1_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_2_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_3_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_4_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_5_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_6_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_7_mcs_out ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10778 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10793 ;
    wire new_AGEMA_signal_10794 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10797 ;
    wire new_AGEMA_signal_10798 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10801 ;
    wire new_AGEMA_signal_10802 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10805 ;
    wire new_AGEMA_signal_10806 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10809 ;
    wire new_AGEMA_signal_10810 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10813 ;
    wire new_AGEMA_signal_10814 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10817 ;
    wire new_AGEMA_signal_10818 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10821 ;
    wire new_AGEMA_signal_10822 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10825 ;
    wire new_AGEMA_signal_10826 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10829 ;
    wire new_AGEMA_signal_10830 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10833 ;
    wire new_AGEMA_signal_10834 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10837 ;
    wire new_AGEMA_signal_10838 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10841 ;
    wire new_AGEMA_signal_10842 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10845 ;
    wire new_AGEMA_signal_10846 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10849 ;
    wire new_AGEMA_signal_10850 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10853 ;
    wire new_AGEMA_signal_10854 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10857 ;
    wire new_AGEMA_signal_10858 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10861 ;
    wire new_AGEMA_signal_10862 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10865 ;
    wire new_AGEMA_signal_10866 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10874 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11197 ;
    wire new_AGEMA_signal_11198 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11201 ;
    wire new_AGEMA_signal_11202 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11205 ;
    wire new_AGEMA_signal_11206 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11209 ;
    wire new_AGEMA_signal_11210 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11213 ;
    wire new_AGEMA_signal_11214 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11217 ;
    wire new_AGEMA_signal_11218 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11221 ;
    wire new_AGEMA_signal_11222 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11225 ;
    wire new_AGEMA_signal_11226 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11229 ;
    wire new_AGEMA_signal_11230 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11233 ;
    wire new_AGEMA_signal_11234 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11237 ;
    wire new_AGEMA_signal_11238 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11241 ;
    wire new_AGEMA_signal_11242 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11245 ;
    wire new_AGEMA_signal_11246 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11249 ;
    wire new_AGEMA_signal_11250 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11253 ;
    wire new_AGEMA_signal_11254 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11257 ;
    wire new_AGEMA_signal_11258 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11261 ;
    wire new_AGEMA_signal_11262 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11265 ;
    wire new_AGEMA_signal_11266 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11269 ;
    wire new_AGEMA_signal_11270 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11273 ;
    wire new_AGEMA_signal_11274 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11277 ;
    wire new_AGEMA_signal_11278 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11281 ;
    wire new_AGEMA_signal_11282 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11285 ;
    wire new_AGEMA_signal_11286 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11289 ;
    wire new_AGEMA_signal_11290 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11293 ;
    wire new_AGEMA_signal_11294 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11297 ;
    wire new_AGEMA_signal_11298 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11301 ;
    wire new_AGEMA_signal_11302 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11305 ;
    wire new_AGEMA_signal_11306 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11309 ;
    wire new_AGEMA_signal_11310 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11313 ;
    wire new_AGEMA_signal_11314 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11317 ;
    wire new_AGEMA_signal_11318 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11321 ;
    wire new_AGEMA_signal_11322 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11645 ;
    wire new_AGEMA_signal_11646 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11649 ;
    wire new_AGEMA_signal_11650 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11653 ;
    wire new_AGEMA_signal_11654 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11657 ;
    wire new_AGEMA_signal_11658 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11661 ;
    wire new_AGEMA_signal_11662 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11665 ;
    wire new_AGEMA_signal_11666 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11669 ;
    wire new_AGEMA_signal_11670 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11673 ;
    wire new_AGEMA_signal_11674 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11677 ;
    wire new_AGEMA_signal_11678 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11681 ;
    wire new_AGEMA_signal_11682 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11685 ;
    wire new_AGEMA_signal_11686 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11689 ;
    wire new_AGEMA_signal_11690 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11693 ;
    wire new_AGEMA_signal_11694 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11697 ;
    wire new_AGEMA_signal_11698 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11701 ;
    wire new_AGEMA_signal_11702 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11705 ;
    wire new_AGEMA_signal_11706 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11709 ;
    wire new_AGEMA_signal_11710 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11713 ;
    wire new_AGEMA_signal_11714 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11717 ;
    wire new_AGEMA_signal_11718 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11721 ;
    wire new_AGEMA_signal_11722 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11725 ;
    wire new_AGEMA_signal_11726 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11729 ;
    wire new_AGEMA_signal_11730 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11733 ;
    wire new_AGEMA_signal_11734 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11737 ;
    wire new_AGEMA_signal_11738 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11741 ;
    wire new_AGEMA_signal_11742 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11745 ;
    wire new_AGEMA_signal_11746 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11749 ;
    wire new_AGEMA_signal_11750 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11753 ;
    wire new_AGEMA_signal_11754 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11757 ;
    wire new_AGEMA_signal_11758 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11761 ;
    wire new_AGEMA_signal_11762 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11765 ;
    wire new_AGEMA_signal_11766 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11769 ;
    wire new_AGEMA_signal_11770 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12087 ;
    wire new_AGEMA_signal_12088 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12091 ;
    wire new_AGEMA_signal_12092 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12095 ;
    wire new_AGEMA_signal_12096 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12099 ;
    wire new_AGEMA_signal_12100 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12103 ;
    wire new_AGEMA_signal_12104 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12107 ;
    wire new_AGEMA_signal_12108 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12111 ;
    wire new_AGEMA_signal_12112 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12115 ;
    wire new_AGEMA_signal_12116 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12119 ;
    wire new_AGEMA_signal_12120 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12123 ;
    wire new_AGEMA_signal_12124 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12127 ;
    wire new_AGEMA_signal_12128 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12131 ;
    wire new_AGEMA_signal_12132 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12135 ;
    wire new_AGEMA_signal_12136 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12139 ;
    wire new_AGEMA_signal_12140 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12143 ;
    wire new_AGEMA_signal_12144 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12147 ;
    wire new_AGEMA_signal_12148 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12151 ;
    wire new_AGEMA_signal_12152 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12155 ;
    wire new_AGEMA_signal_12156 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12159 ;
    wire new_AGEMA_signal_12160 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12163 ;
    wire new_AGEMA_signal_12164 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12167 ;
    wire new_AGEMA_signal_12168 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12171 ;
    wire new_AGEMA_signal_12172 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12175 ;
    wire new_AGEMA_signal_12176 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12179 ;
    wire new_AGEMA_signal_12180 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12183 ;
    wire new_AGEMA_signal_12184 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12187 ;
    wire new_AGEMA_signal_12188 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12191 ;
    wire new_AGEMA_signal_12192 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12195 ;
    wire new_AGEMA_signal_12196 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12199 ;
    wire new_AGEMA_signal_12200 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12313 ;
    wire new_AGEMA_signal_12314 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12317 ;
    wire new_AGEMA_signal_12318 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12321 ;
    wire new_AGEMA_signal_12322 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12325 ;
    wire new_AGEMA_signal_12326 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12329 ;
    wire new_AGEMA_signal_12330 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12333 ;
    wire new_AGEMA_signal_12334 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12337 ;
    wire new_AGEMA_signal_12338 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12341 ;
    wire new_AGEMA_signal_12342 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12345 ;
    wire new_AGEMA_signal_12346 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12349 ;
    wire new_AGEMA_signal_12350 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12353 ;
    wire new_AGEMA_signal_12354 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12357 ;
    wire new_AGEMA_signal_12358 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12361 ;
    wire new_AGEMA_signal_12362 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12365 ;
    wire new_AGEMA_signal_12366 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12369 ;
    wire new_AGEMA_signal_12370 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12373 ;
    wire new_AGEMA_signal_12374 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12377 ;
    wire new_AGEMA_signal_12378 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12381 ;
    wire new_AGEMA_signal_12382 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12385 ;
    wire new_AGEMA_signal_12386 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12389 ;
    wire new_AGEMA_signal_12390 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12393 ;
    wire new_AGEMA_signal_12394 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12397 ;
    wire new_AGEMA_signal_12398 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12401 ;
    wire new_AGEMA_signal_12402 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12405 ;
    wire new_AGEMA_signal_12406 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12409 ;
    wire new_AGEMA_signal_12410 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12413 ;
    wire new_AGEMA_signal_12414 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12417 ;
    wire new_AGEMA_signal_12418 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12421 ;
    wire new_AGEMA_signal_12422 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12425 ;
    wire new_AGEMA_signal_12426 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12429 ;
    wire new_AGEMA_signal_12430 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12433 ;
    wire new_AGEMA_signal_12434 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12437 ;
    wire new_AGEMA_signal_12438 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12441 ;
    wire new_AGEMA_signal_12442 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12445 ;
    wire new_AGEMA_signal_12446 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12449 ;
    wire new_AGEMA_signal_12450 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12453 ;
    wire new_AGEMA_signal_12454 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12457 ;
    wire new_AGEMA_signal_12458 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12461 ;
    wire new_AGEMA_signal_12462 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12465 ;
    wire new_AGEMA_signal_12466 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12469 ;
    wire new_AGEMA_signal_12470 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12473 ;
    wire new_AGEMA_signal_12474 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12477 ;
    wire new_AGEMA_signal_12478 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12481 ;
    wire new_AGEMA_signal_12482 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12485 ;
    wire new_AGEMA_signal_12486 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12489 ;
    wire new_AGEMA_signal_12490 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12493 ;
    wire new_AGEMA_signal_12494 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12497 ;
    wire new_AGEMA_signal_12498 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12501 ;
    wire new_AGEMA_signal_12502 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12505 ;
    wire new_AGEMA_signal_12506 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12509 ;
    wire new_AGEMA_signal_12510 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12513 ;
    wire new_AGEMA_signal_12514 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12517 ;
    wire new_AGEMA_signal_12518 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12521 ;
    wire new_AGEMA_signal_12522 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12525 ;
    wire new_AGEMA_signal_12526 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12529 ;
    wire new_AGEMA_signal_12530 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12533 ;
    wire new_AGEMA_signal_12534 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12537 ;
    wire new_AGEMA_signal_12538 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12541 ;
    wire new_AGEMA_signal_12542 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12545 ;
    wire new_AGEMA_signal_12546 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12549 ;
    wire new_AGEMA_signal_12550 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12553 ;
    wire new_AGEMA_signal_12554 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12557 ;
    wire new_AGEMA_signal_12558 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12561 ;
    wire new_AGEMA_signal_12562 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12565 ;
    wire new_AGEMA_signal_12566 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12569 ;
    wire new_AGEMA_signal_12570 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12573 ;
    wire new_AGEMA_signal_12574 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12577 ;
    wire new_AGEMA_signal_12578 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12581 ;
    wire new_AGEMA_signal_12582 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12585 ;
    wire new_AGEMA_signal_12586 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12589 ;
    wire new_AGEMA_signal_12590 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12593 ;
    wire new_AGEMA_signal_12594 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12597 ;
    wire new_AGEMA_signal_12598 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12601 ;
    wire new_AGEMA_signal_12602 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12605 ;
    wire new_AGEMA_signal_12606 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12609 ;
    wire new_AGEMA_signal_12610 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12613 ;
    wire new_AGEMA_signal_12614 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12617 ;
    wire new_AGEMA_signal_12618 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12621 ;
    wire new_AGEMA_signal_12622 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12625 ;
    wire new_AGEMA_signal_12626 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12629 ;
    wire new_AGEMA_signal_12630 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12633 ;
    wire new_AGEMA_signal_12634 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12637 ;
    wire new_AGEMA_signal_12638 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12641 ;
    wire new_AGEMA_signal_12642 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12645 ;
    wire new_AGEMA_signal_12646 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12649 ;
    wire new_AGEMA_signal_12650 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12653 ;
    wire new_AGEMA_signal_12654 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12657 ;
    wire new_AGEMA_signal_12658 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12661 ;
    wire new_AGEMA_signal_12662 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12665 ;
    wire new_AGEMA_signal_12666 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12669 ;
    wire new_AGEMA_signal_12670 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12673 ;
    wire new_AGEMA_signal_12674 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12677 ;
    wire new_AGEMA_signal_12678 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12681 ;
    wire new_AGEMA_signal_12682 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12685 ;
    wire new_AGEMA_signal_12686 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12689 ;
    wire new_AGEMA_signal_12690 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12693 ;
    wire new_AGEMA_signal_12694 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12697 ;
    wire new_AGEMA_signal_12698 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12701 ;
    wire new_AGEMA_signal_12702 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12705 ;
    wire new_AGEMA_signal_12706 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12709 ;
    wire new_AGEMA_signal_12710 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12713 ;
    wire new_AGEMA_signal_12714 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12717 ;
    wire new_AGEMA_signal_12718 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12721 ;
    wire new_AGEMA_signal_12722 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12725 ;
    wire new_AGEMA_signal_12726 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12729 ;
    wire new_AGEMA_signal_12730 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12733 ;
    wire new_AGEMA_signal_12734 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12737 ;
    wire new_AGEMA_signal_12738 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12741 ;
    wire new_AGEMA_signal_12742 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12745 ;
    wire new_AGEMA_signal_12746 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12749 ;
    wire new_AGEMA_signal_12750 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12753 ;
    wire new_AGEMA_signal_12754 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12757 ;
    wire new_AGEMA_signal_12758 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12761 ;
    wire new_AGEMA_signal_12762 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12765 ;
    wire new_AGEMA_signal_12766 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12769 ;
    wire new_AGEMA_signal_12770 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12773 ;
    wire new_AGEMA_signal_12774 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12777 ;
    wire new_AGEMA_signal_12778 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12781 ;
    wire new_AGEMA_signal_12782 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12785 ;
    wire new_AGEMA_signal_12786 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12789 ;
    wire new_AGEMA_signal_12790 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12793 ;
    wire new_AGEMA_signal_12794 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12797 ;
    wire new_AGEMA_signal_12798 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12801 ;
    wire new_AGEMA_signal_12802 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12805 ;
    wire new_AGEMA_signal_12806 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12809 ;
    wire new_AGEMA_signal_12810 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12813 ;
    wire new_AGEMA_signal_12814 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12817 ;
    wire new_AGEMA_signal_12818 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12821 ;
    wire new_AGEMA_signal_12822 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12825 ;
    wire new_AGEMA_signal_12826 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12829 ;
    wire new_AGEMA_signal_12830 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12833 ;
    wire new_AGEMA_signal_12834 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12837 ;
    wire new_AGEMA_signal_12838 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12841 ;
    wire new_AGEMA_signal_12842 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12845 ;
    wire new_AGEMA_signal_12846 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12849 ;
    wire new_AGEMA_signal_12850 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_12853 ;
    wire new_AGEMA_signal_12854 ;
    wire new_AGEMA_signal_12855 ;
    wire new_AGEMA_signal_12856 ;
    wire new_AGEMA_signal_12857 ;
    wire new_AGEMA_signal_12858 ;
    wire new_AGEMA_signal_12859 ;
    wire new_AGEMA_signal_12860 ;
    wire new_AGEMA_signal_12861 ;
    wire new_AGEMA_signal_12862 ;
    wire new_AGEMA_signal_12863 ;
    wire new_AGEMA_signal_12864 ;
    wire new_AGEMA_signal_12865 ;
    wire new_AGEMA_signal_12866 ;
    wire new_AGEMA_signal_12867 ;
    wire new_AGEMA_signal_12868 ;
    wire new_AGEMA_signal_12869 ;
    wire new_AGEMA_signal_12870 ;
    wire new_AGEMA_signal_12871 ;
    wire new_AGEMA_signal_12872 ;
    wire new_AGEMA_signal_12873 ;
    wire new_AGEMA_signal_12874 ;
    wire new_AGEMA_signal_12875 ;
    wire new_AGEMA_signal_12876 ;
    wire new_AGEMA_signal_12877 ;
    wire new_AGEMA_signal_12878 ;
    wire new_AGEMA_signal_12879 ;
    wire new_AGEMA_signal_12880 ;
    wire new_AGEMA_signal_12881 ;
    wire new_AGEMA_signal_12882 ;
    wire new_AGEMA_signal_12883 ;
    wire new_AGEMA_signal_12884 ;
    wire new_AGEMA_signal_12885 ;
    wire new_AGEMA_signal_12886 ;
    wire new_AGEMA_signal_12887 ;
    wire new_AGEMA_signal_12888 ;
    wire new_AGEMA_signal_12889 ;
    wire new_AGEMA_signal_12890 ;
    wire new_AGEMA_signal_12891 ;
    wire new_AGEMA_signal_12892 ;
    wire new_AGEMA_signal_12893 ;
    wire new_AGEMA_signal_12894 ;
    wire new_AGEMA_signal_12895 ;
    wire new_AGEMA_signal_12896 ;
    wire new_AGEMA_signal_12897 ;
    wire new_AGEMA_signal_12898 ;
    wire new_AGEMA_signal_12899 ;
    wire new_AGEMA_signal_12900 ;
    wire new_AGEMA_signal_12901 ;
    wire new_AGEMA_signal_12902 ;
    wire new_AGEMA_signal_12903 ;
    wire new_AGEMA_signal_12904 ;
    wire new_AGEMA_signal_12905 ;
    wire new_AGEMA_signal_12906 ;
    wire new_AGEMA_signal_12907 ;
    wire new_AGEMA_signal_12908 ;
    wire new_AGEMA_signal_12909 ;
    wire new_AGEMA_signal_12910 ;
    wire new_AGEMA_signal_12911 ;
    wire new_AGEMA_signal_12912 ;
    wire new_AGEMA_signal_12913 ;
    wire new_AGEMA_signal_12914 ;
    wire new_AGEMA_signal_12915 ;
    wire new_AGEMA_signal_12916 ;
    wire new_AGEMA_signal_12917 ;
    wire new_AGEMA_signal_12918 ;
    wire new_AGEMA_signal_12919 ;
    wire new_AGEMA_signal_12920 ;
    wire new_AGEMA_signal_12921 ;
    wire new_AGEMA_signal_12922 ;
    wire new_AGEMA_signal_12923 ;
    wire new_AGEMA_signal_12924 ;
    wire new_AGEMA_signal_12925 ;
    wire new_AGEMA_signal_12926 ;
    wire new_AGEMA_signal_12927 ;
    wire new_AGEMA_signal_12928 ;
    wire new_AGEMA_signal_12929 ;
    wire new_AGEMA_signal_12930 ;
    wire new_AGEMA_signal_12931 ;
    wire new_AGEMA_signal_12932 ;
    wire new_AGEMA_signal_12933 ;
    wire new_AGEMA_signal_12934 ;
    wire new_AGEMA_signal_12935 ;
    wire new_AGEMA_signal_12936 ;
    wire new_AGEMA_signal_12937 ;
    wire new_AGEMA_signal_12938 ;
    wire new_AGEMA_signal_12939 ;
    wire new_AGEMA_signal_12940 ;
    wire new_AGEMA_signal_12941 ;
    wire new_AGEMA_signal_12942 ;
    wire new_AGEMA_signal_12943 ;
    wire new_AGEMA_signal_12944 ;
    wire new_AGEMA_signal_12945 ;
    wire new_AGEMA_signal_12946 ;
    wire new_AGEMA_signal_12947 ;
    wire new_AGEMA_signal_12948 ;
    wire new_AGEMA_signal_12949 ;
    wire new_AGEMA_signal_12950 ;
    wire new_AGEMA_signal_12951 ;
    wire new_AGEMA_signal_12952 ;
    wire new_AGEMA_signal_12953 ;
    wire new_AGEMA_signal_12954 ;
    wire new_AGEMA_signal_12955 ;
    wire new_AGEMA_signal_12956 ;
    wire new_AGEMA_signal_12957 ;
    wire new_AGEMA_signal_12958 ;
    wire new_AGEMA_signal_12959 ;
    wire new_AGEMA_signal_12960 ;
    wire new_AGEMA_signal_12961 ;
    wire new_AGEMA_signal_12962 ;
    wire new_AGEMA_signal_12963 ;
    wire new_AGEMA_signal_12964 ;
    wire new_AGEMA_signal_12965 ;
    wire new_AGEMA_signal_12966 ;
    wire new_AGEMA_signal_12967 ;
    wire new_AGEMA_signal_12968 ;
    wire new_AGEMA_signal_12969 ;
    wire new_AGEMA_signal_12970 ;
    wire new_AGEMA_signal_12971 ;
    wire new_AGEMA_signal_12972 ;
    wire new_AGEMA_signal_12973 ;
    wire new_AGEMA_signal_12974 ;
    wire new_AGEMA_signal_12975 ;
    wire new_AGEMA_signal_12976 ;
    wire new_AGEMA_signal_12977 ;
    wire new_AGEMA_signal_12978 ;
    wire new_AGEMA_signal_12979 ;
    wire new_AGEMA_signal_12980 ;
    wire new_AGEMA_signal_12981 ;
    wire new_AGEMA_signal_12982 ;
    wire new_AGEMA_signal_12983 ;
    wire new_AGEMA_signal_12984 ;
    wire new_AGEMA_signal_12985 ;
    wire new_AGEMA_signal_12986 ;
    wire new_AGEMA_signal_12987 ;
    wire new_AGEMA_signal_12988 ;
    wire new_AGEMA_signal_12989 ;
    wire new_AGEMA_signal_12990 ;
    wire new_AGEMA_signal_12991 ;
    wire new_AGEMA_signal_12992 ;
    wire new_AGEMA_signal_12993 ;
    wire new_AGEMA_signal_12994 ;
    wire new_AGEMA_signal_12995 ;
    wire new_AGEMA_signal_12996 ;
    wire new_AGEMA_signal_12997 ;
    wire new_AGEMA_signal_12998 ;
    wire new_AGEMA_signal_12999 ;
    wire new_AGEMA_signal_13000 ;
    wire new_AGEMA_signal_13001 ;
    wire new_AGEMA_signal_13002 ;
    wire new_AGEMA_signal_13003 ;
    wire new_AGEMA_signal_13004 ;
    wire new_AGEMA_signal_13005 ;
    wire new_AGEMA_signal_13006 ;
    wire new_AGEMA_signal_13007 ;
    wire new_AGEMA_signal_13008 ;
    wire new_AGEMA_signal_13009 ;
    wire new_AGEMA_signal_13010 ;
    wire new_AGEMA_signal_13011 ;
    wire new_AGEMA_signal_13012 ;
    wire new_AGEMA_signal_13013 ;
    wire new_AGEMA_signal_13014 ;
    wire new_AGEMA_signal_13015 ;
    wire new_AGEMA_signal_13016 ;
    wire new_AGEMA_signal_13017 ;
    wire new_AGEMA_signal_13018 ;
    wire new_AGEMA_signal_13019 ;
    wire new_AGEMA_signal_13020 ;
    wire new_AGEMA_signal_13021 ;
    wire new_AGEMA_signal_13022 ;
    wire new_AGEMA_signal_13023 ;
    wire new_AGEMA_signal_13024 ;
    wire new_AGEMA_signal_13025 ;
    wire new_AGEMA_signal_13026 ;
    wire new_AGEMA_signal_13027 ;
    wire new_AGEMA_signal_13028 ;
    wire new_AGEMA_signal_13029 ;
    wire new_AGEMA_signal_13030 ;
    wire new_AGEMA_signal_13031 ;
    wire new_AGEMA_signal_13032 ;
    wire new_AGEMA_signal_13033 ;
    wire new_AGEMA_signal_13034 ;
    wire new_AGEMA_signal_13035 ;
    wire new_AGEMA_signal_13036 ;
    wire new_AGEMA_signal_13037 ;
    wire new_AGEMA_signal_13038 ;
    wire new_AGEMA_signal_13039 ;
    wire new_AGEMA_signal_13040 ;
    wire new_AGEMA_signal_13041 ;
    wire new_AGEMA_signal_13042 ;
    wire new_AGEMA_signal_13043 ;
    wire new_AGEMA_signal_13044 ;
    wire new_AGEMA_signal_13045 ;
    wire new_AGEMA_signal_13046 ;
    wire new_AGEMA_signal_13047 ;
    wire new_AGEMA_signal_13048 ;
    wire new_AGEMA_signal_13049 ;
    wire new_AGEMA_signal_13050 ;
    wire new_AGEMA_signal_13051 ;
    wire new_AGEMA_signal_13052 ;
    wire new_AGEMA_signal_13053 ;
    wire new_AGEMA_signal_13054 ;
    wire new_AGEMA_signal_13055 ;
    wire new_AGEMA_signal_13056 ;
    wire new_AGEMA_signal_13057 ;
    wire new_AGEMA_signal_13058 ;
    wire new_AGEMA_signal_13059 ;
    wire new_AGEMA_signal_13060 ;
    wire new_AGEMA_signal_13061 ;
    wire new_AGEMA_signal_13062 ;
    wire new_AGEMA_signal_13063 ;
    wire new_AGEMA_signal_13064 ;
    wire new_AGEMA_signal_13065 ;
    wire new_AGEMA_signal_13066 ;
    wire new_AGEMA_signal_13067 ;
    wire new_AGEMA_signal_13068 ;
    wire new_AGEMA_signal_13069 ;
    wire new_AGEMA_signal_13070 ;
    wire new_AGEMA_signal_13071 ;
    wire new_AGEMA_signal_13072 ;
    wire new_AGEMA_signal_13073 ;
    wire new_AGEMA_signal_13074 ;
    wire new_AGEMA_signal_13075 ;
    wire new_AGEMA_signal_13076 ;
    wire new_AGEMA_signal_13077 ;
    wire new_AGEMA_signal_13078 ;
    wire new_AGEMA_signal_13079 ;
    wire new_AGEMA_signal_13080 ;
    wire new_AGEMA_signal_13081 ;
    wire new_AGEMA_signal_13082 ;
    wire new_AGEMA_signal_13083 ;
    wire new_AGEMA_signal_13084 ;
    wire new_AGEMA_signal_13085 ;
    wire new_AGEMA_signal_13086 ;
    wire new_AGEMA_signal_13087 ;
    wire new_AGEMA_signal_13088 ;
    wire new_AGEMA_signal_13089 ;
    wire new_AGEMA_signal_13090 ;
    wire new_AGEMA_signal_13091 ;
    wire new_AGEMA_signal_13092 ;
    wire new_AGEMA_signal_13093 ;
    wire new_AGEMA_signal_13094 ;
    wire new_AGEMA_signal_13095 ;
    wire new_AGEMA_signal_13096 ;
    wire new_AGEMA_signal_13097 ;
    wire new_AGEMA_signal_13098 ;
    wire new_AGEMA_signal_13099 ;
    wire new_AGEMA_signal_13100 ;
    wire new_AGEMA_signal_13101 ;
    wire new_AGEMA_signal_13102 ;
    wire new_AGEMA_signal_13103 ;
    wire new_AGEMA_signal_13104 ;
    wire new_AGEMA_signal_13105 ;
    wire new_AGEMA_signal_13106 ;
    wire new_AGEMA_signal_13107 ;
    wire new_AGEMA_signal_13108 ;
    wire new_AGEMA_signal_13109 ;
    wire new_AGEMA_signal_13110 ;
    wire new_AGEMA_signal_13111 ;
    wire new_AGEMA_signal_13112 ;
    wire new_AGEMA_signal_13113 ;
    wire new_AGEMA_signal_13114 ;
    wire new_AGEMA_signal_13115 ;
    wire new_AGEMA_signal_13116 ;
    wire new_AGEMA_signal_13117 ;
    wire new_AGEMA_signal_13118 ;
    wire new_AGEMA_signal_13119 ;
    wire new_AGEMA_signal_13120 ;
    wire new_AGEMA_signal_13121 ;
    wire new_AGEMA_signal_13122 ;
    wire new_AGEMA_signal_13123 ;
    wire new_AGEMA_signal_13124 ;
    wire new_AGEMA_signal_13125 ;
    wire new_AGEMA_signal_13126 ;
    wire new_AGEMA_signal_13127 ;
    wire new_AGEMA_signal_13128 ;
    wire new_AGEMA_signal_13129 ;
    wire new_AGEMA_signal_13130 ;
    wire new_AGEMA_signal_13131 ;
    wire new_AGEMA_signal_13132 ;
    wire new_AGEMA_signal_13133 ;
    wire new_AGEMA_signal_13134 ;
    wire new_AGEMA_signal_13135 ;
    wire new_AGEMA_signal_13136 ;
    wire new_AGEMA_signal_13137 ;
    wire new_AGEMA_signal_13138 ;
    wire new_AGEMA_signal_13139 ;
    wire new_AGEMA_signal_13140 ;
    wire new_AGEMA_signal_13141 ;
    wire new_AGEMA_signal_13142 ;
    wire new_AGEMA_signal_13143 ;
    wire new_AGEMA_signal_13144 ;
    wire new_AGEMA_signal_13145 ;
    wire new_AGEMA_signal_13146 ;
    wire new_AGEMA_signal_13147 ;
    wire new_AGEMA_signal_13148 ;
    wire new_AGEMA_signal_13149 ;
    wire new_AGEMA_signal_13150 ;
    wire new_AGEMA_signal_13151 ;
    wire new_AGEMA_signal_13152 ;
    wire new_AGEMA_signal_13153 ;
    wire new_AGEMA_signal_13154 ;
    wire new_AGEMA_signal_13155 ;
    wire new_AGEMA_signal_13156 ;
    wire new_AGEMA_signal_13157 ;
    wire new_AGEMA_signal_13158 ;
    wire new_AGEMA_signal_13159 ;
    wire new_AGEMA_signal_13160 ;
    wire new_AGEMA_signal_13161 ;
    wire new_AGEMA_signal_13162 ;
    wire new_AGEMA_signal_13163 ;
    wire new_AGEMA_signal_13164 ;
    wire new_AGEMA_signal_13165 ;
    wire new_AGEMA_signal_13166 ;
    wire new_AGEMA_signal_13167 ;
    wire new_AGEMA_signal_13168 ;
    wire new_AGEMA_signal_13169 ;
    wire new_AGEMA_signal_13170 ;
    wire new_AGEMA_signal_13171 ;
    wire new_AGEMA_signal_13172 ;
    wire new_AGEMA_signal_13173 ;
    wire new_AGEMA_signal_13174 ;
    wire new_AGEMA_signal_13175 ;
    wire new_AGEMA_signal_13176 ;
    wire new_AGEMA_signal_13177 ;
    wire new_AGEMA_signal_13178 ;
    wire new_AGEMA_signal_13179 ;
    wire new_AGEMA_signal_13180 ;
    wire new_AGEMA_signal_13181 ;
    wire new_AGEMA_signal_13182 ;
    wire new_AGEMA_signal_13183 ;
    wire new_AGEMA_signal_13184 ;
    wire new_AGEMA_signal_13185 ;
    wire new_AGEMA_signal_13186 ;
    wire new_AGEMA_signal_13187 ;
    wire new_AGEMA_signal_13188 ;
    wire new_AGEMA_signal_13189 ;
    wire new_AGEMA_signal_13190 ;
    wire new_AGEMA_signal_13191 ;
    wire new_AGEMA_signal_13192 ;
    wire new_AGEMA_signal_13193 ;
    wire new_AGEMA_signal_13194 ;
    wire new_AGEMA_signal_13195 ;
    wire new_AGEMA_signal_13196 ;
    wire new_AGEMA_signal_13197 ;
    wire new_AGEMA_signal_13198 ;
    wire new_AGEMA_signal_13199 ;
    wire new_AGEMA_signal_13200 ;
    wire new_AGEMA_signal_13201 ;
    wire new_AGEMA_signal_13202 ;
    wire new_AGEMA_signal_13203 ;
    wire new_AGEMA_signal_13204 ;
    wire new_AGEMA_signal_13205 ;
    wire new_AGEMA_signal_13206 ;
    wire new_AGEMA_signal_13207 ;
    wire new_AGEMA_signal_13208 ;
    wire new_AGEMA_signal_13209 ;
    wire new_AGEMA_signal_13210 ;
    wire new_AGEMA_signal_13211 ;
    wire new_AGEMA_signal_13212 ;
    wire new_AGEMA_signal_13213 ;
    wire new_AGEMA_signal_13214 ;
    wire new_AGEMA_signal_13215 ;
    wire new_AGEMA_signal_13216 ;
    wire new_AGEMA_signal_13217 ;
    wire new_AGEMA_signal_13218 ;
    wire new_AGEMA_signal_13219 ;
    wire new_AGEMA_signal_13220 ;
    wire new_AGEMA_signal_13221 ;
    wire new_AGEMA_signal_13222 ;
    wire new_AGEMA_signal_13223 ;
    wire new_AGEMA_signal_13224 ;
    wire new_AGEMA_signal_13225 ;
    wire new_AGEMA_signal_13226 ;
    wire new_AGEMA_signal_13227 ;
    wire new_AGEMA_signal_13228 ;
    wire new_AGEMA_signal_13229 ;
    wire new_AGEMA_signal_13230 ;
    wire new_AGEMA_signal_13231 ;
    wire new_AGEMA_signal_13232 ;
    wire new_AGEMA_signal_13233 ;
    wire new_AGEMA_signal_13234 ;
    wire new_AGEMA_signal_13235 ;
    wire new_AGEMA_signal_13236 ;
    wire new_AGEMA_signal_13237 ;
    wire new_AGEMA_signal_13238 ;
    wire new_AGEMA_signal_13239 ;
    wire new_AGEMA_signal_13240 ;
    wire new_AGEMA_signal_13241 ;
    wire new_AGEMA_signal_13242 ;
    wire new_AGEMA_signal_13243 ;
    wire new_AGEMA_signal_13244 ;
    wire new_AGEMA_signal_13245 ;
    wire new_AGEMA_signal_13246 ;
    wire new_AGEMA_signal_13247 ;
    wire new_AGEMA_signal_13248 ;
    wire new_AGEMA_signal_13249 ;
    wire new_AGEMA_signal_13250 ;
    wire new_AGEMA_signal_13251 ;
    wire new_AGEMA_signal_13252 ;
    wire new_AGEMA_signal_13253 ;
    wire new_AGEMA_signal_13254 ;
    wire new_AGEMA_signal_13255 ;
    wire new_AGEMA_signal_13256 ;
    wire new_AGEMA_signal_13257 ;
    wire new_AGEMA_signal_13258 ;
    wire new_AGEMA_signal_13259 ;
    wire new_AGEMA_signal_13260 ;
    wire new_AGEMA_signal_13261 ;
    wire new_AGEMA_signal_13262 ;
    wire new_AGEMA_signal_13263 ;
    wire new_AGEMA_signal_13264 ;
    wire new_AGEMA_signal_13265 ;
    wire new_AGEMA_signal_13266 ;
    wire new_AGEMA_signal_13267 ;
    wire new_AGEMA_signal_13268 ;
    wire new_AGEMA_signal_13269 ;
    wire new_AGEMA_signal_13270 ;
    wire new_AGEMA_signal_13271 ;
    wire new_AGEMA_signal_13272 ;
    wire new_AGEMA_signal_13273 ;
    wire new_AGEMA_signal_13274 ;
    wire new_AGEMA_signal_13275 ;
    wire new_AGEMA_signal_13276 ;
    wire new_AGEMA_signal_13277 ;
    wire new_AGEMA_signal_13278 ;
    wire new_AGEMA_signal_13279 ;
    wire new_AGEMA_signal_13280 ;
    wire new_AGEMA_signal_13281 ;
    wire new_AGEMA_signal_13282 ;
    wire new_AGEMA_signal_13283 ;
    wire new_AGEMA_signal_13284 ;
    wire new_AGEMA_signal_13285 ;
    wire new_AGEMA_signal_13286 ;
    wire new_AGEMA_signal_13287 ;
    wire new_AGEMA_signal_13288 ;
    wire new_AGEMA_signal_13289 ;
    wire new_AGEMA_signal_13290 ;
    wire new_AGEMA_signal_13291 ;
    wire new_AGEMA_signal_13292 ;
    wire new_AGEMA_signal_13293 ;
    wire new_AGEMA_signal_13294 ;
    wire new_AGEMA_signal_13295 ;
    wire new_AGEMA_signal_13296 ;
    wire new_AGEMA_signal_13297 ;
    wire new_AGEMA_signal_13298 ;
    wire new_AGEMA_signal_13299 ;
    wire new_AGEMA_signal_13300 ;
    wire new_AGEMA_signal_13301 ;
    wire new_AGEMA_signal_13302 ;
    wire new_AGEMA_signal_13303 ;
    wire new_AGEMA_signal_13304 ;
    wire new_AGEMA_signal_13305 ;
    wire new_AGEMA_signal_13306 ;
    wire new_AGEMA_signal_13307 ;
    wire new_AGEMA_signal_13308 ;
    wire new_AGEMA_signal_13309 ;
    wire new_AGEMA_signal_13310 ;
    wire new_AGEMA_signal_13311 ;
    wire new_AGEMA_signal_13312 ;
    wire new_AGEMA_signal_13313 ;
    wire new_AGEMA_signal_13314 ;
    wire new_AGEMA_signal_13315 ;
    wire new_AGEMA_signal_13316 ;
    wire new_AGEMA_signal_13317 ;
    wire new_AGEMA_signal_13318 ;
    wire new_AGEMA_signal_13319 ;
    wire new_AGEMA_signal_13320 ;
    wire new_AGEMA_signal_13321 ;
    wire new_AGEMA_signal_13322 ;
    wire new_AGEMA_signal_13323 ;
    wire new_AGEMA_signal_13324 ;
    wire new_AGEMA_signal_13325 ;
    wire new_AGEMA_signal_13326 ;
    wire new_AGEMA_signal_13327 ;
    wire new_AGEMA_signal_13328 ;
    wire new_AGEMA_signal_13329 ;
    wire new_AGEMA_signal_13330 ;
    wire new_AGEMA_signal_13331 ;
    wire new_AGEMA_signal_13332 ;
    wire new_AGEMA_signal_13333 ;
    wire new_AGEMA_signal_13334 ;
    wire new_AGEMA_signal_13335 ;
    wire new_AGEMA_signal_13336 ;
    wire new_AGEMA_signal_13337 ;
    wire new_AGEMA_signal_13338 ;
    wire new_AGEMA_signal_13339 ;
    wire new_AGEMA_signal_13340 ;
    wire new_AGEMA_signal_13341 ;
    wire new_AGEMA_signal_13342 ;
    wire new_AGEMA_signal_13343 ;
    wire new_AGEMA_signal_13344 ;
    wire new_AGEMA_signal_13345 ;
    wire new_AGEMA_signal_13346 ;
    wire new_AGEMA_signal_13347 ;
    wire new_AGEMA_signal_13348 ;
    wire new_AGEMA_signal_13349 ;
    wire new_AGEMA_signal_13350 ;
    wire new_AGEMA_signal_13351 ;
    wire new_AGEMA_signal_13352 ;
    wire new_AGEMA_signal_13353 ;
    wire new_AGEMA_signal_13354 ;
    wire new_AGEMA_signal_13355 ;
    wire new_AGEMA_signal_13356 ;
    wire new_AGEMA_signal_13357 ;
    wire new_AGEMA_signal_13358 ;
    wire new_AGEMA_signal_13359 ;
    wire new_AGEMA_signal_13360 ;
    wire new_AGEMA_signal_13361 ;
    wire new_AGEMA_signal_13362 ;
    wire new_AGEMA_signal_13363 ;
    wire new_AGEMA_signal_13364 ;
    wire new_AGEMA_signal_13365 ;
    wire new_AGEMA_signal_13366 ;
    wire new_AGEMA_signal_13367 ;
    wire new_AGEMA_signal_13368 ;
    wire new_AGEMA_signal_13369 ;
    wire new_AGEMA_signal_13370 ;
    wire new_AGEMA_signal_13371 ;
    wire new_AGEMA_signal_13372 ;
    wire new_AGEMA_signal_13373 ;
    wire new_AGEMA_signal_13374 ;
    wire new_AGEMA_signal_13375 ;
    wire new_AGEMA_signal_13376 ;
    wire new_AGEMA_signal_13377 ;
    wire new_AGEMA_signal_13378 ;
    wire new_AGEMA_signal_13379 ;
    wire new_AGEMA_signal_13380 ;
    wire new_AGEMA_signal_13381 ;
    wire new_AGEMA_signal_13382 ;
    wire new_AGEMA_signal_13383 ;
    wire new_AGEMA_signal_13384 ;
    wire new_AGEMA_signal_13385 ;
    wire new_AGEMA_signal_13386 ;
    wire new_AGEMA_signal_13387 ;
    wire new_AGEMA_signal_13388 ;
    wire new_AGEMA_signal_13389 ;
    wire new_AGEMA_signal_13390 ;
    wire new_AGEMA_signal_13391 ;
    wire new_AGEMA_signal_13392 ;
    wire new_AGEMA_signal_13393 ;
    wire new_AGEMA_signal_13394 ;
    wire new_AGEMA_signal_13395 ;
    wire new_AGEMA_signal_13396 ;
    wire new_AGEMA_signal_13397 ;
    wire new_AGEMA_signal_13398 ;
    wire new_AGEMA_signal_13399 ;
    wire new_AGEMA_signal_13400 ;
    wire new_AGEMA_signal_13401 ;
    wire new_AGEMA_signal_13402 ;
    wire new_AGEMA_signal_13403 ;
    wire new_AGEMA_signal_13404 ;
    wire new_AGEMA_signal_13405 ;
    wire new_AGEMA_signal_13406 ;
    wire new_AGEMA_signal_13407 ;
    wire new_AGEMA_signal_13408 ;
    wire new_AGEMA_signal_13409 ;
    wire new_AGEMA_signal_13410 ;
    wire new_AGEMA_signal_13411 ;
    wire new_AGEMA_signal_13412 ;
    wire new_AGEMA_signal_13413 ;
    wire new_AGEMA_signal_13414 ;
    wire new_AGEMA_signal_13415 ;
    wire new_AGEMA_signal_13416 ;
    wire new_AGEMA_signal_13417 ;
    wire new_AGEMA_signal_13418 ;
    wire new_AGEMA_signal_13419 ;
    wire new_AGEMA_signal_13420 ;
    wire new_AGEMA_signal_13421 ;
    wire new_AGEMA_signal_13422 ;
    wire new_AGEMA_signal_13423 ;
    wire new_AGEMA_signal_13424 ;
    wire new_AGEMA_signal_13425 ;
    wire new_AGEMA_signal_13426 ;
    wire new_AGEMA_signal_13427 ;
    wire new_AGEMA_signal_13428 ;
    wire new_AGEMA_signal_13429 ;
    wire new_AGEMA_signal_13430 ;
    wire new_AGEMA_signal_13431 ;
    wire new_AGEMA_signal_13432 ;
    wire new_AGEMA_signal_13433 ;
    wire new_AGEMA_signal_13434 ;
    wire new_AGEMA_signal_13435 ;
    wire new_AGEMA_signal_13436 ;
    wire new_AGEMA_signal_13437 ;
    wire new_AGEMA_signal_13438 ;
    wire new_AGEMA_signal_13439 ;
    wire new_AGEMA_signal_13440 ;
    wire new_AGEMA_signal_13441 ;
    wire new_AGEMA_signal_13442 ;
    wire new_AGEMA_signal_13443 ;
    wire new_AGEMA_signal_13444 ;
    wire new_AGEMA_signal_13445 ;
    wire new_AGEMA_signal_13446 ;
    wire new_AGEMA_signal_13447 ;
    wire new_AGEMA_signal_13448 ;
    wire new_AGEMA_signal_13449 ;
    wire new_AGEMA_signal_13450 ;
    wire new_AGEMA_signal_13451 ;
    wire new_AGEMA_signal_13452 ;
    wire new_AGEMA_signal_13453 ;
    wire new_AGEMA_signal_13454 ;
    wire new_AGEMA_signal_13455 ;
    wire new_AGEMA_signal_13456 ;
    wire new_AGEMA_signal_13457 ;
    wire new_AGEMA_signal_13458 ;
    wire new_AGEMA_signal_13459 ;
    wire new_AGEMA_signal_13460 ;
    wire new_AGEMA_signal_13461 ;
    wire new_AGEMA_signal_13462 ;
    wire new_AGEMA_signal_13463 ;
    wire new_AGEMA_signal_13464 ;
    wire new_AGEMA_signal_13465 ;
    wire new_AGEMA_signal_13466 ;
    wire new_AGEMA_signal_13467 ;
    wire new_AGEMA_signal_13468 ;
    wire new_AGEMA_signal_13469 ;
    wire new_AGEMA_signal_13470 ;
    wire new_AGEMA_signal_13471 ;
    wire new_AGEMA_signal_13472 ;
    wire new_AGEMA_signal_13473 ;
    wire new_AGEMA_signal_13474 ;
    wire new_AGEMA_signal_13475 ;
    wire new_AGEMA_signal_13476 ;
    wire new_AGEMA_signal_13477 ;
    wire new_AGEMA_signal_13478 ;
    wire new_AGEMA_signal_13479 ;
    wire new_AGEMA_signal_13480 ;
    wire new_AGEMA_signal_13481 ;
    wire new_AGEMA_signal_13482 ;
    wire new_AGEMA_signal_13483 ;
    wire new_AGEMA_signal_13484 ;
    wire new_AGEMA_signal_13485 ;
    wire new_AGEMA_signal_13486 ;
    wire new_AGEMA_signal_13487 ;
    wire new_AGEMA_signal_13488 ;
    wire new_AGEMA_signal_13489 ;
    wire new_AGEMA_signal_13490 ;
    wire new_AGEMA_signal_13491 ;
    wire new_AGEMA_signal_13492 ;
    wire new_AGEMA_signal_13493 ;
    wire new_AGEMA_signal_13494 ;
    wire new_AGEMA_signal_13495 ;
    wire new_AGEMA_signal_13496 ;
    wire new_AGEMA_signal_13497 ;
    wire new_AGEMA_signal_13498 ;
    wire new_AGEMA_signal_13499 ;
    wire new_AGEMA_signal_13500 ;
    wire new_AGEMA_signal_13501 ;
    wire new_AGEMA_signal_13502 ;
    wire new_AGEMA_signal_13503 ;
    wire new_AGEMA_signal_13504 ;
    wire new_AGEMA_signal_13505 ;
    wire new_AGEMA_signal_13506 ;
    wire new_AGEMA_signal_13507 ;
    wire new_AGEMA_signal_13508 ;
    wire new_AGEMA_signal_13509 ;
    wire new_AGEMA_signal_13510 ;
    wire new_AGEMA_signal_13511 ;
    wire new_AGEMA_signal_13512 ;
    wire new_AGEMA_signal_13513 ;
    wire new_AGEMA_signal_13514 ;
    wire new_AGEMA_signal_13515 ;
    wire new_AGEMA_signal_13516 ;
    wire new_AGEMA_signal_13517 ;
    wire new_AGEMA_signal_13518 ;
    wire new_AGEMA_signal_13519 ;
    wire new_AGEMA_signal_13520 ;
    wire new_AGEMA_signal_13521 ;
    wire new_AGEMA_signal_13522 ;
    wire new_AGEMA_signal_13523 ;
    wire new_AGEMA_signal_13524 ;
    wire new_AGEMA_signal_13525 ;
    wire new_AGEMA_signal_13526 ;
    wire new_AGEMA_signal_13527 ;
    wire new_AGEMA_signal_13528 ;
    wire new_AGEMA_signal_13529 ;
    wire new_AGEMA_signal_13530 ;
    wire new_AGEMA_signal_13531 ;
    wire new_AGEMA_signal_13532 ;
    wire new_AGEMA_signal_13533 ;
    wire new_AGEMA_signal_13534 ;
    wire new_AGEMA_signal_13535 ;
    wire new_AGEMA_signal_13536 ;
    wire new_AGEMA_signal_13537 ;
    wire new_AGEMA_signal_13538 ;
    wire new_AGEMA_signal_13539 ;
    wire new_AGEMA_signal_13540 ;
    wire new_AGEMA_signal_13541 ;
    wire new_AGEMA_signal_13542 ;
    wire new_AGEMA_signal_13543 ;
    wire new_AGEMA_signal_13544 ;
    wire new_AGEMA_signal_13545 ;
    wire new_AGEMA_signal_13546 ;
    wire new_AGEMA_signal_13547 ;
    wire new_AGEMA_signal_13548 ;
    wire new_AGEMA_signal_13549 ;
    wire new_AGEMA_signal_13550 ;
    wire new_AGEMA_signal_13551 ;
    wire new_AGEMA_signal_13552 ;
    wire new_AGEMA_signal_13553 ;
    wire new_AGEMA_signal_13554 ;
    wire new_AGEMA_signal_13555 ;
    wire new_AGEMA_signal_13558 ;
    wire new_AGEMA_signal_13559 ;
    wire new_AGEMA_signal_13560 ;
    wire new_AGEMA_signal_13561 ;
    wire new_AGEMA_signal_13566 ;
    wire new_AGEMA_signal_13567 ;
    wire new_AGEMA_signal_13568 ;
    wire new_AGEMA_signal_13569 ;
    wire new_AGEMA_signal_13570 ;
    wire new_AGEMA_signal_13571 ;
    wire new_AGEMA_signal_13572 ;
    wire new_AGEMA_signal_13573 ;
    wire new_AGEMA_signal_13574 ;
    wire new_AGEMA_signal_13575 ;
    wire new_AGEMA_signal_13576 ;
    wire new_AGEMA_signal_13577 ;
    wire new_AGEMA_signal_13578 ;
    wire new_AGEMA_signal_13579 ;
    wire new_AGEMA_signal_13580 ;
    wire new_AGEMA_signal_13581 ;
    wire new_AGEMA_signal_13582 ;
    wire new_AGEMA_signal_13583 ;
    wire new_AGEMA_signal_13584 ;
    wire new_AGEMA_signal_13585 ;
    wire new_AGEMA_signal_13586 ;
    wire new_AGEMA_signal_13587 ;
    wire new_AGEMA_signal_13588 ;
    wire new_AGEMA_signal_13589 ;
    wire new_AGEMA_signal_13590 ;
    wire new_AGEMA_signal_13591 ;
    wire new_AGEMA_signal_13592 ;
    wire new_AGEMA_signal_13593 ;
    wire new_AGEMA_signal_13594 ;
    wire new_AGEMA_signal_13595 ;
    wire new_AGEMA_signal_13596 ;
    wire new_AGEMA_signal_13597 ;
    wire new_AGEMA_signal_13598 ;
    wire new_AGEMA_signal_13599 ;
    wire new_AGEMA_signal_13600 ;
    wire new_AGEMA_signal_13601 ;
    wire new_AGEMA_signal_13602 ;
    wire new_AGEMA_signal_13603 ;
    wire new_AGEMA_signal_13604 ;
    wire new_AGEMA_signal_13605 ;
    wire new_AGEMA_signal_13606 ;
    wire new_AGEMA_signal_13607 ;
    wire new_AGEMA_signal_13608 ;
    wire new_AGEMA_signal_13609 ;
    wire new_AGEMA_signal_13610 ;
    wire new_AGEMA_signal_13611 ;
    wire new_AGEMA_signal_13612 ;
    wire new_AGEMA_signal_13613 ;
    wire new_AGEMA_signal_13614 ;
    wire new_AGEMA_signal_13615 ;
    wire new_AGEMA_signal_13616 ;
    wire new_AGEMA_signal_13617 ;
    wire new_AGEMA_signal_13618 ;
    wire new_AGEMA_signal_13619 ;
    wire new_AGEMA_signal_13620 ;
    wire new_AGEMA_signal_13621 ;
    wire new_AGEMA_signal_13622 ;
    wire new_AGEMA_signal_13623 ;
    wire new_AGEMA_signal_13624 ;
    wire new_AGEMA_signal_13625 ;
    wire new_AGEMA_signal_13626 ;
    wire new_AGEMA_signal_13627 ;
    wire new_AGEMA_signal_13628 ;
    wire new_AGEMA_signal_13629 ;
    wire new_AGEMA_signal_13630 ;
    wire new_AGEMA_signal_13631 ;
    wire new_AGEMA_signal_13632 ;
    wire new_AGEMA_signal_13633 ;
    wire new_AGEMA_signal_13634 ;
    wire new_AGEMA_signal_13635 ;
    wire new_AGEMA_signal_13636 ;
    wire new_AGEMA_signal_13637 ;
    wire new_AGEMA_signal_13638 ;
    wire new_AGEMA_signal_13639 ;
    wire new_AGEMA_signal_13640 ;
    wire new_AGEMA_signal_13641 ;
    wire new_AGEMA_signal_13642 ;
    wire new_AGEMA_signal_13643 ;
    wire new_AGEMA_signal_13644 ;
    wire new_AGEMA_signal_13645 ;
    wire new_AGEMA_signal_13646 ;
    wire new_AGEMA_signal_13647 ;
    wire new_AGEMA_signal_13648 ;
    wire new_AGEMA_signal_13649 ;
    wire new_AGEMA_signal_13650 ;
    wire new_AGEMA_signal_13651 ;
    wire new_AGEMA_signal_13652 ;
    wire new_AGEMA_signal_13653 ;
    wire new_AGEMA_signal_13654 ;
    wire new_AGEMA_signal_13655 ;
    wire new_AGEMA_signal_13656 ;
    wire new_AGEMA_signal_13657 ;
    wire new_AGEMA_signal_13658 ;
    wire new_AGEMA_signal_13659 ;
    wire new_AGEMA_signal_13660 ;
    wire new_AGEMA_signal_13661 ;
    wire new_AGEMA_signal_13662 ;
    wire new_AGEMA_signal_13663 ;
    wire new_AGEMA_signal_13664 ;
    wire new_AGEMA_signal_13665 ;
    wire new_AGEMA_signal_13666 ;
    wire new_AGEMA_signal_13667 ;
    wire new_AGEMA_signal_13668 ;
    wire new_AGEMA_signal_13669 ;
    wire new_AGEMA_signal_13670 ;
    wire new_AGEMA_signal_13671 ;
    wire new_AGEMA_signal_13672 ;
    wire new_AGEMA_signal_13673 ;
    wire new_AGEMA_signal_13674 ;
    wire new_AGEMA_signal_13675 ;
    wire new_AGEMA_signal_13676 ;
    wire new_AGEMA_signal_13677 ;
    wire new_AGEMA_signal_13678 ;
    wire new_AGEMA_signal_13679 ;
    wire new_AGEMA_signal_13680 ;
    wire new_AGEMA_signal_13681 ;
    wire new_AGEMA_signal_13682 ;
    wire new_AGEMA_signal_13683 ;
    wire new_AGEMA_signal_13684 ;
    wire new_AGEMA_signal_13685 ;
    wire new_AGEMA_signal_13686 ;
    wire new_AGEMA_signal_13687 ;
    wire new_AGEMA_signal_13688 ;
    wire new_AGEMA_signal_13689 ;
    wire new_AGEMA_signal_13690 ;
    wire new_AGEMA_signal_13691 ;
    wire new_AGEMA_signal_13692 ;
    wire new_AGEMA_signal_13693 ;
    wire new_AGEMA_signal_13694 ;
    wire new_AGEMA_signal_13695 ;
    wire new_AGEMA_signal_13696 ;
    wire new_AGEMA_signal_13697 ;
    wire new_AGEMA_signal_13698 ;
    wire new_AGEMA_signal_13699 ;
    wire new_AGEMA_signal_13700 ;
    wire new_AGEMA_signal_13701 ;
    wire new_AGEMA_signal_13702 ;
    wire new_AGEMA_signal_13703 ;
    wire new_AGEMA_signal_13704 ;
    wire new_AGEMA_signal_13705 ;
    wire new_AGEMA_signal_13706 ;
    wire new_AGEMA_signal_13707 ;
    wire new_AGEMA_signal_13708 ;
    wire new_AGEMA_signal_13709 ;
    wire new_AGEMA_signal_13710 ;
    wire new_AGEMA_signal_13711 ;
    wire new_AGEMA_signal_13712 ;
    wire new_AGEMA_signal_13713 ;
    wire new_AGEMA_signal_13714 ;
    wire new_AGEMA_signal_13715 ;
    wire new_AGEMA_signal_13716 ;
    wire new_AGEMA_signal_13717 ;
    wire new_AGEMA_signal_13718 ;
    wire new_AGEMA_signal_13719 ;
    wire new_AGEMA_signal_13720 ;
    wire new_AGEMA_signal_13721 ;
    wire new_AGEMA_signal_13722 ;
    wire new_AGEMA_signal_13723 ;
    wire new_AGEMA_signal_13724 ;
    wire new_AGEMA_signal_13725 ;
    wire new_AGEMA_signal_13726 ;
    wire new_AGEMA_signal_13727 ;
    wire new_AGEMA_signal_13728 ;
    wire new_AGEMA_signal_13729 ;
    wire new_AGEMA_signal_13730 ;
    wire new_AGEMA_signal_13731 ;
    wire new_AGEMA_signal_13732 ;
    wire new_AGEMA_signal_13733 ;
    wire new_AGEMA_signal_13734 ;
    wire new_AGEMA_signal_13735 ;
    wire new_AGEMA_signal_13736 ;
    wire new_AGEMA_signal_13737 ;
    wire new_AGEMA_signal_13738 ;
    wire new_AGEMA_signal_13739 ;
    wire new_AGEMA_signal_13740 ;
    wire new_AGEMA_signal_13741 ;
    wire new_AGEMA_signal_13742 ;
    wire new_AGEMA_signal_13743 ;
    wire new_AGEMA_signal_13744 ;
    wire new_AGEMA_signal_13745 ;
    wire new_AGEMA_signal_13746 ;
    wire new_AGEMA_signal_13747 ;
    wire new_AGEMA_signal_13748 ;
    wire new_AGEMA_signal_13749 ;
    wire new_AGEMA_signal_13750 ;
    wire new_AGEMA_signal_13751 ;
    wire new_AGEMA_signal_13752 ;
    wire new_AGEMA_signal_13753 ;
    wire new_AGEMA_signal_13754 ;
    wire new_AGEMA_signal_13755 ;
    wire new_AGEMA_signal_13756 ;
    wire new_AGEMA_signal_13757 ;
    wire new_AGEMA_signal_13758 ;
    wire new_AGEMA_signal_13759 ;
    wire new_AGEMA_signal_13760 ;
    wire new_AGEMA_signal_13761 ;
    wire new_AGEMA_signal_13762 ;
    wire new_AGEMA_signal_13763 ;
    wire new_AGEMA_signal_13764 ;
    wire new_AGEMA_signal_13765 ;
    wire new_AGEMA_signal_13766 ;
    wire new_AGEMA_signal_13767 ;
    wire new_AGEMA_signal_13768 ;
    wire new_AGEMA_signal_13769 ;
    wire new_AGEMA_signal_13770 ;
    wire new_AGEMA_signal_13771 ;
    wire new_AGEMA_signal_13772 ;
    wire new_AGEMA_signal_13773 ;
    wire new_AGEMA_signal_13776 ;
    wire new_AGEMA_signal_13777 ;
    wire new_AGEMA_signal_13778 ;
    wire new_AGEMA_signal_13779 ;
    wire new_AGEMA_signal_13784 ;
    wire new_AGEMA_signal_13785 ;
    wire new_AGEMA_signal_13786 ;
    wire new_AGEMA_signal_13787 ;
    wire new_AGEMA_signal_13788 ;
    wire new_AGEMA_signal_13789 ;
    wire new_AGEMA_signal_13790 ;
    wire new_AGEMA_signal_13791 ;
    wire new_AGEMA_signal_13792 ;
    wire new_AGEMA_signal_13793 ;
    wire new_AGEMA_signal_13794 ;
    wire new_AGEMA_signal_13795 ;
    wire new_AGEMA_signal_13796 ;
    wire new_AGEMA_signal_13797 ;
    wire new_AGEMA_signal_13798 ;
    wire new_AGEMA_signal_13799 ;
    wire new_AGEMA_signal_13800 ;
    wire new_AGEMA_signal_13801 ;
    wire new_AGEMA_signal_13802 ;
    wire new_AGEMA_signal_13803 ;
    wire new_AGEMA_signal_13804 ;
    wire new_AGEMA_signal_13805 ;
    wire new_AGEMA_signal_13806 ;
    wire new_AGEMA_signal_13807 ;
    wire new_AGEMA_signal_13808 ;
    wire new_AGEMA_signal_13809 ;
    wire new_AGEMA_signal_13810 ;
    wire new_AGEMA_signal_13811 ;
    wire new_AGEMA_signal_13812 ;
    wire new_AGEMA_signal_13813 ;
    wire new_AGEMA_signal_13814 ;
    wire new_AGEMA_signal_13815 ;
    wire new_AGEMA_signal_13816 ;
    wire new_AGEMA_signal_13817 ;
    wire new_AGEMA_signal_13818 ;
    wire new_AGEMA_signal_13819 ;
    wire new_AGEMA_signal_13820 ;
    wire new_AGEMA_signal_13821 ;
    wire new_AGEMA_signal_13822 ;
    wire new_AGEMA_signal_13823 ;
    wire new_AGEMA_signal_13824 ;
    wire new_AGEMA_signal_13825 ;
    wire new_AGEMA_signal_13826 ;
    wire new_AGEMA_signal_13827 ;
    wire new_AGEMA_signal_13828 ;
    wire new_AGEMA_signal_13829 ;
    wire new_AGEMA_signal_13830 ;
    wire new_AGEMA_signal_13831 ;
    wire new_AGEMA_signal_13832 ;
    wire new_AGEMA_signal_13833 ;
    wire new_AGEMA_signal_13834 ;
    wire new_AGEMA_signal_13835 ;
    wire new_AGEMA_signal_13836 ;
    wire new_AGEMA_signal_13837 ;
    wire new_AGEMA_signal_13838 ;
    wire new_AGEMA_signal_13839 ;
    wire new_AGEMA_signal_13840 ;
    wire new_AGEMA_signal_13841 ;
    wire new_AGEMA_signal_13842 ;
    wire new_AGEMA_signal_13843 ;
    wire new_AGEMA_signal_13844 ;
    wire new_AGEMA_signal_13845 ;
    wire new_AGEMA_signal_13846 ;
    wire new_AGEMA_signal_13847 ;
    wire new_AGEMA_signal_13848 ;
    wire new_AGEMA_signal_13849 ;
    wire new_AGEMA_signal_13850 ;
    wire new_AGEMA_signal_13851 ;
    wire new_AGEMA_signal_13852 ;
    wire new_AGEMA_signal_13853 ;
    wire new_AGEMA_signal_13854 ;
    wire new_AGEMA_signal_13855 ;
    wire new_AGEMA_signal_13856 ;
    wire new_AGEMA_signal_13857 ;
    wire new_AGEMA_signal_13858 ;
    wire new_AGEMA_signal_13859 ;
    wire new_AGEMA_signal_13860 ;
    wire new_AGEMA_signal_13861 ;
    wire new_AGEMA_signal_13862 ;
    wire new_AGEMA_signal_13863 ;
    wire new_AGEMA_signal_13864 ;
    wire new_AGEMA_signal_13865 ;
    wire new_AGEMA_signal_13866 ;
    wire new_AGEMA_signal_13867 ;
    wire new_AGEMA_signal_13868 ;
    wire new_AGEMA_signal_13869 ;
    wire new_AGEMA_signal_13870 ;
    wire new_AGEMA_signal_13871 ;
    wire new_AGEMA_signal_13872 ;
    wire new_AGEMA_signal_13873 ;
    wire new_AGEMA_signal_13874 ;
    wire new_AGEMA_signal_13875 ;
    wire new_AGEMA_signal_13876 ;
    wire new_AGEMA_signal_13877 ;
    wire new_AGEMA_signal_13878 ;
    wire new_AGEMA_signal_13879 ;
    wire new_AGEMA_signal_13880 ;
    wire new_AGEMA_signal_13881 ;
    wire new_AGEMA_signal_13882 ;
    wire new_AGEMA_signal_13883 ;
    wire new_AGEMA_signal_13884 ;
    wire new_AGEMA_signal_13885 ;
    wire new_AGEMA_signal_13886 ;
    wire new_AGEMA_signal_13887 ;
    wire new_AGEMA_signal_13888 ;
    wire new_AGEMA_signal_13889 ;
    wire new_AGEMA_signal_13890 ;
    wire new_AGEMA_signal_13891 ;
    wire new_AGEMA_signal_13892 ;
    wire new_AGEMA_signal_13893 ;
    wire new_AGEMA_signal_13894 ;
    wire new_AGEMA_signal_13895 ;
    wire new_AGEMA_signal_13896 ;
    wire new_AGEMA_signal_13897 ;
    wire new_AGEMA_signal_13898 ;
    wire new_AGEMA_signal_13899 ;
    wire new_AGEMA_signal_13900 ;
    wire new_AGEMA_signal_13901 ;
    wire new_AGEMA_signal_13902 ;
    wire new_AGEMA_signal_13903 ;
    wire new_AGEMA_signal_13904 ;
    wire new_AGEMA_signal_13905 ;
    wire new_AGEMA_signal_13906 ;
    wire new_AGEMA_signal_13907 ;
    wire new_AGEMA_signal_13908 ;
    wire new_AGEMA_signal_13909 ;
    wire new_AGEMA_signal_13910 ;
    wire new_AGEMA_signal_13911 ;
    wire new_AGEMA_signal_13912 ;
    wire new_AGEMA_signal_13913 ;
    wire new_AGEMA_signal_13914 ;
    wire new_AGEMA_signal_13915 ;
    wire new_AGEMA_signal_13916 ;
    wire new_AGEMA_signal_13917 ;
    wire new_AGEMA_signal_13918 ;
    wire new_AGEMA_signal_13919 ;
    wire new_AGEMA_signal_13920 ;
    wire new_AGEMA_signal_13921 ;
    wire new_AGEMA_signal_13922 ;
    wire new_AGEMA_signal_13923 ;
    wire new_AGEMA_signal_13924 ;
    wire new_AGEMA_signal_13925 ;
    wire new_AGEMA_signal_13926 ;
    wire new_AGEMA_signal_13927 ;
    wire new_AGEMA_signal_13928 ;
    wire new_AGEMA_signal_13929 ;
    wire new_AGEMA_signal_13930 ;
    wire new_AGEMA_signal_13931 ;
    wire new_AGEMA_signal_13932 ;
    wire new_AGEMA_signal_13933 ;
    wire new_AGEMA_signal_13934 ;
    wire new_AGEMA_signal_13935 ;
    wire new_AGEMA_signal_13936 ;
    wire new_AGEMA_signal_13937 ;
    wire new_AGEMA_signal_13938 ;
    wire new_AGEMA_signal_13939 ;
    wire new_AGEMA_signal_13944 ;
    wire new_AGEMA_signal_13945 ;
    wire new_AGEMA_signal_13946 ;
    wire new_AGEMA_signal_13947 ;
    wire new_AGEMA_signal_13948 ;
    wire new_AGEMA_signal_13949 ;
    wire new_AGEMA_signal_13950 ;
    wire new_AGEMA_signal_13951 ;
    wire new_AGEMA_signal_13952 ;
    wire new_AGEMA_signal_13953 ;
    wire new_AGEMA_signal_13954 ;
    wire new_AGEMA_signal_13955 ;
    wire new_AGEMA_signal_13956 ;
    wire new_AGEMA_signal_13957 ;
    wire new_AGEMA_signal_13958 ;
    wire new_AGEMA_signal_13959 ;
    wire new_AGEMA_signal_13960 ;
    wire new_AGEMA_signal_13961 ;
    wire new_AGEMA_signal_13962 ;
    wire new_AGEMA_signal_13963 ;
    wire new_AGEMA_signal_13988 ;
    wire new_AGEMA_signal_13989 ;
    wire new_AGEMA_signal_13990 ;
    wire new_AGEMA_signal_13991 ;
    wire new_AGEMA_signal_13992 ;
    wire new_AGEMA_signal_13993 ;
    wire new_AGEMA_signal_13994 ;
    wire new_AGEMA_signal_13995 ;
    wire new_AGEMA_signal_13996 ;
    wire new_AGEMA_signal_13997 ;
    wire new_AGEMA_signal_13998 ;
    wire new_AGEMA_signal_13999 ;
    wire new_AGEMA_signal_14002 ;
    wire new_AGEMA_signal_14003 ;
    wire new_AGEMA_signal_14004 ;
    wire new_AGEMA_signal_14005 ;
    wire new_AGEMA_signal_14006 ;
    wire new_AGEMA_signal_14007 ;
    wire new_AGEMA_signal_14008 ;
    wire new_AGEMA_signal_14009 ;
    wire new_AGEMA_signal_14010 ;
    wire new_AGEMA_signal_14011 ;
    wire new_AGEMA_signal_14012 ;
    wire new_AGEMA_signal_14013 ;
    wire new_AGEMA_signal_14014 ;
    wire new_AGEMA_signal_14015 ;
    wire new_AGEMA_signal_14016 ;
    wire new_AGEMA_signal_14017 ;
    wire new_AGEMA_signal_14018 ;
    wire new_AGEMA_signal_14019 ;
    wire new_AGEMA_signal_14020 ;
    wire new_AGEMA_signal_14021 ;
    wire new_AGEMA_signal_14022 ;
    wire new_AGEMA_signal_14023 ;
    wire new_AGEMA_signal_14024 ;
    wire new_AGEMA_signal_14025 ;
    wire new_AGEMA_signal_14026 ;
    wire new_AGEMA_signal_14027 ;
    wire new_AGEMA_signal_14028 ;
    wire new_AGEMA_signal_14029 ;
    wire new_AGEMA_signal_14030 ;
    wire new_AGEMA_signal_14031 ;
    wire new_AGEMA_signal_14032 ;
    wire new_AGEMA_signal_14033 ;
    wire new_AGEMA_signal_14034 ;
    wire new_AGEMA_signal_14035 ;
    wire new_AGEMA_signal_14036 ;
    wire new_AGEMA_signal_14037 ;
    wire new_AGEMA_signal_14038 ;
    wire new_AGEMA_signal_14039 ;
    wire new_AGEMA_signal_14040 ;
    wire new_AGEMA_signal_14041 ;
    wire new_AGEMA_signal_14042 ;
    wire new_AGEMA_signal_14043 ;
    wire new_AGEMA_signal_14044 ;
    wire new_AGEMA_signal_14045 ;
    wire new_AGEMA_signal_14046 ;
    wire new_AGEMA_signal_14047 ;
    wire new_AGEMA_signal_14048 ;
    wire new_AGEMA_signal_14049 ;
    wire new_AGEMA_signal_14050 ;
    wire new_AGEMA_signal_14051 ;
    wire new_AGEMA_signal_14052 ;
    wire new_AGEMA_signal_14053 ;
    wire new_AGEMA_signal_14054 ;
    wire new_AGEMA_signal_14055 ;
    wire new_AGEMA_signal_14056 ;
    wire new_AGEMA_signal_14057 ;
    wire new_AGEMA_signal_14058 ;
    wire new_AGEMA_signal_14059 ;
    wire new_AGEMA_signal_14060 ;
    wire new_AGEMA_signal_14061 ;
    wire new_AGEMA_signal_14062 ;
    wire new_AGEMA_signal_14063 ;
    wire new_AGEMA_signal_14064 ;
    wire new_AGEMA_signal_14065 ;
    wire new_AGEMA_signal_14066 ;
    wire new_AGEMA_signal_14067 ;
    wire new_AGEMA_signal_14068 ;
    wire new_AGEMA_signal_14069 ;
    wire new_AGEMA_signal_14070 ;
    wire new_AGEMA_signal_14071 ;
    wire new_AGEMA_signal_14072 ;
    wire new_AGEMA_signal_14073 ;
    wire new_AGEMA_signal_14074 ;
    wire new_AGEMA_signal_14075 ;
    wire new_AGEMA_signal_14076 ;
    wire new_AGEMA_signal_14077 ;
    wire new_AGEMA_signal_14078 ;
    wire new_AGEMA_signal_14079 ;
    wire new_AGEMA_signal_14080 ;
    wire new_AGEMA_signal_14081 ;
    wire new_AGEMA_signal_14082 ;
    wire new_AGEMA_signal_14083 ;
    wire new_AGEMA_signal_14084 ;
    wire new_AGEMA_signal_14085 ;
    wire new_AGEMA_signal_14088 ;
    wire new_AGEMA_signal_14089 ;
    wire new_AGEMA_signal_14090 ;
    wire new_AGEMA_signal_14091 ;
    wire new_AGEMA_signal_14092 ;
    wire new_AGEMA_signal_14093 ;
    wire new_AGEMA_signal_14094 ;
    wire new_AGEMA_signal_14095 ;
    wire new_AGEMA_signal_14096 ;
    wire new_AGEMA_signal_14097 ;
    wire new_AGEMA_signal_14098 ;
    wire new_AGEMA_signal_14099 ;
    wire new_AGEMA_signal_14100 ;
    wire new_AGEMA_signal_14101 ;
    wire new_AGEMA_signal_14102 ;
    wire new_AGEMA_signal_14103 ;
    wire new_AGEMA_signal_14104 ;
    wire new_AGEMA_signal_14105 ;
    wire new_AGEMA_signal_14106 ;
    wire new_AGEMA_signal_14107 ;
    wire new_AGEMA_signal_14108 ;
    wire new_AGEMA_signal_14109 ;
    wire new_AGEMA_signal_14110 ;
    wire new_AGEMA_signal_14111 ;
    wire new_AGEMA_signal_14112 ;
    wire new_AGEMA_signal_14113 ;
    wire new_AGEMA_signal_14114 ;
    wire new_AGEMA_signal_14115 ;
    wire new_AGEMA_signal_14116 ;
    wire new_AGEMA_signal_14117 ;
    wire new_AGEMA_signal_14118 ;
    wire new_AGEMA_signal_14119 ;
    wire new_AGEMA_signal_14120 ;
    wire new_AGEMA_signal_14121 ;
    wire new_AGEMA_signal_14124 ;
    wire new_AGEMA_signal_14125 ;
    wire new_AGEMA_signal_14126 ;
    wire new_AGEMA_signal_14127 ;
    wire new_AGEMA_signal_14128 ;
    wire new_AGEMA_signal_14129 ;
    wire new_AGEMA_signal_14130 ;
    wire new_AGEMA_signal_14131 ;
    wire new_AGEMA_signal_14132 ;
    wire new_AGEMA_signal_14133 ;
    wire new_AGEMA_signal_14134 ;
    wire new_AGEMA_signal_14135 ;
    wire new_AGEMA_signal_14136 ;
    wire new_AGEMA_signal_14137 ;
    wire new_AGEMA_signal_14138 ;
    wire new_AGEMA_signal_14139 ;
    wire new_AGEMA_signal_14140 ;
    wire new_AGEMA_signal_14141 ;
    wire new_AGEMA_signal_14142 ;
    wire new_AGEMA_signal_14143 ;
    wire new_AGEMA_signal_14144 ;
    wire new_AGEMA_signal_14145 ;
    wire new_AGEMA_signal_14146 ;
    wire new_AGEMA_signal_14147 ;
    wire new_AGEMA_signal_14148 ;
    wire new_AGEMA_signal_14149 ;
    wire new_AGEMA_signal_14150 ;
    wire new_AGEMA_signal_14151 ;
    wire new_AGEMA_signal_14152 ;
    wire new_AGEMA_signal_14153 ;
    wire new_AGEMA_signal_14154 ;
    wire new_AGEMA_signal_14155 ;
    wire new_AGEMA_signal_14156 ;
    wire new_AGEMA_signal_14157 ;
    wire new_AGEMA_signal_14158 ;
    wire new_AGEMA_signal_14159 ;
    wire new_AGEMA_signal_14160 ;
    wire new_AGEMA_signal_14161 ;
    wire new_AGEMA_signal_14162 ;
    wire new_AGEMA_signal_14163 ;
    wire new_AGEMA_signal_14164 ;
    wire new_AGEMA_signal_14165 ;
    wire new_AGEMA_signal_14166 ;
    wire new_AGEMA_signal_14167 ;
    wire new_AGEMA_signal_14168 ;
    wire new_AGEMA_signal_14169 ;
    wire new_AGEMA_signal_14170 ;
    wire new_AGEMA_signal_14171 ;
    wire new_AGEMA_signal_14172 ;
    wire new_AGEMA_signal_14173 ;
    wire new_AGEMA_signal_14174 ;
    wire new_AGEMA_signal_14175 ;
    wire new_AGEMA_signal_14176 ;
    wire new_AGEMA_signal_14177 ;
    wire new_AGEMA_signal_14178 ;
    wire new_AGEMA_signal_14179 ;
    wire new_AGEMA_signal_14180 ;
    wire new_AGEMA_signal_14181 ;
    wire new_AGEMA_signal_14182 ;
    wire new_AGEMA_signal_14183 ;
    wire new_AGEMA_signal_14184 ;
    wire new_AGEMA_signal_14185 ;
    wire new_AGEMA_signal_14188 ;
    wire new_AGEMA_signal_14189 ;
    wire new_AGEMA_signal_14190 ;
    wire new_AGEMA_signal_14191 ;
    wire new_AGEMA_signal_14192 ;
    wire new_AGEMA_signal_14193 ;
    wire new_AGEMA_signal_14194 ;
    wire new_AGEMA_signal_14195 ;
    wire new_AGEMA_signal_14196 ;
    wire new_AGEMA_signal_14197 ;
    wire new_AGEMA_signal_14198 ;
    wire new_AGEMA_signal_14199 ;
    wire new_AGEMA_signal_14200 ;
    wire new_AGEMA_signal_14201 ;
    wire new_AGEMA_signal_14202 ;
    wire new_AGEMA_signal_14203 ;
    wire new_AGEMA_signal_14204 ;
    wire new_AGEMA_signal_14205 ;
    wire new_AGEMA_signal_14206 ;
    wire new_AGEMA_signal_14207 ;
    wire new_AGEMA_signal_14208 ;
    wire new_AGEMA_signal_14209 ;
    wire new_AGEMA_signal_14210 ;
    wire new_AGEMA_signal_14211 ;
    wire new_AGEMA_signal_14212 ;
    wire new_AGEMA_signal_14213 ;
    wire new_AGEMA_signal_14214 ;
    wire new_AGEMA_signal_14215 ;
    wire new_AGEMA_signal_14216 ;
    wire new_AGEMA_signal_14217 ;
    wire new_AGEMA_signal_14218 ;
    wire new_AGEMA_signal_14219 ;
    wire new_AGEMA_signal_14220 ;
    wire new_AGEMA_signal_14221 ;
    wire new_AGEMA_signal_14222 ;
    wire new_AGEMA_signal_14223 ;
    wire new_AGEMA_signal_14224 ;
    wire new_AGEMA_signal_14225 ;
    wire new_AGEMA_signal_14226 ;
    wire new_AGEMA_signal_14227 ;
    wire new_AGEMA_signal_14228 ;
    wire new_AGEMA_signal_14229 ;
    wire new_AGEMA_signal_14230 ;
    wire new_AGEMA_signal_14231 ;
    wire new_AGEMA_signal_14232 ;
    wire new_AGEMA_signal_14233 ;
    wire new_AGEMA_signal_14234 ;
    wire new_AGEMA_signal_14235 ;
    wire new_AGEMA_signal_14236 ;
    wire new_AGEMA_signal_14237 ;
    wire new_AGEMA_signal_14238 ;
    wire new_AGEMA_signal_14239 ;
    wire new_AGEMA_signal_14240 ;
    wire new_AGEMA_signal_14241 ;
    wire new_AGEMA_signal_14242 ;
    wire new_AGEMA_signal_14243 ;
    wire new_AGEMA_signal_14244 ;
    wire new_AGEMA_signal_14245 ;
    wire new_AGEMA_signal_14246 ;
    wire new_AGEMA_signal_14247 ;
    wire new_AGEMA_signal_14248 ;
    wire new_AGEMA_signal_14249 ;
    wire new_AGEMA_signal_14250 ;
    wire new_AGEMA_signal_14251 ;
    wire new_AGEMA_signal_14252 ;
    wire new_AGEMA_signal_14253 ;
    wire new_AGEMA_signal_14254 ;
    wire new_AGEMA_signal_14255 ;
    wire new_AGEMA_signal_14256 ;
    wire new_AGEMA_signal_14257 ;
    wire new_AGEMA_signal_14258 ;
    wire new_AGEMA_signal_14259 ;
    wire new_AGEMA_signal_14260 ;
    wire new_AGEMA_signal_14261 ;
    wire new_AGEMA_signal_14262 ;
    wire new_AGEMA_signal_14263 ;
    wire new_AGEMA_signal_14264 ;
    wire new_AGEMA_signal_14265 ;
    wire new_AGEMA_signal_14266 ;
    wire new_AGEMA_signal_14267 ;
    wire new_AGEMA_signal_14268 ;
    wire new_AGEMA_signal_14269 ;
    wire new_AGEMA_signal_14270 ;
    wire new_AGEMA_signal_14271 ;
    wire new_AGEMA_signal_14274 ;
    wire new_AGEMA_signal_14275 ;
    wire new_AGEMA_signal_14276 ;
    wire new_AGEMA_signal_14277 ;
    wire new_AGEMA_signal_14278 ;
    wire new_AGEMA_signal_14279 ;
    wire new_AGEMA_signal_14280 ;
    wire new_AGEMA_signal_14281 ;
    wire new_AGEMA_signal_14282 ;
    wire new_AGEMA_signal_14283 ;
    wire new_AGEMA_signal_14284 ;
    wire new_AGEMA_signal_14285 ;
    wire new_AGEMA_signal_14286 ;
    wire new_AGEMA_signal_14287 ;
    wire new_AGEMA_signal_14288 ;
    wire new_AGEMA_signal_14289 ;
    wire new_AGEMA_signal_14290 ;
    wire new_AGEMA_signal_14291 ;
    wire new_AGEMA_signal_14292 ;
    wire new_AGEMA_signal_14293 ;
    wire new_AGEMA_signal_14294 ;
    wire new_AGEMA_signal_14295 ;
    wire new_AGEMA_signal_14296 ;
    wire new_AGEMA_signal_14297 ;
    wire new_AGEMA_signal_14298 ;
    wire new_AGEMA_signal_14299 ;
    wire new_AGEMA_signal_14300 ;
    wire new_AGEMA_signal_14301 ;
    wire new_AGEMA_signal_14302 ;
    wire new_AGEMA_signal_14303 ;
    wire new_AGEMA_signal_14304 ;
    wire new_AGEMA_signal_14305 ;
    wire new_AGEMA_signal_14306 ;
    wire new_AGEMA_signal_14307 ;
    wire new_AGEMA_signal_14310 ;
    wire new_AGEMA_signal_14311 ;
    wire new_AGEMA_signal_14312 ;
    wire new_AGEMA_signal_14313 ;
    wire new_AGEMA_signal_14314 ;
    wire new_AGEMA_signal_14315 ;
    wire new_AGEMA_signal_14316 ;
    wire new_AGEMA_signal_14317 ;
    wire new_AGEMA_signal_14318 ;
    wire new_AGEMA_signal_14319 ;
    wire new_AGEMA_signal_14320 ;
    wire new_AGEMA_signal_14321 ;
    wire new_AGEMA_signal_14322 ;
    wire new_AGEMA_signal_14323 ;
    wire new_AGEMA_signal_14324 ;
    wire new_AGEMA_signal_14325 ;
    wire new_AGEMA_signal_14326 ;
    wire new_AGEMA_signal_14327 ;
    wire new_AGEMA_signal_14328 ;
    wire new_AGEMA_signal_14329 ;
    wire new_AGEMA_signal_14330 ;
    wire new_AGEMA_signal_14331 ;
    wire new_AGEMA_signal_14332 ;
    wire new_AGEMA_signal_14333 ;
    wire new_AGEMA_signal_14334 ;
    wire new_AGEMA_signal_14335 ;
    wire new_AGEMA_signal_14336 ;
    wire new_AGEMA_signal_14337 ;
    wire new_AGEMA_signal_14338 ;
    wire new_AGEMA_signal_14339 ;
    wire new_AGEMA_signal_14340 ;
    wire new_AGEMA_signal_14341 ;
    wire new_AGEMA_signal_14342 ;
    wire new_AGEMA_signal_14343 ;
    wire new_AGEMA_signal_14344 ;
    wire new_AGEMA_signal_14345 ;
    wire new_AGEMA_signal_14346 ;
    wire new_AGEMA_signal_14347 ;
    wire new_AGEMA_signal_14348 ;
    wire new_AGEMA_signal_14349 ;
    wire new_AGEMA_signal_14350 ;
    wire new_AGEMA_signal_14351 ;
    wire new_AGEMA_signal_14352 ;
    wire new_AGEMA_signal_14353 ;
    wire new_AGEMA_signal_14354 ;
    wire new_AGEMA_signal_14355 ;
    wire new_AGEMA_signal_14356 ;
    wire new_AGEMA_signal_14357 ;
    wire new_AGEMA_signal_14358 ;
    wire new_AGEMA_signal_14359 ;
    wire new_AGEMA_signal_14360 ;
    wire new_AGEMA_signal_14361 ;
    wire new_AGEMA_signal_14362 ;
    wire new_AGEMA_signal_14363 ;
    wire new_AGEMA_signal_14364 ;
    wire new_AGEMA_signal_14365 ;
    wire new_AGEMA_signal_14366 ;
    wire new_AGEMA_signal_14367 ;
    wire new_AGEMA_signal_14368 ;
    wire new_AGEMA_signal_14369 ;
    wire new_AGEMA_signal_14370 ;
    wire new_AGEMA_signal_14371 ;
    wire new_AGEMA_signal_14372 ;
    wire new_AGEMA_signal_14373 ;
    wire new_AGEMA_signal_14374 ;
    wire new_AGEMA_signal_14375 ;
    wire new_AGEMA_signal_14376 ;
    wire new_AGEMA_signal_14377 ;
    wire new_AGEMA_signal_14378 ;
    wire new_AGEMA_signal_14379 ;
    wire new_AGEMA_signal_14380 ;
    wire new_AGEMA_signal_14381 ;
    wire new_AGEMA_signal_14382 ;
    wire new_AGEMA_signal_14383 ;
    wire new_AGEMA_signal_14410 ;
    wire new_AGEMA_signal_14411 ;
    wire new_AGEMA_signal_14412 ;
    wire new_AGEMA_signal_14413 ;
    wire new_AGEMA_signal_14414 ;
    wire new_AGEMA_signal_14415 ;
    wire new_AGEMA_signal_14416 ;
    wire new_AGEMA_signal_14417 ;
    wire new_AGEMA_signal_14418 ;
    wire new_AGEMA_signal_14419 ;
    wire new_AGEMA_signal_14420 ;
    wire new_AGEMA_signal_14421 ;
    wire new_AGEMA_signal_14422 ;
    wire new_AGEMA_signal_14423 ;
    wire new_AGEMA_signal_14424 ;
    wire new_AGEMA_signal_14425 ;
    wire new_AGEMA_signal_14426 ;
    wire new_AGEMA_signal_14427 ;
    wire new_AGEMA_signal_14428 ;
    wire new_AGEMA_signal_14429 ;
    wire new_AGEMA_signal_14430 ;
    wire new_AGEMA_signal_14431 ;
    wire new_AGEMA_signal_14432 ;
    wire new_AGEMA_signal_14433 ;
    wire new_AGEMA_signal_14434 ;
    wire new_AGEMA_signal_14435 ;
    wire new_AGEMA_signal_14436 ;
    wire new_AGEMA_signal_14437 ;
    wire new_AGEMA_signal_14438 ;
    wire new_AGEMA_signal_14439 ;
    wire new_AGEMA_signal_14440 ;
    wire new_AGEMA_signal_14441 ;
    wire new_AGEMA_signal_14442 ;
    wire new_AGEMA_signal_14443 ;
    wire new_AGEMA_signal_14444 ;
    wire new_AGEMA_signal_14445 ;
    wire new_AGEMA_signal_14446 ;
    wire new_AGEMA_signal_14447 ;
    wire new_AGEMA_signal_14448 ;
    wire new_AGEMA_signal_14449 ;
    wire new_AGEMA_signal_14450 ;
    wire new_AGEMA_signal_14451 ;
    wire new_AGEMA_signal_14452 ;
    wire new_AGEMA_signal_14453 ;
    wire new_AGEMA_signal_14454 ;
    wire new_AGEMA_signal_14455 ;
    wire new_AGEMA_signal_14456 ;
    wire new_AGEMA_signal_14457 ;
    wire new_AGEMA_signal_14458 ;
    wire new_AGEMA_signal_14459 ;
    wire new_AGEMA_signal_14460 ;
    wire new_AGEMA_signal_14461 ;
    wire new_AGEMA_signal_14462 ;
    wire new_AGEMA_signal_14463 ;
    wire new_AGEMA_signal_14464 ;
    wire new_AGEMA_signal_14465 ;
    wire new_AGEMA_signal_14466 ;
    wire new_AGEMA_signal_14467 ;
    wire new_AGEMA_signal_14468 ;
    wire new_AGEMA_signal_14469 ;
    wire new_AGEMA_signal_14470 ;
    wire new_AGEMA_signal_14471 ;
    wire new_AGEMA_signal_14472 ;
    wire new_AGEMA_signal_14473 ;
    wire new_AGEMA_signal_14476 ;
    wire new_AGEMA_signal_14477 ;
    wire new_AGEMA_signal_14478 ;
    wire new_AGEMA_signal_14479 ;
    wire new_AGEMA_signal_14480 ;
    wire new_AGEMA_signal_14481 ;
    wire new_AGEMA_signal_14482 ;
    wire new_AGEMA_signal_14483 ;
    wire new_AGEMA_signal_14484 ;
    wire new_AGEMA_signal_14485 ;
    wire new_AGEMA_signal_14486 ;
    wire new_AGEMA_signal_14487 ;
    wire new_AGEMA_signal_14488 ;
    wire new_AGEMA_signal_14489 ;
    wire new_AGEMA_signal_14490 ;
    wire new_AGEMA_signal_14491 ;
    wire new_AGEMA_signal_14492 ;
    wire new_AGEMA_signal_14493 ;
    wire new_AGEMA_signal_14494 ;
    wire new_AGEMA_signal_14495 ;
    wire new_AGEMA_signal_14496 ;
    wire new_AGEMA_signal_14497 ;
    wire new_AGEMA_signal_14498 ;
    wire new_AGEMA_signal_14499 ;
    wire new_AGEMA_signal_14500 ;
    wire new_AGEMA_signal_14501 ;
    wire new_AGEMA_signal_14502 ;
    wire new_AGEMA_signal_14503 ;
    wire new_AGEMA_signal_14504 ;
    wire new_AGEMA_signal_14505 ;
    wire new_AGEMA_signal_14506 ;
    wire new_AGEMA_signal_14507 ;
    wire new_AGEMA_signal_14508 ;
    wire new_AGEMA_signal_14509 ;
    wire new_AGEMA_signal_14510 ;
    wire new_AGEMA_signal_14511 ;
    wire new_AGEMA_signal_14512 ;
    wire new_AGEMA_signal_14513 ;
    wire new_AGEMA_signal_14514 ;
    wire new_AGEMA_signal_14515 ;
    wire new_AGEMA_signal_14516 ;
    wire new_AGEMA_signal_14517 ;
    wire new_AGEMA_signal_14518 ;
    wire new_AGEMA_signal_14519 ;
    wire new_AGEMA_signal_14522 ;
    wire new_AGEMA_signal_14523 ;
    wire new_AGEMA_signal_14524 ;
    wire new_AGEMA_signal_14525 ;
    wire new_AGEMA_signal_14526 ;
    wire new_AGEMA_signal_14527 ;
    wire new_AGEMA_signal_14528 ;
    wire new_AGEMA_signal_14529 ;
    wire new_AGEMA_signal_14530 ;
    wire new_AGEMA_signal_14531 ;
    wire new_AGEMA_signal_14532 ;
    wire new_AGEMA_signal_14533 ;
    wire new_AGEMA_signal_14534 ;
    wire new_AGEMA_signal_14535 ;
    wire new_AGEMA_signal_14536 ;
    wire new_AGEMA_signal_14537 ;
    wire new_AGEMA_signal_14538 ;
    wire new_AGEMA_signal_14539 ;
    wire new_AGEMA_signal_14540 ;
    wire new_AGEMA_signal_14541 ;
    wire new_AGEMA_signal_14542 ;
    wire new_AGEMA_signal_14543 ;
    wire new_AGEMA_signal_14544 ;
    wire new_AGEMA_signal_14545 ;
    wire new_AGEMA_signal_14546 ;
    wire new_AGEMA_signal_14547 ;
    wire new_AGEMA_signal_14548 ;
    wire new_AGEMA_signal_14549 ;
    wire new_AGEMA_signal_14550 ;
    wire new_AGEMA_signal_14551 ;
    wire new_AGEMA_signal_14552 ;
    wire new_AGEMA_signal_14553 ;
    wire new_AGEMA_signal_14554 ;
    wire new_AGEMA_signal_14555 ;
    wire new_AGEMA_signal_14556 ;
    wire new_AGEMA_signal_14557 ;
    wire new_AGEMA_signal_14558 ;
    wire new_AGEMA_signal_14559 ;
    wire new_AGEMA_signal_14560 ;
    wire new_AGEMA_signal_14561 ;
    wire new_AGEMA_signal_14562 ;
    wire new_AGEMA_signal_14563 ;
    wire new_AGEMA_signal_14564 ;
    wire new_AGEMA_signal_14565 ;
    wire new_AGEMA_signal_14566 ;
    wire new_AGEMA_signal_14567 ;
    wire new_AGEMA_signal_14570 ;
    wire new_AGEMA_signal_14571 ;
    wire new_AGEMA_signal_14572 ;
    wire new_AGEMA_signal_14573 ;
    wire new_AGEMA_signal_14574 ;
    wire new_AGEMA_signal_14575 ;
    wire new_AGEMA_signal_14576 ;
    wire new_AGEMA_signal_14577 ;
    wire new_AGEMA_signal_14578 ;
    wire new_AGEMA_signal_14579 ;
    wire new_AGEMA_signal_14580 ;
    wire new_AGEMA_signal_14581 ;
    wire new_AGEMA_signal_14582 ;
    wire new_AGEMA_signal_14583 ;
    wire new_AGEMA_signal_14584 ;
    wire new_AGEMA_signal_14585 ;
    wire new_AGEMA_signal_14586 ;
    wire new_AGEMA_signal_14587 ;
    wire new_AGEMA_signal_14588 ;
    wire new_AGEMA_signal_14589 ;
    wire new_AGEMA_signal_14590 ;
    wire new_AGEMA_signal_14591 ;
    wire new_AGEMA_signal_14592 ;
    wire new_AGEMA_signal_14593 ;
    wire new_AGEMA_signal_14594 ;
    wire new_AGEMA_signal_14595 ;
    wire new_AGEMA_signal_14596 ;
    wire new_AGEMA_signal_14597 ;
    wire new_AGEMA_signal_14598 ;
    wire new_AGEMA_signal_14599 ;
    wire new_AGEMA_signal_14600 ;
    wire new_AGEMA_signal_14601 ;
    wire new_AGEMA_signal_14602 ;
    wire new_AGEMA_signal_14603 ;
    wire new_AGEMA_signal_14604 ;
    wire new_AGEMA_signal_14605 ;
    wire new_AGEMA_signal_14608 ;
    wire new_AGEMA_signal_14609 ;
    wire new_AGEMA_signal_14610 ;
    wire new_AGEMA_signal_14611 ;
    wire new_AGEMA_signal_14612 ;
    wire new_AGEMA_signal_14613 ;
    wire new_AGEMA_signal_14614 ;
    wire new_AGEMA_signal_14615 ;
    wire new_AGEMA_signal_14616 ;
    wire new_AGEMA_signal_14617 ;
    wire new_AGEMA_signal_14618 ;
    wire new_AGEMA_signal_14619 ;
    wire new_AGEMA_signal_14620 ;
    wire new_AGEMA_signal_14621 ;
    wire new_AGEMA_signal_14622 ;
    wire new_AGEMA_signal_14623 ;
    wire new_AGEMA_signal_14624 ;
    wire new_AGEMA_signal_14625 ;
    wire new_AGEMA_signal_14626 ;
    wire new_AGEMA_signal_14627 ;
    wire new_AGEMA_signal_14628 ;
    wire new_AGEMA_signal_14629 ;
    wire new_AGEMA_signal_14630 ;
    wire new_AGEMA_signal_14631 ;
    wire new_AGEMA_signal_14632 ;
    wire new_AGEMA_signal_14633 ;
    wire new_AGEMA_signal_14634 ;
    wire new_AGEMA_signal_14635 ;
    wire new_AGEMA_signal_14636 ;
    wire new_AGEMA_signal_14637 ;
    wire new_AGEMA_signal_14638 ;
    wire new_AGEMA_signal_14639 ;
    wire new_AGEMA_signal_14640 ;
    wire new_AGEMA_signal_14641 ;
    wire new_AGEMA_signal_14642 ;
    wire new_AGEMA_signal_14643 ;
    wire new_AGEMA_signal_14644 ;
    wire new_AGEMA_signal_14645 ;
    wire new_AGEMA_signal_14646 ;
    wire new_AGEMA_signal_14647 ;
    wire new_AGEMA_signal_14648 ;
    wire new_AGEMA_signal_14649 ;
    wire new_AGEMA_signal_14650 ;
    wire new_AGEMA_signal_14651 ;
    wire new_AGEMA_signal_14652 ;
    wire new_AGEMA_signal_14653 ;
    wire new_AGEMA_signal_14654 ;
    wire new_AGEMA_signal_14655 ;
    wire new_AGEMA_signal_14656 ;
    wire new_AGEMA_signal_14657 ;
    wire new_AGEMA_signal_14658 ;
    wire new_AGEMA_signal_14659 ;
    wire new_AGEMA_signal_14660 ;
    wire new_AGEMA_signal_14661 ;
    wire new_AGEMA_signal_14662 ;
    wire new_AGEMA_signal_14663 ;
    wire new_AGEMA_signal_14664 ;
    wire new_AGEMA_signal_14665 ;
    wire new_AGEMA_signal_14666 ;
    wire new_AGEMA_signal_14667 ;
    wire new_AGEMA_signal_14668 ;
    wire new_AGEMA_signal_14669 ;
    wire new_AGEMA_signal_14670 ;
    wire new_AGEMA_signal_14671 ;
    wire new_AGEMA_signal_14674 ;
    wire new_AGEMA_signal_14675 ;
    wire new_AGEMA_signal_14676 ;
    wire new_AGEMA_signal_14677 ;
    wire new_AGEMA_signal_14678 ;
    wire new_AGEMA_signal_14679 ;
    wire new_AGEMA_signal_14680 ;
    wire new_AGEMA_signal_14681 ;
    wire new_AGEMA_signal_14682 ;
    wire new_AGEMA_signal_14683 ;
    wire new_AGEMA_signal_14684 ;
    wire new_AGEMA_signal_14685 ;
    wire new_AGEMA_signal_14686 ;
    wire new_AGEMA_signal_14687 ;
    wire new_AGEMA_signal_14688 ;
    wire new_AGEMA_signal_14689 ;
    wire new_AGEMA_signal_14690 ;
    wire new_AGEMA_signal_14691 ;
    wire new_AGEMA_signal_14692 ;
    wire new_AGEMA_signal_14693 ;
    wire new_AGEMA_signal_14694 ;
    wire new_AGEMA_signal_14695 ;
    wire new_AGEMA_signal_14696 ;
    wire new_AGEMA_signal_14697 ;
    wire new_AGEMA_signal_14698 ;
    wire new_AGEMA_signal_14699 ;
    wire new_AGEMA_signal_14700 ;
    wire new_AGEMA_signal_14701 ;
    wire new_AGEMA_signal_14702 ;
    wire new_AGEMA_signal_14703 ;
    wire new_AGEMA_signal_14704 ;
    wire new_AGEMA_signal_14705 ;
    wire new_AGEMA_signal_14706 ;
    wire new_AGEMA_signal_14707 ;
    wire new_AGEMA_signal_14708 ;
    wire new_AGEMA_signal_14709 ;
    wire new_AGEMA_signal_14710 ;
    wire new_AGEMA_signal_14711 ;
    wire new_AGEMA_signal_14712 ;
    wire new_AGEMA_signal_14713 ;
    wire new_AGEMA_signal_14714 ;
    wire new_AGEMA_signal_14715 ;
    wire new_AGEMA_signal_14716 ;
    wire new_AGEMA_signal_14717 ;
    wire new_AGEMA_signal_14720 ;
    wire new_AGEMA_signal_14721 ;
    wire new_AGEMA_signal_14722 ;
    wire new_AGEMA_signal_14723 ;
    wire new_AGEMA_signal_14724 ;
    wire new_AGEMA_signal_14725 ;
    wire new_AGEMA_signal_14726 ;
    wire new_AGEMA_signal_14727 ;
    wire new_AGEMA_signal_14728 ;
    wire new_AGEMA_signal_14729 ;
    wire new_AGEMA_signal_14730 ;
    wire new_AGEMA_signal_14731 ;
    wire new_AGEMA_signal_14732 ;
    wire new_AGEMA_signal_14733 ;
    wire new_AGEMA_signal_14734 ;
    wire new_AGEMA_signal_14735 ;
    wire new_AGEMA_signal_14736 ;
    wire new_AGEMA_signal_14737 ;
    wire new_AGEMA_signal_14738 ;
    wire new_AGEMA_signal_14739 ;
    wire new_AGEMA_signal_14740 ;
    wire new_AGEMA_signal_14741 ;
    wire new_AGEMA_signal_14742 ;
    wire new_AGEMA_signal_14743 ;
    wire new_AGEMA_signal_14744 ;
    wire new_AGEMA_signal_14745 ;
    wire new_AGEMA_signal_14746 ;
    wire new_AGEMA_signal_14747 ;
    wire new_AGEMA_signal_14748 ;
    wire new_AGEMA_signal_14749 ;
    wire new_AGEMA_signal_14750 ;
    wire new_AGEMA_signal_14751 ;
    wire new_AGEMA_signal_14752 ;
    wire new_AGEMA_signal_14753 ;
    wire new_AGEMA_signal_14754 ;
    wire new_AGEMA_signal_14755 ;
    wire new_AGEMA_signal_14756 ;
    wire new_AGEMA_signal_14757 ;
    wire new_AGEMA_signal_14758 ;
    wire new_AGEMA_signal_14759 ;
    wire new_AGEMA_signal_14760 ;
    wire new_AGEMA_signal_14761 ;
    wire new_AGEMA_signal_14762 ;
    wire new_AGEMA_signal_14763 ;
    wire new_AGEMA_signal_14764 ;
    wire new_AGEMA_signal_14765 ;
    wire new_AGEMA_signal_14768 ;
    wire new_AGEMA_signal_14769 ;
    wire new_AGEMA_signal_14770 ;
    wire new_AGEMA_signal_14771 ;
    wire new_AGEMA_signal_14772 ;
    wire new_AGEMA_signal_14773 ;
    wire new_AGEMA_signal_14774 ;
    wire new_AGEMA_signal_14775 ;
    wire new_AGEMA_signal_14776 ;
    wire new_AGEMA_signal_14777 ;
    wire new_AGEMA_signal_14778 ;
    wire new_AGEMA_signal_14779 ;
    wire new_AGEMA_signal_14780 ;
    wire new_AGEMA_signal_14781 ;
    wire new_AGEMA_signal_14782 ;
    wire new_AGEMA_signal_14783 ;
    wire new_AGEMA_signal_14784 ;
    wire new_AGEMA_signal_14785 ;
    wire new_AGEMA_signal_14786 ;
    wire new_AGEMA_signal_14787 ;
    wire new_AGEMA_signal_14788 ;
    wire new_AGEMA_signal_14789 ;
    wire new_AGEMA_signal_14790 ;
    wire new_AGEMA_signal_14791 ;
    wire new_AGEMA_signal_14792 ;
    wire new_AGEMA_signal_14793 ;
    wire new_AGEMA_signal_14794 ;
    wire new_AGEMA_signal_14795 ;
    wire new_AGEMA_signal_14796 ;
    wire new_AGEMA_signal_14797 ;
    wire new_AGEMA_signal_14798 ;
    wire new_AGEMA_signal_14799 ;
    wire new_AGEMA_signal_14800 ;
    wire new_AGEMA_signal_14801 ;
    wire new_AGEMA_signal_14802 ;
    wire new_AGEMA_signal_14803 ;
    wire new_AGEMA_signal_14824 ;
    wire new_AGEMA_signal_14825 ;
    wire new_AGEMA_signal_14826 ;
    wire new_AGEMA_signal_14827 ;
    wire new_AGEMA_signal_14828 ;
    wire new_AGEMA_signal_14829 ;
    wire new_AGEMA_signal_14830 ;
    wire new_AGEMA_signal_14831 ;
    wire new_AGEMA_signal_14832 ;
    wire new_AGEMA_signal_14833 ;
    wire new_AGEMA_signal_14834 ;
    wire new_AGEMA_signal_14835 ;
    wire new_AGEMA_signal_14836 ;
    wire new_AGEMA_signal_14837 ;
    wire new_AGEMA_signal_14838 ;
    wire new_AGEMA_signal_14839 ;
    wire new_AGEMA_signal_14840 ;
    wire new_AGEMA_signal_14841 ;
    wire new_AGEMA_signal_14842 ;
    wire new_AGEMA_signal_14843 ;
    wire new_AGEMA_signal_14844 ;
    wire new_AGEMA_signal_14845 ;
    wire new_AGEMA_signal_14846 ;
    wire new_AGEMA_signal_14847 ;
    wire new_AGEMA_signal_14848 ;
    wire new_AGEMA_signal_14849 ;
    wire new_AGEMA_signal_14850 ;
    wire new_AGEMA_signal_14851 ;
    wire new_AGEMA_signal_14852 ;
    wire new_AGEMA_signal_14853 ;
    wire new_AGEMA_signal_14854 ;
    wire new_AGEMA_signal_14855 ;
    wire new_AGEMA_signal_14856 ;
    wire new_AGEMA_signal_14857 ;
    wire new_AGEMA_signal_14858 ;
    wire new_AGEMA_signal_14859 ;
    wire new_AGEMA_signal_14892 ;
    wire new_AGEMA_signal_14893 ;
    wire new_AGEMA_signal_14896 ;
    wire new_AGEMA_signal_14897 ;
    wire new_AGEMA_signal_14898 ;
    wire new_AGEMA_signal_14899 ;
    wire new_AGEMA_signal_14900 ;
    wire new_AGEMA_signal_14901 ;
    wire new_AGEMA_signal_14902 ;
    wire new_AGEMA_signal_14903 ;
    wire new_AGEMA_signal_14904 ;
    wire new_AGEMA_signal_14905 ;
    wire new_AGEMA_signal_14910 ;
    wire new_AGEMA_signal_14911 ;
    wire new_AGEMA_signal_14912 ;
    wire new_AGEMA_signal_14913 ;
    wire new_AGEMA_signal_14914 ;
    wire new_AGEMA_signal_14915 ;
    wire new_AGEMA_signal_14916 ;
    wire new_AGEMA_signal_14917 ;
    wire new_AGEMA_signal_14918 ;
    wire new_AGEMA_signal_14919 ;
    wire new_AGEMA_signal_14920 ;
    wire new_AGEMA_signal_14921 ;
    wire new_AGEMA_signal_14922 ;
    wire new_AGEMA_signal_14923 ;
    wire new_AGEMA_signal_14924 ;
    wire new_AGEMA_signal_14925 ;
    wire new_AGEMA_signal_14926 ;
    wire new_AGEMA_signal_14927 ;
    wire new_AGEMA_signal_14928 ;
    wire new_AGEMA_signal_14929 ;
    wire new_AGEMA_signal_14930 ;
    wire new_AGEMA_signal_14931 ;
    wire new_AGEMA_signal_14932 ;
    wire new_AGEMA_signal_14933 ;
    wire new_AGEMA_signal_14934 ;
    wire new_AGEMA_signal_14935 ;
    wire new_AGEMA_signal_14938 ;
    wire new_AGEMA_signal_14939 ;
    wire new_AGEMA_signal_14944 ;
    wire new_AGEMA_signal_14945 ;
    wire new_AGEMA_signal_14946 ;
    wire new_AGEMA_signal_14947 ;
    wire new_AGEMA_signal_14950 ;
    wire new_AGEMA_signal_14951 ;
    wire new_AGEMA_signal_14952 ;
    wire new_AGEMA_signal_14953 ;
    wire new_AGEMA_signal_14954 ;
    wire new_AGEMA_signal_14955 ;
    wire new_AGEMA_signal_14956 ;
    wire new_AGEMA_signal_14957 ;
    wire new_AGEMA_signal_14958 ;
    wire new_AGEMA_signal_14959 ;
    wire new_AGEMA_signal_14960 ;
    wire new_AGEMA_signal_14961 ;
    wire new_AGEMA_signal_14962 ;
    wire new_AGEMA_signal_14963 ;
    wire new_AGEMA_signal_14966 ;
    wire new_AGEMA_signal_14967 ;
    wire new_AGEMA_signal_14970 ;
    wire new_AGEMA_signal_14971 ;
    wire new_AGEMA_signal_14972 ;
    wire new_AGEMA_signal_14973 ;
    wire new_AGEMA_signal_14974 ;
    wire new_AGEMA_signal_14975 ;
    wire new_AGEMA_signal_14976 ;
    wire new_AGEMA_signal_14977 ;
    wire new_AGEMA_signal_14978 ;
    wire new_AGEMA_signal_14979 ;
    wire new_AGEMA_signal_14980 ;
    wire new_AGEMA_signal_14981 ;
    wire new_AGEMA_signal_14982 ;
    wire new_AGEMA_signal_14983 ;
    wire new_AGEMA_signal_14988 ;
    wire new_AGEMA_signal_14989 ;
    wire new_AGEMA_signal_14994 ;
    wire new_AGEMA_signal_14995 ;
    wire new_AGEMA_signal_14996 ;
    wire new_AGEMA_signal_14997 ;
    wire new_AGEMA_signal_14998 ;
    wire new_AGEMA_signal_14999 ;
    wire new_AGEMA_signal_15000 ;
    wire new_AGEMA_signal_15001 ;
    wire new_AGEMA_signal_15002 ;
    wire new_AGEMA_signal_15003 ;
    wire new_AGEMA_signal_15004 ;
    wire new_AGEMA_signal_15005 ;
    wire new_AGEMA_signal_15006 ;
    wire new_AGEMA_signal_15007 ;
    wire new_AGEMA_signal_15008 ;
    wire new_AGEMA_signal_15009 ;
    wire new_AGEMA_signal_15010 ;
    wire new_AGEMA_signal_15011 ;
    wire new_AGEMA_signal_15012 ;
    wire new_AGEMA_signal_15013 ;
    wire new_AGEMA_signal_15014 ;
    wire new_AGEMA_signal_15015 ;
    wire new_AGEMA_signal_15016 ;
    wire new_AGEMA_signal_15017 ;
    wire new_AGEMA_signal_15018 ;
    wire new_AGEMA_signal_15019 ;
    wire new_AGEMA_signal_15020 ;
    wire new_AGEMA_signal_15021 ;
    wire new_AGEMA_signal_15022 ;
    wire new_AGEMA_signal_15023 ;
    wire new_AGEMA_signal_15024 ;
    wire new_AGEMA_signal_15025 ;
    wire new_AGEMA_signal_15026 ;
    wire new_AGEMA_signal_15027 ;
    wire new_AGEMA_signal_15028 ;
    wire new_AGEMA_signal_15029 ;
    wire new_AGEMA_signal_15030 ;
    wire new_AGEMA_signal_15031 ;
    wire new_AGEMA_signal_15032 ;
    wire new_AGEMA_signal_15033 ;
    wire new_AGEMA_signal_15034 ;
    wire new_AGEMA_signal_15035 ;
    wire new_AGEMA_signal_15040 ;
    wire new_AGEMA_signal_15041 ;
    wire new_AGEMA_signal_15044 ;
    wire new_AGEMA_signal_15045 ;
    wire new_AGEMA_signal_15046 ;
    wire new_AGEMA_signal_15047 ;
    wire new_AGEMA_signal_15048 ;
    wire new_AGEMA_signal_15049 ;
    wire new_AGEMA_signal_15050 ;
    wire new_AGEMA_signal_15051 ;
    wire new_AGEMA_signal_15052 ;
    wire new_AGEMA_signal_15053 ;
    wire new_AGEMA_signal_15056 ;
    wire new_AGEMA_signal_15057 ;
    wire new_AGEMA_signal_15062 ;
    wire new_AGEMA_signal_15063 ;
    wire new_AGEMA_signal_15064 ;
    wire new_AGEMA_signal_15065 ;
    wire new_AGEMA_signal_15066 ;
    wire new_AGEMA_signal_15067 ;
    wire new_AGEMA_signal_15068 ;
    wire new_AGEMA_signal_15069 ;
    wire new_AGEMA_signal_15070 ;
    wire new_AGEMA_signal_15071 ;
    wire new_AGEMA_signal_15072 ;
    wire new_AGEMA_signal_15073 ;
    wire new_AGEMA_signal_15074 ;
    wire new_AGEMA_signal_15075 ;
    wire new_AGEMA_signal_15076 ;
    wire new_AGEMA_signal_15077 ;
    wire new_AGEMA_signal_15078 ;
    wire new_AGEMA_signal_15079 ;
    wire new_AGEMA_signal_15080 ;
    wire new_AGEMA_signal_15081 ;
    wire new_AGEMA_signal_15082 ;
    wire new_AGEMA_signal_15083 ;
    wire new_AGEMA_signal_15086 ;
    wire new_AGEMA_signal_15087 ;
    wire new_AGEMA_signal_15088 ;
    wire new_AGEMA_signal_15089 ;
    wire new_AGEMA_signal_15090 ;
    wire new_AGEMA_signal_15091 ;
    wire new_AGEMA_signal_15092 ;
    wire new_AGEMA_signal_15093 ;
    wire new_AGEMA_signal_15094 ;
    wire new_AGEMA_signal_15095 ;
    wire new_AGEMA_signal_15100 ;
    wire new_AGEMA_signal_15101 ;
    wire new_AGEMA_signal_15102 ;
    wire new_AGEMA_signal_15103 ;
    wire new_AGEMA_signal_15104 ;
    wire new_AGEMA_signal_15105 ;
    wire new_AGEMA_signal_15106 ;
    wire new_AGEMA_signal_15107 ;
    wire new_AGEMA_signal_15108 ;
    wire new_AGEMA_signal_15109 ;
    wire new_AGEMA_signal_15110 ;
    wire new_AGEMA_signal_15111 ;
    wire new_AGEMA_signal_15112 ;
    wire new_AGEMA_signal_15113 ;
    wire new_AGEMA_signal_15114 ;
    wire new_AGEMA_signal_15115 ;
    wire new_AGEMA_signal_15116 ;
    wire new_AGEMA_signal_15117 ;
    wire new_AGEMA_signal_15118 ;
    wire new_AGEMA_signal_15119 ;
    wire new_AGEMA_signal_15120 ;
    wire new_AGEMA_signal_15121 ;
    wire new_AGEMA_signal_15122 ;
    wire new_AGEMA_signal_15123 ;
    wire new_AGEMA_signal_15124 ;
    wire new_AGEMA_signal_15125 ;
    wire new_AGEMA_signal_15128 ;
    wire new_AGEMA_signal_15129 ;
    wire new_AGEMA_signal_15134 ;
    wire new_AGEMA_signal_15135 ;
    wire new_AGEMA_signal_15136 ;
    wire new_AGEMA_signal_15137 ;
    wire new_AGEMA_signal_15140 ;
    wire new_AGEMA_signal_15141 ;
    wire new_AGEMA_signal_15142 ;
    wire new_AGEMA_signal_15143 ;
    wire new_AGEMA_signal_15144 ;
    wire new_AGEMA_signal_15145 ;
    wire new_AGEMA_signal_15146 ;
    wire new_AGEMA_signal_15147 ;
    wire new_AGEMA_signal_15148 ;
    wire new_AGEMA_signal_15149 ;
    wire new_AGEMA_signal_15150 ;
    wire new_AGEMA_signal_15151 ;
    wire new_AGEMA_signal_15152 ;
    wire new_AGEMA_signal_15153 ;
    wire new_AGEMA_signal_15156 ;
    wire new_AGEMA_signal_15157 ;
    wire new_AGEMA_signal_15160 ;
    wire new_AGEMA_signal_15161 ;
    wire new_AGEMA_signal_15162 ;
    wire new_AGEMA_signal_15163 ;
    wire new_AGEMA_signal_15164 ;
    wire new_AGEMA_signal_15165 ;
    wire new_AGEMA_signal_15166 ;
    wire new_AGEMA_signal_15167 ;
    wire new_AGEMA_signal_15168 ;
    wire new_AGEMA_signal_15169 ;
    wire new_AGEMA_signal_15170 ;
    wire new_AGEMA_signal_15171 ;
    wire new_AGEMA_signal_15172 ;
    wire new_AGEMA_signal_15173 ;
    wire new_AGEMA_signal_15178 ;
    wire new_AGEMA_signal_15179 ;
    wire new_AGEMA_signal_15184 ;
    wire new_AGEMA_signal_15185 ;
    wire new_AGEMA_signal_15186 ;
    wire new_AGEMA_signal_15187 ;
    wire new_AGEMA_signal_15188 ;
    wire new_AGEMA_signal_15189 ;
    wire new_AGEMA_signal_15190 ;
    wire new_AGEMA_signal_15191 ;
    wire new_AGEMA_signal_15192 ;
    wire new_AGEMA_signal_15193 ;
    wire new_AGEMA_signal_15194 ;
    wire new_AGEMA_signal_15195 ;
    wire new_AGEMA_signal_15196 ;
    wire new_AGEMA_signal_15197 ;
    wire new_AGEMA_signal_15198 ;
    wire new_AGEMA_signal_15199 ;
    wire new_AGEMA_signal_15200 ;
    wire new_AGEMA_signal_15201 ;
    wire new_AGEMA_signal_15202 ;
    wire new_AGEMA_signal_15203 ;
    wire new_AGEMA_signal_15204 ;
    wire new_AGEMA_signal_15205 ;
    wire new_AGEMA_signal_15206 ;
    wire new_AGEMA_signal_15207 ;
    wire new_AGEMA_signal_15208 ;
    wire new_AGEMA_signal_15209 ;
    wire new_AGEMA_signal_15210 ;
    wire new_AGEMA_signal_15211 ;
    wire new_AGEMA_signal_15212 ;
    wire new_AGEMA_signal_15213 ;
    wire new_AGEMA_signal_15214 ;
    wire new_AGEMA_signal_15215 ;
    wire new_AGEMA_signal_15216 ;
    wire new_AGEMA_signal_15217 ;
    wire new_AGEMA_signal_15218 ;
    wire new_AGEMA_signal_15219 ;
    wire new_AGEMA_signal_15220 ;
    wire new_AGEMA_signal_15221 ;
    wire new_AGEMA_signal_15222 ;
    wire new_AGEMA_signal_15223 ;
    wire new_AGEMA_signal_15224 ;
    wire new_AGEMA_signal_15225 ;
    wire new_AGEMA_signal_15230 ;
    wire new_AGEMA_signal_15231 ;
    wire new_AGEMA_signal_15234 ;
    wire new_AGEMA_signal_15235 ;
    wire new_AGEMA_signal_15236 ;
    wire new_AGEMA_signal_15237 ;
    wire new_AGEMA_signal_15238 ;
    wire new_AGEMA_signal_15239 ;
    wire new_AGEMA_signal_15240 ;
    wire new_AGEMA_signal_15241 ;
    wire new_AGEMA_signal_15242 ;
    wire new_AGEMA_signal_15243 ;
    wire new_AGEMA_signal_15246 ;
    wire new_AGEMA_signal_15247 ;
    wire new_AGEMA_signal_15252 ;
    wire new_AGEMA_signal_15253 ;
    wire new_AGEMA_signal_15254 ;
    wire new_AGEMA_signal_15255 ;
    wire new_AGEMA_signal_15256 ;
    wire new_AGEMA_signal_15257 ;
    wire new_AGEMA_signal_15258 ;
    wire new_AGEMA_signal_15259 ;
    wire new_AGEMA_signal_15260 ;
    wire new_AGEMA_signal_15261 ;
    wire new_AGEMA_signal_15262 ;
    wire new_AGEMA_signal_15263 ;
    wire new_AGEMA_signal_15264 ;
    wire new_AGEMA_signal_15265 ;
    wire new_AGEMA_signal_15266 ;
    wire new_AGEMA_signal_15267 ;
    wire new_AGEMA_signal_15268 ;
    wire new_AGEMA_signal_15269 ;
    wire new_AGEMA_signal_15270 ;
    wire new_AGEMA_signal_15271 ;
    wire new_AGEMA_signal_15296 ;
    wire new_AGEMA_signal_15297 ;
    wire new_AGEMA_signal_15298 ;
    wire new_AGEMA_signal_15299 ;
    wire new_AGEMA_signal_15300 ;
    wire new_AGEMA_signal_15301 ;
    wire new_AGEMA_signal_15302 ;
    wire new_AGEMA_signal_15303 ;
    wire new_AGEMA_signal_15304 ;
    wire new_AGEMA_signal_15305 ;
    wire new_AGEMA_signal_15306 ;
    wire new_AGEMA_signal_15307 ;
    wire new_AGEMA_signal_15308 ;
    wire new_AGEMA_signal_15309 ;
    wire new_AGEMA_signal_15310 ;
    wire new_AGEMA_signal_15311 ;
    wire new_AGEMA_signal_15312 ;
    wire new_AGEMA_signal_15313 ;
    wire new_AGEMA_signal_15314 ;
    wire new_AGEMA_signal_15315 ;
    wire new_AGEMA_signal_15316 ;
    wire new_AGEMA_signal_15317 ;
    wire new_AGEMA_signal_15318 ;
    wire new_AGEMA_signal_15319 ;
    wire new_AGEMA_signal_15320 ;
    wire new_AGEMA_signal_15321 ;
    wire new_AGEMA_signal_15322 ;
    wire new_AGEMA_signal_15323 ;
    wire new_AGEMA_signal_15324 ;
    wire new_AGEMA_signal_15325 ;
    wire new_AGEMA_signal_15326 ;
    wire new_AGEMA_signal_15327 ;
    wire new_AGEMA_signal_15328 ;
    wire new_AGEMA_signal_15329 ;
    wire new_AGEMA_signal_15330 ;
    wire new_AGEMA_signal_15331 ;
    wire new_AGEMA_signal_15484 ;
    wire new_AGEMA_signal_15485 ;
    wire new_AGEMA_signal_15488 ;
    wire new_AGEMA_signal_15489 ;
    wire new_AGEMA_signal_15490 ;
    wire new_AGEMA_signal_15491 ;
    wire new_AGEMA_signal_15494 ;
    wire new_AGEMA_signal_15495 ;
    wire new_AGEMA_signal_15496 ;
    wire new_AGEMA_signal_15497 ;
    wire new_AGEMA_signal_15498 ;
    wire new_AGEMA_signal_15499 ;
    wire new_AGEMA_signal_15500 ;
    wire new_AGEMA_signal_15501 ;
    wire new_AGEMA_signal_15502 ;
    wire new_AGEMA_signal_15503 ;
    wire new_AGEMA_signal_15504 ;
    wire new_AGEMA_signal_15505 ;
    wire new_AGEMA_signal_15508 ;
    wire new_AGEMA_signal_15509 ;
    wire new_AGEMA_signal_15510 ;
    wire new_AGEMA_signal_15511 ;
    wire new_AGEMA_signal_15514 ;
    wire new_AGEMA_signal_15515 ;
    wire new_AGEMA_signal_15518 ;
    wire new_AGEMA_signal_15519 ;
    wire new_AGEMA_signal_15520 ;
    wire new_AGEMA_signal_15521 ;
    wire new_AGEMA_signal_15524 ;
    wire new_AGEMA_signal_15525 ;
    wire new_AGEMA_signal_15526 ;
    wire new_AGEMA_signal_15527 ;
    wire new_AGEMA_signal_15528 ;
    wire new_AGEMA_signal_15529 ;
    wire new_AGEMA_signal_15530 ;
    wire new_AGEMA_signal_15531 ;
    wire new_AGEMA_signal_15532 ;
    wire new_AGEMA_signal_15533 ;
    wire new_AGEMA_signal_15536 ;
    wire new_AGEMA_signal_15537 ;
    wire new_AGEMA_signal_15538 ;
    wire new_AGEMA_signal_15539 ;
    wire new_AGEMA_signal_15544 ;
    wire new_AGEMA_signal_15545 ;
    wire new_AGEMA_signal_15546 ;
    wire new_AGEMA_signal_15547 ;
    wire new_AGEMA_signal_15548 ;
    wire new_AGEMA_signal_15549 ;
    wire new_AGEMA_signal_15550 ;
    wire new_AGEMA_signal_15551 ;
    wire new_AGEMA_signal_15554 ;
    wire new_AGEMA_signal_15555 ;
    wire new_AGEMA_signal_15556 ;
    wire new_AGEMA_signal_15557 ;
    wire new_AGEMA_signal_15558 ;
    wire new_AGEMA_signal_15559 ;
    wire new_AGEMA_signal_15560 ;
    wire new_AGEMA_signal_15561 ;
    wire new_AGEMA_signal_15562 ;
    wire new_AGEMA_signal_15563 ;
    wire new_AGEMA_signal_15564 ;
    wire new_AGEMA_signal_15565 ;
    wire new_AGEMA_signal_15566 ;
    wire new_AGEMA_signal_15567 ;
    wire new_AGEMA_signal_15568 ;
    wire new_AGEMA_signal_15569 ;
    wire new_AGEMA_signal_15570 ;
    wire new_AGEMA_signal_15571 ;
    wire new_AGEMA_signal_15572 ;
    wire new_AGEMA_signal_15573 ;
    wire new_AGEMA_signal_15574 ;
    wire new_AGEMA_signal_15575 ;
    wire new_AGEMA_signal_15578 ;
    wire new_AGEMA_signal_15579 ;
    wire new_AGEMA_signal_15580 ;
    wire new_AGEMA_signal_15581 ;
    wire new_AGEMA_signal_15584 ;
    wire new_AGEMA_signal_15585 ;
    wire new_AGEMA_signal_15586 ;
    wire new_AGEMA_signal_15587 ;
    wire new_AGEMA_signal_15592 ;
    wire new_AGEMA_signal_15593 ;
    wire new_AGEMA_signal_15594 ;
    wire new_AGEMA_signal_15595 ;
    wire new_AGEMA_signal_15598 ;
    wire new_AGEMA_signal_15599 ;
    wire new_AGEMA_signal_15600 ;
    wire new_AGEMA_signal_15601 ;
    wire new_AGEMA_signal_15602 ;
    wire new_AGEMA_signal_15603 ;
    wire new_AGEMA_signal_15604 ;
    wire new_AGEMA_signal_15605 ;
    wire new_AGEMA_signal_15606 ;
    wire new_AGEMA_signal_15607 ;
    wire new_AGEMA_signal_15608 ;
    wire new_AGEMA_signal_15609 ;
    wire new_AGEMA_signal_15610 ;
    wire new_AGEMA_signal_15611 ;
    wire new_AGEMA_signal_15612 ;
    wire new_AGEMA_signal_15613 ;
    wire new_AGEMA_signal_15620 ;
    wire new_AGEMA_signal_15621 ;
    wire new_AGEMA_signal_15622 ;
    wire new_AGEMA_signal_15623 ;
    wire new_AGEMA_signal_15626 ;
    wire new_AGEMA_signal_15627 ;
    wire new_AGEMA_signal_15628 ;
    wire new_AGEMA_signal_15629 ;
    wire new_AGEMA_signal_15632 ;
    wire new_AGEMA_signal_15633 ;
    wire new_AGEMA_signal_15634 ;
    wire new_AGEMA_signal_15635 ;
    wire new_AGEMA_signal_15636 ;
    wire new_AGEMA_signal_15637 ;
    wire new_AGEMA_signal_15638 ;
    wire new_AGEMA_signal_15639 ;
    wire new_AGEMA_signal_15640 ;
    wire new_AGEMA_signal_15641 ;
    wire new_AGEMA_signal_15642 ;
    wire new_AGEMA_signal_15643 ;
    wire new_AGEMA_signal_15646 ;
    wire new_AGEMA_signal_15647 ;
    wire new_AGEMA_signal_15648 ;
    wire new_AGEMA_signal_15649 ;
    wire new_AGEMA_signal_15652 ;
    wire new_AGEMA_signal_15653 ;
    wire new_AGEMA_signal_15656 ;
    wire new_AGEMA_signal_15657 ;
    wire new_AGEMA_signal_15658 ;
    wire new_AGEMA_signal_15659 ;
    wire new_AGEMA_signal_15662 ;
    wire new_AGEMA_signal_15663 ;
    wire new_AGEMA_signal_15664 ;
    wire new_AGEMA_signal_15665 ;
    wire new_AGEMA_signal_15666 ;
    wire new_AGEMA_signal_15667 ;
    wire new_AGEMA_signal_15668 ;
    wire new_AGEMA_signal_15669 ;
    wire new_AGEMA_signal_15670 ;
    wire new_AGEMA_signal_15671 ;
    wire new_AGEMA_signal_15674 ;
    wire new_AGEMA_signal_15675 ;
    wire new_AGEMA_signal_15676 ;
    wire new_AGEMA_signal_15677 ;
    wire new_AGEMA_signal_15682 ;
    wire new_AGEMA_signal_15683 ;
    wire new_AGEMA_signal_15684 ;
    wire new_AGEMA_signal_15685 ;
    wire new_AGEMA_signal_15686 ;
    wire new_AGEMA_signal_15687 ;
    wire new_AGEMA_signal_15688 ;
    wire new_AGEMA_signal_15689 ;
    wire new_AGEMA_signal_15692 ;
    wire new_AGEMA_signal_15693 ;
    wire new_AGEMA_signal_15694 ;
    wire new_AGEMA_signal_15695 ;
    wire new_AGEMA_signal_15696 ;
    wire new_AGEMA_signal_15697 ;
    wire new_AGEMA_signal_15698 ;
    wire new_AGEMA_signal_15699 ;
    wire new_AGEMA_signal_15700 ;
    wire new_AGEMA_signal_15701 ;
    wire new_AGEMA_signal_15702 ;
    wire new_AGEMA_signal_15703 ;
    wire new_AGEMA_signal_15704 ;
    wire new_AGEMA_signal_15705 ;
    wire new_AGEMA_signal_15706 ;
    wire new_AGEMA_signal_15707 ;
    wire new_AGEMA_signal_15708 ;
    wire new_AGEMA_signal_15709 ;
    wire new_AGEMA_signal_15710 ;
    wire new_AGEMA_signal_15711 ;
    wire new_AGEMA_signal_15712 ;
    wire new_AGEMA_signal_15713 ;
    wire new_AGEMA_signal_15716 ;
    wire new_AGEMA_signal_15717 ;
    wire new_AGEMA_signal_15718 ;
    wire new_AGEMA_signal_15719 ;
    wire new_AGEMA_signal_15722 ;
    wire new_AGEMA_signal_15723 ;
    wire new_AGEMA_signal_15724 ;
    wire new_AGEMA_signal_15725 ;
    wire new_AGEMA_signal_15730 ;
    wire new_AGEMA_signal_15731 ;
    wire new_AGEMA_signal_15732 ;
    wire new_AGEMA_signal_15733 ;
    wire new_AGEMA_signal_15736 ;
    wire new_AGEMA_signal_15737 ;
    wire new_AGEMA_signal_15738 ;
    wire new_AGEMA_signal_15739 ;
    wire new_AGEMA_signal_15740 ;
    wire new_AGEMA_signal_15741 ;
    wire new_AGEMA_signal_15742 ;
    wire new_AGEMA_signal_15743 ;
    wire new_AGEMA_signal_15744 ;
    wire new_AGEMA_signal_15745 ;
    wire new_AGEMA_signal_15746 ;
    wire new_AGEMA_signal_15747 ;
    wire new_AGEMA_signal_15748 ;
    wire new_AGEMA_signal_15749 ;
    wire new_AGEMA_signal_15750 ;
    wire new_AGEMA_signal_15751 ;
    wire new_AGEMA_signal_15758 ;
    wire new_AGEMA_signal_15759 ;
    wire new_AGEMA_signal_15796 ;
    wire new_AGEMA_signal_15797 ;
    wire new_AGEMA_signal_15798 ;
    wire new_AGEMA_signal_15799 ;
    wire new_AGEMA_signal_15800 ;
    wire new_AGEMA_signal_15801 ;
    wire new_AGEMA_signal_15802 ;
    wire new_AGEMA_signal_15803 ;
    wire new_AGEMA_signal_15804 ;
    wire new_AGEMA_signal_15805 ;
    wire new_AGEMA_signal_15806 ;
    wire new_AGEMA_signal_15807 ;
    wire new_AGEMA_signal_15808 ;
    wire new_AGEMA_signal_15809 ;
    wire new_AGEMA_signal_15810 ;
    wire new_AGEMA_signal_15811 ;
    wire new_AGEMA_signal_15812 ;
    wire new_AGEMA_signal_15813 ;
    wire new_AGEMA_signal_15814 ;
    wire new_AGEMA_signal_15815 ;
    wire new_AGEMA_signal_15816 ;
    wire new_AGEMA_signal_15817 ;
    wire new_AGEMA_signal_15818 ;
    wire new_AGEMA_signal_15819 ;
    wire new_AGEMA_signal_15820 ;
    wire new_AGEMA_signal_15821 ;
    wire new_AGEMA_signal_15822 ;
    wire new_AGEMA_signal_15823 ;
    wire new_AGEMA_signal_15824 ;
    wire new_AGEMA_signal_15825 ;
    wire new_AGEMA_signal_15826 ;
    wire new_AGEMA_signal_15827 ;
    wire new_AGEMA_signal_15828 ;
    wire new_AGEMA_signal_15829 ;
    wire new_AGEMA_signal_15830 ;
    wire new_AGEMA_signal_15831 ;
    wire new_AGEMA_signal_15832 ;
    wire new_AGEMA_signal_15833 ;
    wire new_AGEMA_signal_15834 ;
    wire new_AGEMA_signal_15835 ;
    wire new_AGEMA_signal_15836 ;
    wire new_AGEMA_signal_15837 ;
    wire new_AGEMA_signal_15838 ;
    wire new_AGEMA_signal_15839 ;
    wire new_AGEMA_signal_15840 ;
    wire new_AGEMA_signal_15841 ;
    wire new_AGEMA_signal_15842 ;
    wire new_AGEMA_signal_15843 ;
    wire new_AGEMA_signal_15844 ;
    wire new_AGEMA_signal_15845 ;
    wire new_AGEMA_signal_15846 ;
    wire new_AGEMA_signal_15847 ;
    wire new_AGEMA_signal_15848 ;
    wire new_AGEMA_signal_15849 ;
    wire new_AGEMA_signal_15850 ;
    wire new_AGEMA_signal_15851 ;
    wire new_AGEMA_signal_15996 ;
    wire new_AGEMA_signal_15997 ;
    wire new_AGEMA_signal_16004 ;
    wire new_AGEMA_signal_16005 ;
    wire new_AGEMA_signal_16006 ;
    wire new_AGEMA_signal_16007 ;
    wire new_AGEMA_signal_16008 ;
    wire new_AGEMA_signal_16009 ;
    wire new_AGEMA_signal_16010 ;
    wire new_AGEMA_signal_16011 ;
    wire new_AGEMA_signal_16012 ;
    wire new_AGEMA_signal_16013 ;
    wire new_AGEMA_signal_16014 ;
    wire new_AGEMA_signal_16015 ;
    wire new_AGEMA_signal_16018 ;
    wire new_AGEMA_signal_16019 ;
    wire new_AGEMA_signal_16020 ;
    wire new_AGEMA_signal_16021 ;
    wire new_AGEMA_signal_16024 ;
    wire new_AGEMA_signal_16025 ;
    wire new_AGEMA_signal_16026 ;
    wire new_AGEMA_signal_16027 ;
    wire new_AGEMA_signal_16028 ;
    wire new_AGEMA_signal_16029 ;
    wire new_AGEMA_signal_16030 ;
    wire new_AGEMA_signal_16031 ;
    wire new_AGEMA_signal_16032 ;
    wire new_AGEMA_signal_16033 ;
    wire new_AGEMA_signal_16040 ;
    wire new_AGEMA_signal_16041 ;
    wire new_AGEMA_signal_16042 ;
    wire new_AGEMA_signal_16043 ;
    wire new_AGEMA_signal_16044 ;
    wire new_AGEMA_signal_16045 ;
    wire new_AGEMA_signal_16046 ;
    wire new_AGEMA_signal_16047 ;
    wire new_AGEMA_signal_16054 ;
    wire new_AGEMA_signal_16055 ;
    wire new_AGEMA_signal_16058 ;
    wire new_AGEMA_signal_16059 ;
    wire new_AGEMA_signal_16060 ;
    wire new_AGEMA_signal_16061 ;
    wire new_AGEMA_signal_16062 ;
    wire new_AGEMA_signal_16063 ;
    wire new_AGEMA_signal_16064 ;
    wire new_AGEMA_signal_16065 ;
    wire new_AGEMA_signal_16066 ;
    wire new_AGEMA_signal_16067 ;
    wire new_AGEMA_signal_16070 ;
    wire new_AGEMA_signal_16071 ;
    wire new_AGEMA_signal_16078 ;
    wire new_AGEMA_signal_16079 ;
    wire new_AGEMA_signal_16080 ;
    wire new_AGEMA_signal_16081 ;
    wire new_AGEMA_signal_16082 ;
    wire new_AGEMA_signal_16083 ;
    wire new_AGEMA_signal_16084 ;
    wire new_AGEMA_signal_16085 ;
    wire new_AGEMA_signal_16086 ;
    wire new_AGEMA_signal_16087 ;
    wire new_AGEMA_signal_16088 ;
    wire new_AGEMA_signal_16089 ;
    wire new_AGEMA_signal_16092 ;
    wire new_AGEMA_signal_16093 ;
    wire new_AGEMA_signal_16094 ;
    wire new_AGEMA_signal_16095 ;
    wire new_AGEMA_signal_16098 ;
    wire new_AGEMA_signal_16099 ;
    wire new_AGEMA_signal_16100 ;
    wire new_AGEMA_signal_16101 ;
    wire new_AGEMA_signal_16102 ;
    wire new_AGEMA_signal_16103 ;
    wire new_AGEMA_signal_16104 ;
    wire new_AGEMA_signal_16105 ;
    wire new_AGEMA_signal_16106 ;
    wire new_AGEMA_signal_16107 ;
    wire new_AGEMA_signal_16114 ;
    wire new_AGEMA_signal_16115 ;
    wire new_AGEMA_signal_16116 ;
    wire new_AGEMA_signal_16117 ;
    wire new_AGEMA_signal_16118 ;
    wire new_AGEMA_signal_16119 ;
    wire new_AGEMA_signal_16120 ;
    wire new_AGEMA_signal_16121 ;
    wire new_AGEMA_signal_16128 ;
    wire new_AGEMA_signal_16129 ;
    wire new_AGEMA_signal_16132 ;
    wire new_AGEMA_signal_16133 ;
    wire new_AGEMA_signal_16134 ;
    wire new_AGEMA_signal_16135 ;
    wire new_AGEMA_signal_16136 ;
    wire new_AGEMA_signal_16137 ;
    wire new_AGEMA_signal_16138 ;
    wire new_AGEMA_signal_16139 ;
    wire new_AGEMA_signal_16140 ;
    wire new_AGEMA_signal_16141 ;
    wire new_AGEMA_signal_16180 ;
    wire new_AGEMA_signal_16181 ;
    wire new_AGEMA_signal_16182 ;
    wire new_AGEMA_signal_16183 ;
    wire new_AGEMA_signal_16184 ;
    wire new_AGEMA_signal_16185 ;
    wire new_AGEMA_signal_16186 ;
    wire new_AGEMA_signal_16187 ;
    wire new_AGEMA_signal_16188 ;
    wire new_AGEMA_signal_16189 ;
    wire new_AGEMA_signal_16190 ;
    wire new_AGEMA_signal_16191 ;
    wire new_AGEMA_signal_16192 ;
    wire new_AGEMA_signal_16193 ;
    wire new_AGEMA_signal_16194 ;
    wire new_AGEMA_signal_16195 ;
    wire new_AGEMA_signal_16196 ;
    wire new_AGEMA_signal_16197 ;
    wire new_AGEMA_signal_16198 ;
    wire new_AGEMA_signal_16199 ;
    wire new_AGEMA_signal_16200 ;
    wire new_AGEMA_signal_16201 ;
    wire new_AGEMA_signal_16202 ;
    wire new_AGEMA_signal_16203 ;
    wire new_AGEMA_signal_16204 ;
    wire new_AGEMA_signal_16205 ;
    wire new_AGEMA_signal_16206 ;
    wire new_AGEMA_signal_16207 ;
    wire new_AGEMA_signal_16208 ;
    wire new_AGEMA_signal_16209 ;
    wire new_AGEMA_signal_16210 ;
    wire new_AGEMA_signal_16211 ;
    wire new_AGEMA_signal_16212 ;
    wire new_AGEMA_signal_16213 ;
    wire new_AGEMA_signal_16214 ;
    wire new_AGEMA_signal_16215 ;
    wire new_AGEMA_signal_16216 ;
    wire new_AGEMA_signal_16217 ;
    wire new_AGEMA_signal_16218 ;
    wire new_AGEMA_signal_16219 ;
    wire new_AGEMA_signal_16220 ;
    wire new_AGEMA_signal_16221 ;
    wire new_AGEMA_signal_16222 ;
    wire new_AGEMA_signal_16223 ;
    wire new_AGEMA_signal_16224 ;
    wire new_AGEMA_signal_16225 ;
    wire new_AGEMA_signal_16226 ;
    wire new_AGEMA_signal_16227 ;
    wire new_AGEMA_signal_16228 ;
    wire new_AGEMA_signal_16229 ;
    wire new_AGEMA_signal_16230 ;
    wire new_AGEMA_signal_16231 ;
    wire new_AGEMA_signal_16232 ;
    wire new_AGEMA_signal_16233 ;
    wire new_AGEMA_signal_16234 ;
    wire new_AGEMA_signal_16235 ;
    wire new_AGEMA_signal_16236 ;
    wire new_AGEMA_signal_16237 ;
    wire new_AGEMA_signal_16238 ;
    wire new_AGEMA_signal_16239 ;
    wire new_AGEMA_signal_16240 ;
    wire new_AGEMA_signal_16241 ;
    wire new_AGEMA_signal_16242 ;
    wire new_AGEMA_signal_16243 ;
    wire new_AGEMA_signal_16244 ;
    wire new_AGEMA_signal_16245 ;
    wire new_AGEMA_signal_16246 ;
    wire new_AGEMA_signal_16247 ;
    wire new_AGEMA_signal_16248 ;
    wire new_AGEMA_signal_16249 ;
    wire new_AGEMA_signal_16250 ;
    wire new_AGEMA_signal_16251 ;
    wire new_AGEMA_signal_16362 ;
    wire new_AGEMA_signal_16363 ;
    wire new_AGEMA_signal_16364 ;
    wire new_AGEMA_signal_16365 ;
    wire new_AGEMA_signal_16366 ;
    wire new_AGEMA_signal_16367 ;
    wire new_AGEMA_signal_16374 ;
    wire new_AGEMA_signal_16375 ;
    wire new_AGEMA_signal_16376 ;
    wire new_AGEMA_signal_16377 ;
    wire new_AGEMA_signal_16378 ;
    wire new_AGEMA_signal_16379 ;
    wire new_AGEMA_signal_16436 ;
    wire new_AGEMA_signal_16437 ;
    wire new_AGEMA_signal_16438 ;
    wire new_AGEMA_signal_16439 ;
    wire new_AGEMA_signal_16464 ;
    wire new_AGEMA_signal_16465 ;
    wire new_AGEMA_signal_16468 ;
    wire new_AGEMA_signal_16469 ;
    wire new_AGEMA_signal_16544 ;
    wire new_AGEMA_signal_16545 ;
    wire new_AGEMA_signal_16546 ;
    wire new_AGEMA_signal_16547 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_0_U1 ( .s (p256_sel), .b ({w0_s2[0], w0_s1[0], w0_s0[0]}), .a ({w1_s2[0], w1_s1[0], w1_s0[0]}), .c ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, addc_in[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_1_U1 ( .s (p256_sel), .b ({w0_s2[1], w0_s1[1], w0_s0[1]}), .a ({w1_s2[1], w1_s1[1], w1_s0[1]}), .c ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, addc_in[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_2_U1 ( .s (p256_sel), .b ({w0_s2[2], w0_s1[2], w0_s0[2]}), .a ({w1_s2[2], w1_s1[2], w1_s0[2]}), .c ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, addc_in[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_3_U1 ( .s (p256_sel), .b ({w0_s2[3], w0_s1[3], w0_s0[3]}), .a ({w1_s2[3], w1_s1[3], w1_s0[3]}), .c ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, addc_in[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_4_U1 ( .s (p256_sel), .b ({w0_s2[4], w0_s1[4], w0_s0[4]}), .a ({w1_s2[4], w1_s1[4], w1_s0[4]}), .c ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, addc_in[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_5_U1 ( .s (p256_sel), .b ({w0_s2[5], w0_s1[5], w0_s0[5]}), .a ({w1_s2[5], w1_s1[5], w1_s0[5]}), .c ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, addc_in[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_6_U1 ( .s (p256_sel), .b ({w0_s2[6], w0_s1[6], w0_s0[6]}), .a ({w1_s2[6], w1_s1[6], w1_s0[6]}), .c ({new_AGEMA_signal_5773, new_AGEMA_signal_5772, addc_in[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_7_U1 ( .s (p256_sel), .b ({w0_s2[7], w0_s1[7], w0_s0[7]}), .a ({w1_s2[7], w1_s1[7], w1_s0[7]}), .c ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, addc_in[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_8_U1 ( .s (p256_sel), .b ({w0_s2[8], w0_s1[8], w0_s0[8]}), .a ({w1_s2[8], w1_s1[8], w1_s0[8]}), .c ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, addc_in[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_9_U1 ( .s (p256_sel), .b ({w0_s2[9], w0_s1[9], w0_s0[9]}), .a ({w1_s2[9], w1_s1[9], w1_s0[9]}), .c ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, addc_in[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_10_U1 ( .s (p256_sel), .b ({w0_s2[10], w0_s1[10], w0_s0[10]}), .a ({w1_s2[10], w1_s1[10], w1_s0[10]}), .c ({new_AGEMA_signal_5797, new_AGEMA_signal_5796, addc_in[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_11_U1 ( .s (p256_sel), .b ({w0_s2[11], w0_s1[11], w0_s0[11]}), .a ({w1_s2[11], w1_s1[11], w1_s0[11]}), .c ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, addc_in[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_12_U1 ( .s (p256_sel), .b ({w0_s2[12], w0_s1[12], w0_s0[12]}), .a ({w1_s2[12], w1_s1[12], w1_s0[12]}), .c ({new_AGEMA_signal_5809, new_AGEMA_signal_5808, addc_in[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_13_U1 ( .s (p256_sel), .b ({w0_s2[13], w0_s1[13], w0_s0[13]}), .a ({w1_s2[13], w1_s1[13], w1_s0[13]}), .c ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, addc_in[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_14_U1 ( .s (p256_sel), .b ({w0_s2[14], w0_s1[14], w0_s0[14]}), .a ({w1_s2[14], w1_s1[14], w1_s0[14]}), .c ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, addc_in[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_15_U1 ( .s (p256_sel), .b ({w0_s2[15], w0_s1[15], w0_s0[15]}), .a ({w1_s2[15], w1_s1[15], w1_s0[15]}), .c ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, addc_in[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_16_U1 ( .s (p256_sel), .b ({w0_s2[16], w0_s1[16], w0_s0[16]}), .a ({w1_s2[16], w1_s1[16], w1_s0[16]}), .c ({new_AGEMA_signal_5833, new_AGEMA_signal_5832, addc_in[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_17_U1 ( .s (p256_sel), .b ({w0_s2[17], w0_s1[17], w0_s0[17]}), .a ({w1_s2[17], w1_s1[17], w1_s0[17]}), .c ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, addc_in[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_18_U1 ( .s (p256_sel), .b ({w0_s2[18], w0_s1[18], w0_s0[18]}), .a ({w1_s2[18], w1_s1[18], w1_s0[18]}), .c ({new_AGEMA_signal_5845, new_AGEMA_signal_5844, addc_in[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_19_U1 ( .s (p256_sel), .b ({w0_s2[19], w0_s1[19], w0_s0[19]}), .a ({w1_s2[19], w1_s1[19], w1_s0[19]}), .c ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, addc_in[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_20_U1 ( .s (p256_sel), .b ({w0_s2[20], w0_s1[20], w0_s0[20]}), .a ({w1_s2[20], w1_s1[20], w1_s0[20]}), .c ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, addc_in[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_21_U1 ( .s (p256_sel), .b ({w0_s2[21], w0_s1[21], w0_s0[21]}), .a ({w1_s2[21], w1_s1[21], w1_s0[21]}), .c ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, addc_in[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_22_U1 ( .s (p256_sel), .b ({w0_s2[22], w0_s1[22], w0_s0[22]}), .a ({w1_s2[22], w1_s1[22], w1_s0[22]}), .c ({new_AGEMA_signal_5869, new_AGEMA_signal_5868, addc_in[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_23_U1 ( .s (p256_sel), .b ({w0_s2[23], w0_s1[23], w0_s0[23]}), .a ({w1_s2[23], w1_s1[23], w1_s0[23]}), .c ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, addc_in[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_24_U1 ( .s (p256_sel), .b ({w0_s2[24], w0_s1[24], w0_s0[24]}), .a ({w1_s2[24], w1_s1[24], w1_s0[24]}), .c ({new_AGEMA_signal_5881, new_AGEMA_signal_5880, addc_in[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_25_U1 ( .s (p256_sel), .b ({w0_s2[25], w0_s1[25], w0_s0[25]}), .a ({w1_s2[25], w1_s1[25], w1_s0[25]}), .c ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, addc_in[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_26_U1 ( .s (p256_sel), .b ({w0_s2[26], w0_s1[26], w0_s0[26]}), .a ({w1_s2[26], w1_s1[26], w1_s0[26]}), .c ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, addc_in[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_27_U1 ( .s (p256_sel), .b ({w0_s2[27], w0_s1[27], w0_s0[27]}), .a ({w1_s2[27], w1_s1[27], w1_s0[27]}), .c ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, addc_in[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_28_U1 ( .s (p256_sel), .b ({w0_s2[28], w0_s1[28], w0_s0[28]}), .a ({w1_s2[28], w1_s1[28], w1_s0[28]}), .c ({new_AGEMA_signal_5905, new_AGEMA_signal_5904, addc_in[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_29_U1 ( .s (p256_sel), .b ({w0_s2[29], w0_s1[29], w0_s0[29]}), .a ({w1_s2[29], w1_s1[29], w1_s0[29]}), .c ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, addc_in[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_30_U1 ( .s (p256_sel), .b ({w0_s2[30], w0_s1[30], w0_s0[30]}), .a ({w1_s2[30], w1_s1[30], w1_s0[30]}), .c ({new_AGEMA_signal_5917, new_AGEMA_signal_5916, addc_in[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_31_U1 ( .s (p256_sel), .b ({w0_s2[31], w0_s1[31], w0_s0[31]}), .a ({w1_s2[31], w1_s1[31], w1_s0[31]}), .c ({new_AGEMA_signal_5923, new_AGEMA_signal_5922, addc_in[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_32_U1 ( .s (p256_sel), .b ({w0_s2[32], w0_s1[32], w0_s0[32]}), .a ({w1_s2[32], w1_s1[32], w1_s0[32]}), .c ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, addc_in[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_33_U1 ( .s (p256_sel), .b ({w0_s2[33], w0_s1[33], w0_s0[33]}), .a ({w1_s2[33], w1_s1[33], w1_s0[33]}), .c ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, addc_in[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_34_U1 ( .s (p256_sel), .b ({w0_s2[34], w0_s1[34], w0_s0[34]}), .a ({w1_s2[34], w1_s1[34], w1_s0[34]}), .c ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, addc_in[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_35_U1 ( .s (p256_sel), .b ({w0_s2[35], w0_s1[35], w0_s0[35]}), .a ({w1_s2[35], w1_s1[35], w1_s0[35]}), .c ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, addc_in[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_36_U1 ( .s (p256_sel), .b ({w0_s2[36], w0_s1[36], w0_s0[36]}), .a ({w1_s2[36], w1_s1[36], w1_s0[36]}), .c ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, addc_in[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_37_U1 ( .s (p256_sel), .b ({w0_s2[37], w0_s1[37], w0_s0[37]}), .a ({w1_s2[37], w1_s1[37], w1_s0[37]}), .c ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, addc_in[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_38_U1 ( .s (p256_sel), .b ({w0_s2[38], w0_s1[38], w0_s0[38]}), .a ({w1_s2[38], w1_s1[38], w1_s0[38]}), .c ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, addc_in[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_39_U1 ( .s (p256_sel), .b ({w0_s2[39], w0_s1[39], w0_s0[39]}), .a ({w1_s2[39], w1_s1[39], w1_s0[39]}), .c ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, addc_in[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_40_U1 ( .s (p256_sel), .b ({w0_s2[40], w0_s1[40], w0_s0[40]}), .a ({w1_s2[40], w1_s1[40], w1_s0[40]}), .c ({new_AGEMA_signal_5977, new_AGEMA_signal_5976, addc_in[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_41_U1 ( .s (p256_sel), .b ({w0_s2[41], w0_s1[41], w0_s0[41]}), .a ({w1_s2[41], w1_s1[41], w1_s0[41]}), .c ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, addc_in[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_42_U1 ( .s (p256_sel), .b ({w0_s2[42], w0_s1[42], w0_s0[42]}), .a ({w1_s2[42], w1_s1[42], w1_s0[42]}), .c ({new_AGEMA_signal_5989, new_AGEMA_signal_5988, addc_in[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_43_U1 ( .s (p256_sel), .b ({w0_s2[43], w0_s1[43], w0_s0[43]}), .a ({w1_s2[43], w1_s1[43], w1_s0[43]}), .c ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, addc_in[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_44_U1 ( .s (p256_sel), .b ({w0_s2[44], w0_s1[44], w0_s0[44]}), .a ({w1_s2[44], w1_s1[44], w1_s0[44]}), .c ({new_AGEMA_signal_6001, new_AGEMA_signal_6000, addc_in[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_45_U1 ( .s (p256_sel), .b ({w0_s2[45], w0_s1[45], w0_s0[45]}), .a ({w1_s2[45], w1_s1[45], w1_s0[45]}), .c ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, addc_in[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_46_U1 ( .s (p256_sel), .b ({w0_s2[46], w0_s1[46], w0_s0[46]}), .a ({w1_s2[46], w1_s1[46], w1_s0[46]}), .c ({new_AGEMA_signal_6013, new_AGEMA_signal_6012, addc_in[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_47_U1 ( .s (p256_sel), .b ({w0_s2[47], w0_s1[47], w0_s0[47]}), .a ({w1_s2[47], w1_s1[47], w1_s0[47]}), .c ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, addc_in[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_48_U1 ( .s (p256_sel), .b ({w0_s2[48], w0_s1[48], w0_s0[48]}), .a ({w1_s2[48], w1_s1[48], w1_s0[48]}), .c ({new_AGEMA_signal_6025, new_AGEMA_signal_6024, addc_in[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_49_U1 ( .s (p256_sel), .b ({w0_s2[49], w0_s1[49], w0_s0[49]}), .a ({w1_s2[49], w1_s1[49], w1_s0[49]}), .c ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, addc_in[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_50_U1 ( .s (p256_sel), .b ({w0_s2[50], w0_s1[50], w0_s0[50]}), .a ({w1_s2[50], w1_s1[50], w1_s0[50]}), .c ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, addc_in[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_51_U1 ( .s (p256_sel), .b ({w0_s2[51], w0_s1[51], w0_s0[51]}), .a ({w1_s2[51], w1_s1[51], w1_s0[51]}), .c ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, addc_in[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_52_U1 ( .s (p256_sel), .b ({w0_s2[52], w0_s1[52], w0_s0[52]}), .a ({w1_s2[52], w1_s1[52], w1_s0[52]}), .c ({new_AGEMA_signal_6049, new_AGEMA_signal_6048, addc_in[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_53_U1 ( .s (p256_sel), .b ({w0_s2[53], w0_s1[53], w0_s0[53]}), .a ({w1_s2[53], w1_s1[53], w1_s0[53]}), .c ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, addc_in[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_54_U1 ( .s (p256_sel), .b ({w0_s2[54], w0_s1[54], w0_s0[54]}), .a ({w1_s2[54], w1_s1[54], w1_s0[54]}), .c ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, addc_in[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_55_U1 ( .s (p256_sel), .b ({w0_s2[55], w0_s1[55], w0_s0[55]}), .a ({w1_s2[55], w1_s1[55], w1_s0[55]}), .c ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, addc_in[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_56_U1 ( .s (p256_sel), .b ({w0_s2[56], w0_s1[56], w0_s0[56]}), .a ({w1_s2[56], w1_s1[56], w1_s0[56]}), .c ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, addc_in[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_57_U1 ( .s (p256_sel), .b ({w0_s2[57], w0_s1[57], w0_s0[57]}), .a ({w1_s2[57], w1_s1[57], w1_s0[57]}), .c ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, addc_in[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_58_U1 ( .s (p256_sel), .b ({w0_s2[58], w0_s1[58], w0_s0[58]}), .a ({w1_s2[58], w1_s1[58], w1_s0[58]}), .c ({new_AGEMA_signal_6085, new_AGEMA_signal_6084, addc_in[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_59_U1 ( .s (p256_sel), .b ({w0_s2[59], w0_s1[59], w0_s0[59]}), .a ({w1_s2[59], w1_s1[59], w1_s0[59]}), .c ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, addc_in[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_60_U1 ( .s (p256_sel), .b ({w0_s2[60], w0_s1[60], w0_s0[60]}), .a ({w1_s2[60], w1_s1[60], w1_s0[60]}), .c ({new_AGEMA_signal_6097, new_AGEMA_signal_6096, addc_in[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_61_U1 ( .s (p256_sel), .b ({w0_s2[61], w0_s1[61], w0_s0[61]}), .a ({w1_s2[61], w1_s1[61], w1_s0[61]}), .c ({new_AGEMA_signal_6103, new_AGEMA_signal_6102, addc_in[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_62_U1 ( .s (p256_sel), .b ({w0_s2[62], w0_s1[62], w0_s0[62]}), .a ({w1_s2[62], w1_s1[62], w1_s0[62]}), .c ({new_AGEMA_signal_6109, new_AGEMA_signal_6108, addc_in[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_63_U1 ( .s (p256_sel), .b ({w0_s2[63], w0_s1[63], w0_s0[63]}), .a ({w1_s2[63], w1_s1[63], w1_s0[63]}), .c ({new_AGEMA_signal_6115, new_AGEMA_signal_6114, addc_in[63]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_64_U1 ( .s (p256_sel), .b ({w0_s2[64], w0_s1[64], w0_s0[64]}), .a ({w1_s2[64], w1_s1[64], w1_s0[64]}), .c ({new_AGEMA_signal_6121, new_AGEMA_signal_6120, addc_in[64]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_65_U1 ( .s (p256_sel), .b ({w0_s2[65], w0_s1[65], w0_s0[65]}), .a ({w1_s2[65], w1_s1[65], w1_s0[65]}), .c ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, addc_in[65]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_66_U1 ( .s (p256_sel), .b ({w0_s2[66], w0_s1[66], w0_s0[66]}), .a ({w1_s2[66], w1_s1[66], w1_s0[66]}), .c ({new_AGEMA_signal_6133, new_AGEMA_signal_6132, addc_in[66]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_67_U1 ( .s (p256_sel), .b ({w0_s2[67], w0_s1[67], w0_s0[67]}), .a ({w1_s2[67], w1_s1[67], w1_s0[67]}), .c ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, addc_in[67]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_68_U1 ( .s (p256_sel), .b ({w0_s2[68], w0_s1[68], w0_s0[68]}), .a ({w1_s2[68], w1_s1[68], w1_s0[68]}), .c ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, addc_in[68]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_69_U1 ( .s (p256_sel), .b ({w0_s2[69], w0_s1[69], w0_s0[69]}), .a ({w1_s2[69], w1_s1[69], w1_s0[69]}), .c ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, addc_in[69]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_70_U1 ( .s (p256_sel), .b ({w0_s2[70], w0_s1[70], w0_s0[70]}), .a ({w1_s2[70], w1_s1[70], w1_s0[70]}), .c ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, addc_in[70]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_71_U1 ( .s (p256_sel), .b ({w0_s2[71], w0_s1[71], w0_s0[71]}), .a ({w1_s2[71], w1_s1[71], w1_s0[71]}), .c ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, addc_in[71]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_72_U1 ( .s (p256_sel), .b ({w0_s2[72], w0_s1[72], w0_s0[72]}), .a ({w1_s2[72], w1_s1[72], w1_s0[72]}), .c ({new_AGEMA_signal_6169, new_AGEMA_signal_6168, addc_in[72]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_73_U1 ( .s (p256_sel), .b ({w0_s2[73], w0_s1[73], w0_s0[73]}), .a ({w1_s2[73], w1_s1[73], w1_s0[73]}), .c ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, addc_in[73]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_74_U1 ( .s (p256_sel), .b ({w0_s2[74], w0_s1[74], w0_s0[74]}), .a ({w1_s2[74], w1_s1[74], w1_s0[74]}), .c ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, addc_in[74]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_75_U1 ( .s (p256_sel), .b ({w0_s2[75], w0_s1[75], w0_s0[75]}), .a ({w1_s2[75], w1_s1[75], w1_s0[75]}), .c ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, addc_in[75]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_76_U1 ( .s (p256_sel), .b ({w0_s2[76], w0_s1[76], w0_s0[76]}), .a ({w1_s2[76], w1_s1[76], w1_s0[76]}), .c ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, addc_in[76]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_77_U1 ( .s (p256_sel), .b ({w0_s2[77], w0_s1[77], w0_s0[77]}), .a ({w1_s2[77], w1_s1[77], w1_s0[77]}), .c ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, addc_in[77]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_78_U1 ( .s (p256_sel), .b ({w0_s2[78], w0_s1[78], w0_s0[78]}), .a ({w1_s2[78], w1_s1[78], w1_s0[78]}), .c ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, addc_in[78]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_79_U1 ( .s (p256_sel), .b ({w0_s2[79], w0_s1[79], w0_s0[79]}), .a ({w1_s2[79], w1_s1[79], w1_s0[79]}), .c ({new_AGEMA_signal_6211, new_AGEMA_signal_6210, addc_in[79]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_80_U1 ( .s (p256_sel), .b ({w0_s2[80], w0_s1[80], w0_s0[80]}), .a ({w1_s2[80], w1_s1[80], w1_s0[80]}), .c ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, addc_in[80]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_81_U1 ( .s (p256_sel), .b ({w0_s2[81], w0_s1[81], w0_s0[81]}), .a ({w1_s2[81], w1_s1[81], w1_s0[81]}), .c ({new_AGEMA_signal_6223, new_AGEMA_signal_6222, addc_in[81]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_82_U1 ( .s (p256_sel), .b ({w0_s2[82], w0_s1[82], w0_s0[82]}), .a ({w1_s2[82], w1_s1[82], w1_s0[82]}), .c ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, addc_in[82]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_83_U1 ( .s (p256_sel), .b ({w0_s2[83], w0_s1[83], w0_s0[83]}), .a ({w1_s2[83], w1_s1[83], w1_s0[83]}), .c ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, addc_in[83]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_84_U1 ( .s (p256_sel), .b ({w0_s2[84], w0_s1[84], w0_s0[84]}), .a ({w1_s2[84], w1_s1[84], w1_s0[84]}), .c ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, addc_in[84]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_85_U1 ( .s (p256_sel), .b ({w0_s2[85], w0_s1[85], w0_s0[85]}), .a ({w1_s2[85], w1_s1[85], w1_s0[85]}), .c ({new_AGEMA_signal_6247, new_AGEMA_signal_6246, addc_in[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_86_U1 ( .s (p256_sel), .b ({w0_s2[86], w0_s1[86], w0_s0[86]}), .a ({w1_s2[86], w1_s1[86], w1_s0[86]}), .c ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, addc_in[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_87_U1 ( .s (p256_sel), .b ({w0_s2[87], w0_s1[87], w0_s0[87]}), .a ({w1_s2[87], w1_s1[87], w1_s0[87]}), .c ({new_AGEMA_signal_6259, new_AGEMA_signal_6258, addc_in[87]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_88_U1 ( .s (p256_sel), .b ({w0_s2[88], w0_s1[88], w0_s0[88]}), .a ({w1_s2[88], w1_s1[88], w1_s0[88]}), .c ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, addc_in[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_89_U1 ( .s (p256_sel), .b ({w0_s2[89], w0_s1[89], w0_s0[89]}), .a ({w1_s2[89], w1_s1[89], w1_s0[89]}), .c ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, addc_in[89]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_90_U1 ( .s (p256_sel), .b ({w0_s2[90], w0_s1[90], w0_s0[90]}), .a ({w1_s2[90], w1_s1[90], w1_s0[90]}), .c ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, addc_in[90]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_91_U1 ( .s (p256_sel), .b ({w0_s2[91], w0_s1[91], w0_s0[91]}), .a ({w1_s2[91], w1_s1[91], w1_s0[91]}), .c ({new_AGEMA_signal_6283, new_AGEMA_signal_6282, addc_in[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_92_U1 ( .s (p256_sel), .b ({w0_s2[92], w0_s1[92], w0_s0[92]}), .a ({w1_s2[92], w1_s1[92], w1_s0[92]}), .c ({new_AGEMA_signal_6289, new_AGEMA_signal_6288, addc_in[92]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_93_U1 ( .s (p256_sel), .b ({w0_s2[93], w0_s1[93], w0_s0[93]}), .a ({w1_s2[93], w1_s1[93], w1_s0[93]}), .c ({new_AGEMA_signal_6295, new_AGEMA_signal_6294, addc_in[93]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_94_U1 ( .s (p256_sel), .b ({w0_s2[94], w0_s1[94], w0_s0[94]}), .a ({w1_s2[94], w1_s1[94], w1_s0[94]}), .c ({new_AGEMA_signal_6301, new_AGEMA_signal_6300, addc_in[94]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_95_U1 ( .s (p256_sel), .b ({w0_s2[95], w0_s1[95], w0_s0[95]}), .a ({w1_s2[95], w1_s1[95], w1_s0[95]}), .c ({new_AGEMA_signal_6307, new_AGEMA_signal_6306, addc_in[95]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_96_U1 ( .s (p256_sel), .b ({w0_s2[96], w0_s1[96], w0_s0[96]}), .a ({w1_s2[96], w1_s1[96], w1_s0[96]}), .c ({new_AGEMA_signal_6313, new_AGEMA_signal_6312, addc_in[96]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_97_U1 ( .s (p256_sel), .b ({w0_s2[97], w0_s1[97], w0_s0[97]}), .a ({w1_s2[97], w1_s1[97], w1_s0[97]}), .c ({new_AGEMA_signal_6319, new_AGEMA_signal_6318, addc_in[97]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_98_U1 ( .s (p256_sel), .b ({w0_s2[98], w0_s1[98], w0_s0[98]}), .a ({w1_s2[98], w1_s1[98], w1_s0[98]}), .c ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, addc_in[98]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_99_U1 ( .s (p256_sel), .b ({w0_s2[99], w0_s1[99], w0_s0[99]}), .a ({w1_s2[99], w1_s1[99], w1_s0[99]}), .c ({new_AGEMA_signal_6331, new_AGEMA_signal_6330, addc_in[99]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_100_U1 ( .s (p256_sel), .b ({w0_s2[100], w0_s1[100], w0_s0[100]}), .a ({w1_s2[100], w1_s1[100], w1_s0[100]}), .c ({new_AGEMA_signal_6337, new_AGEMA_signal_6336, addc_in[100]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_101_U1 ( .s (p256_sel), .b ({w0_s2[101], w0_s1[101], w0_s0[101]}), .a ({w1_s2[101], w1_s1[101], w1_s0[101]}), .c ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, addc_in[101]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_102_U1 ( .s (p256_sel), .b ({w0_s2[102], w0_s1[102], w0_s0[102]}), .a ({w1_s2[102], w1_s1[102], w1_s0[102]}), .c ({new_AGEMA_signal_6349, new_AGEMA_signal_6348, addc_in[102]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_103_U1 ( .s (p256_sel), .b ({w0_s2[103], w0_s1[103], w0_s0[103]}), .a ({w1_s2[103], w1_s1[103], w1_s0[103]}), .c ({new_AGEMA_signal_6355, new_AGEMA_signal_6354, addc_in[103]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_104_U1 ( .s (p256_sel), .b ({w0_s2[104], w0_s1[104], w0_s0[104]}), .a ({w1_s2[104], w1_s1[104], w1_s0[104]}), .c ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, addc_in[104]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_105_U1 ( .s (p256_sel), .b ({w0_s2[105], w0_s1[105], w0_s0[105]}), .a ({w1_s2[105], w1_s1[105], w1_s0[105]}), .c ({new_AGEMA_signal_6367, new_AGEMA_signal_6366, addc_in[105]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_106_U1 ( .s (p256_sel), .b ({w0_s2[106], w0_s1[106], w0_s0[106]}), .a ({w1_s2[106], w1_s1[106], w1_s0[106]}), .c ({new_AGEMA_signal_6373, new_AGEMA_signal_6372, addc_in[106]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_107_U1 ( .s (p256_sel), .b ({w0_s2[107], w0_s1[107], w0_s0[107]}), .a ({w1_s2[107], w1_s1[107], w1_s0[107]}), .c ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, addc_in[107]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_108_U1 ( .s (p256_sel), .b ({w0_s2[108], w0_s1[108], w0_s0[108]}), .a ({w1_s2[108], w1_s1[108], w1_s0[108]}), .c ({new_AGEMA_signal_6385, new_AGEMA_signal_6384, addc_in[108]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_109_U1 ( .s (p256_sel), .b ({w0_s2[109], w0_s1[109], w0_s0[109]}), .a ({w1_s2[109], w1_s1[109], w1_s0[109]}), .c ({new_AGEMA_signal_6391, new_AGEMA_signal_6390, addc_in[109]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_110_U1 ( .s (p256_sel), .b ({w0_s2[110], w0_s1[110], w0_s0[110]}), .a ({w1_s2[110], w1_s1[110], w1_s0[110]}), .c ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, addc_in[110]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_111_U1 ( .s (p256_sel), .b ({w0_s2[111], w0_s1[111], w0_s0[111]}), .a ({w1_s2[111], w1_s1[111], w1_s0[111]}), .c ({new_AGEMA_signal_6403, new_AGEMA_signal_6402, addc_in[111]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_112_U1 ( .s (p256_sel), .b ({w0_s2[112], w0_s1[112], w0_s0[112]}), .a ({w1_s2[112], w1_s1[112], w1_s0[112]}), .c ({new_AGEMA_signal_6409, new_AGEMA_signal_6408, addc_in[112]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_113_U1 ( .s (p256_sel), .b ({w0_s2[113], w0_s1[113], w0_s0[113]}), .a ({w1_s2[113], w1_s1[113], w1_s0[113]}), .c ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, addc_in[113]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_114_U1 ( .s (p256_sel), .b ({w0_s2[114], w0_s1[114], w0_s0[114]}), .a ({w1_s2[114], w1_s1[114], w1_s0[114]}), .c ({new_AGEMA_signal_6421, new_AGEMA_signal_6420, addc_in[114]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_115_U1 ( .s (p256_sel), .b ({w0_s2[115], w0_s1[115], w0_s0[115]}), .a ({w1_s2[115], w1_s1[115], w1_s0[115]}), .c ({new_AGEMA_signal_6427, new_AGEMA_signal_6426, addc_in[115]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_116_U1 ( .s (p256_sel), .b ({w0_s2[116], w0_s1[116], w0_s0[116]}), .a ({w1_s2[116], w1_s1[116], w1_s0[116]}), .c ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, addc_in[116]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_117_U1 ( .s (p256_sel), .b ({w0_s2[117], w0_s1[117], w0_s0[117]}), .a ({w1_s2[117], w1_s1[117], w1_s0[117]}), .c ({new_AGEMA_signal_6439, new_AGEMA_signal_6438, addc_in[117]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_118_U1 ( .s (p256_sel), .b ({w0_s2[118], w0_s1[118], w0_s0[118]}), .a ({w1_s2[118], w1_s1[118], w1_s0[118]}), .c ({new_AGEMA_signal_6445, new_AGEMA_signal_6444, addc_in[118]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_119_U1 ( .s (p256_sel), .b ({w0_s2[119], w0_s1[119], w0_s0[119]}), .a ({w1_s2[119], w1_s1[119], w1_s0[119]}), .c ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, addc_in[119]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_120_U1 ( .s (p256_sel), .b ({w0_s2[120], w0_s1[120], w0_s0[120]}), .a ({w1_s2[120], w1_s1[120], w1_s0[120]}), .c ({new_AGEMA_signal_6457, new_AGEMA_signal_6456, addc_in[120]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_121_U1 ( .s (p256_sel), .b ({w0_s2[121], w0_s1[121], w0_s0[121]}), .a ({w1_s2[121], w1_s1[121], w1_s0[121]}), .c ({new_AGEMA_signal_6463, new_AGEMA_signal_6462, addc_in[121]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_122_U1 ( .s (p256_sel), .b ({w0_s2[122], w0_s1[122], w0_s0[122]}), .a ({w1_s2[122], w1_s1[122], w1_s0[122]}), .c ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, addc_in[122]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_123_U1 ( .s (p256_sel), .b ({w0_s2[123], w0_s1[123], w0_s0[123]}), .a ({w1_s2[123], w1_s1[123], w1_s0[123]}), .c ({new_AGEMA_signal_6475, new_AGEMA_signal_6474, addc_in[123]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_124_U1 ( .s (p256_sel), .b ({w0_s2[124], w0_s1[124], w0_s0[124]}), .a ({w1_s2[124], w1_s1[124], w1_s0[124]}), .c ({new_AGEMA_signal_6481, new_AGEMA_signal_6480, addc_in[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_125_U1 ( .s (p256_sel), .b ({w0_s2[125], w0_s1[125], w0_s0[125]}), .a ({w1_s2[125], w1_s1[125], w1_s0[125]}), .c ({new_AGEMA_signal_6487, new_AGEMA_signal_6486, addc_in[125]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_126_U1 ( .s (p256_sel), .b ({w0_s2[126], w0_s1[126], w0_s0[126]}), .a ({w1_s2[126], w1_s1[126], w1_s0[126]}), .c ({new_AGEMA_signal_6493, new_AGEMA_signal_6492, addc_in[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst1_MUXInst_127_U1 ( .s (p256_sel), .b ({w0_s2[127], w0_s1[127], w0_s0[127]}), .a ({w1_s2[127], w1_s1[127], w1_s0[127]}), .c ({new_AGEMA_signal_6499, new_AGEMA_signal_6498, addc_in[127]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_U8 ( .a ({new_AGEMA_signal_6501, new_AGEMA_signal_6500, add_sub1_0_n8}), .b ({1'b0, 1'b0, add_sub1_0_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, add_sub1_0_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_U7 ( .a ({new_AGEMA_signal_6499, new_AGEMA_signal_6498, addc_in[127]}), .b ({1'b0, 1'b0, p256_sel}), .c ({new_AGEMA_signal_6501, new_AGEMA_signal_6500, add_sub1_0_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_U6 ( .a ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, add_sub1_0_n7}), .b ({1'b0, 1'b0, add_sub1_0_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_7535, new_AGEMA_signal_7534, add_sub1_0_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_U5 ( .a ({new_AGEMA_signal_6493, new_AGEMA_signal_6492, addc_in[126]}), .b ({1'b0, 1'b0, add_sub1_0_addc_rom_ic_out[2]}), .c ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, add_sub1_0_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_U4 ( .a ({new_AGEMA_signal_6503, new_AGEMA_signal_6502, add_sub1_0_n6}), .b ({1'b0, 1'b0, add_sub1_0_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_7537, new_AGEMA_signal_7536, add_sub1_0_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_U3 ( .a ({new_AGEMA_signal_6487, new_AGEMA_signal_6486, addc_in[125]}), .b ({1'b0, 1'b0, add_sub1_0_addc_rom_ic_out[1]}), .c ({new_AGEMA_signal_6503, new_AGEMA_signal_6502, add_sub1_0_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_U2 ( .a ({new_AGEMA_signal_7365, new_AGEMA_signal_7364, add_sub1_0_n5}), .b ({1'b0, 1'b0, add_sub1_0_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_7539, new_AGEMA_signal_7538, add_sub1_0_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_U1 ( .a ({new_AGEMA_signal_6481, new_AGEMA_signal_6480, addc_in[124]}), .b ({1'b0, 1'b0, add_sub1_0_addc_rom_ic_out[0]}), .c ({new_AGEMA_signal_7365, new_AGEMA_signal_7364, add_sub1_0_n5}) ) ;
    XOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U4 ( .A (1'b0), .B (p256_sel), .Z (add_sub1_0_addc_rom_ic_out[1]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_0_addc_rom_ic1_ANF_0_n2), .B (1'b0), .ZN (add_sub1_0_addc_rom_ic_out[0]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U2 ( .A (1'b0), .B (add_sub1_0_addc_rom_ic_out[2]), .ZN (add_sub1_0_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_0_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_0_addc_rom_ic_out[2]) ) ;
    AND2_X1 add_sub1_0_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b0), .A2 (1'b0), .ZN (add_sub1_0_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n21), .B (add_sub1_0_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_0_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n19), .B (add_sub1_0_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t5), .B (add_sub1_0_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t7), .B (add_sub1_0_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n17), .B (add_sub1_0_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_0_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t6), .B (add_sub1_0_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n14), .B (add_sub1_0_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_0_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t5), .B (add_sub1_0_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_0_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_0_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n12), .B (add_sub1_0_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_0_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t0), .B (add_sub1_0_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t4), .B (add_sub1_0_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_0_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_0_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_0_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_0_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, add_sub1_0_addc_out[3]}), .b ({new_AGEMA_signal_7535, new_AGEMA_signal_7534, add_sub1_0_addc_out[2]}), .c ({new_AGEMA_signal_8005, new_AGEMA_signal_8004, add_sub1_0_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_7537, new_AGEMA_signal_7536, add_sub1_0_addc_out[1]}), .b ({new_AGEMA_signal_7535, new_AGEMA_signal_7534, add_sub1_0_addc_out[2]}), .c ({new_AGEMA_signal_8007, new_AGEMA_signal_8006, add_sub1_0_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_6475, new_AGEMA_signal_6474, addc_in[123]}), .b ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, addc_in[122]}), .c ({new_AGEMA_signal_6505, new_AGEMA_signal_6504, add_sub1_0_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_6463, new_AGEMA_signal_6462, addc_in[121]}), .b ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, addc_in[122]}), .c ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, add_sub1_0_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, addc_in[119]}), .b ({new_AGEMA_signal_6445, new_AGEMA_signal_6444, addc_in[118]}), .c ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, add_sub1_0_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_6439, new_AGEMA_signal_6438, addc_in[117]}), .b ({new_AGEMA_signal_6445, new_AGEMA_signal_6444, addc_in[118]}), .c ({new_AGEMA_signal_6521, new_AGEMA_signal_6520, add_sub1_0_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_6427, new_AGEMA_signal_6426, addc_in[115]}), .b ({new_AGEMA_signal_6421, new_AGEMA_signal_6420, addc_in[114]}), .c ({new_AGEMA_signal_6533, new_AGEMA_signal_6532, add_sub1_0_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, addc_in[113]}), .b ({new_AGEMA_signal_6421, new_AGEMA_signal_6420, addc_in[114]}), .c ({new_AGEMA_signal_6535, new_AGEMA_signal_6534, add_sub1_0_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_6403, new_AGEMA_signal_6402, addc_in[111]}), .b ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, addc_in[110]}), .c ({new_AGEMA_signal_6547, new_AGEMA_signal_6546, add_sub1_0_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_6391, new_AGEMA_signal_6390, addc_in[109]}), .b ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, addc_in[110]}), .c ({new_AGEMA_signal_6549, new_AGEMA_signal_6548, add_sub1_0_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, addc_in[107]}), .b ({new_AGEMA_signal_6373, new_AGEMA_signal_6372, addc_in[106]}), .c ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, add_sub1_0_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_6367, new_AGEMA_signal_6366, addc_in[105]}), .b ({new_AGEMA_signal_6373, new_AGEMA_signal_6372, addc_in[106]}), .c ({new_AGEMA_signal_6563, new_AGEMA_signal_6562, add_sub1_0_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_6355, new_AGEMA_signal_6354, addc_in[103]}), .b ({new_AGEMA_signal_6349, new_AGEMA_signal_6348, addc_in[102]}), .c ({new_AGEMA_signal_6575, new_AGEMA_signal_6574, add_sub1_0_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, addc_in[101]}), .b ({new_AGEMA_signal_6349, new_AGEMA_signal_6348, addc_in[102]}), .c ({new_AGEMA_signal_6577, new_AGEMA_signal_6576, add_sub1_0_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_6331, new_AGEMA_signal_6330, addc_in[99]}), .b ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, addc_in[98]}), .c ({new_AGEMA_signal_6589, new_AGEMA_signal_6588, add_sub1_0_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_6319, new_AGEMA_signal_6318, addc_in[97]}), .b ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, addc_in[98]}), .c ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, add_sub1_0_subc_rom_sbox_0_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_U8 ( .a ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, add_sub1_1_n8}), .b ({1'b0, 1'b0, add_sub1_1_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_7555, new_AGEMA_signal_7554, add_sub1_1_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_U7 ( .a ({new_AGEMA_signal_6307, new_AGEMA_signal_6306, addc_in[95]}), .b ({1'b0, 1'b0, p256_sel}), .c ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, add_sub1_1_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_U6 ( .a ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, add_sub1_1_n7}), .b ({1'b0, 1'b0, add_sub1_1_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, add_sub1_1_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_U5 ( .a ({new_AGEMA_signal_6301, new_AGEMA_signal_6300, addc_in[94]}), .b ({1'b0, 1'b0, add_sub1_1_addc_rom_ic_out[2]}), .c ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, add_sub1_1_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_U4 ( .a ({new_AGEMA_signal_6605, new_AGEMA_signal_6604, add_sub1_1_n6}), .b ({1'b0, 1'b0, add_sub1_1_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_7559, new_AGEMA_signal_7558, add_sub1_1_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_U3 ( .a ({new_AGEMA_signal_6295, new_AGEMA_signal_6294, addc_in[93]}), .b ({1'b0, 1'b0, add_sub1_1_addc_rom_ic_out[1]}), .c ({new_AGEMA_signal_6605, new_AGEMA_signal_6604, add_sub1_1_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_U2 ( .a ({new_AGEMA_signal_7395, new_AGEMA_signal_7394, add_sub1_1_n5}), .b ({1'b0, 1'b0, add_sub1_1_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_7561, new_AGEMA_signal_7560, add_sub1_1_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_U1 ( .a ({new_AGEMA_signal_6289, new_AGEMA_signal_6288, addc_in[92]}), .b ({1'b0, 1'b0, add_sub1_1_addc_rom_ic_out[0]}), .c ({new_AGEMA_signal_7395, new_AGEMA_signal_7394, add_sub1_1_n5}) ) ;
    XOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U4 ( .A (1'b0), .B (p256_sel), .Z (add_sub1_1_addc_rom_ic_out[1]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_1_addc_rom_ic1_ANF_0_n2), .B (1'b1), .ZN (add_sub1_1_addc_rom_ic_out[0]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U2 ( .A (1'b0), .B (add_sub1_1_addc_rom_ic_out[2]), .ZN (add_sub1_1_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_1_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_1_addc_rom_ic_out[2]) ) ;
    AND2_X1 add_sub1_1_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b1), .A2 (1'b0), .ZN (add_sub1_1_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n21), .B (add_sub1_1_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_1_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n19), .B (add_sub1_1_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t5), .B (add_sub1_1_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t7), .B (add_sub1_1_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n17), .B (add_sub1_1_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_1_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t6), .B (add_sub1_1_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n14), .B (add_sub1_1_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_1_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t5), .B (add_sub1_1_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_1_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_1_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n12), .B (add_sub1_1_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_1_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t0), .B (add_sub1_1_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t4), .B (add_sub1_1_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_1_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_1_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_1_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_1_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_7555, new_AGEMA_signal_7554, add_sub1_1_addc_out[3]}), .b ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, add_sub1_1_addc_out[2]}), .c ({new_AGEMA_signal_8047, new_AGEMA_signal_8046, add_sub1_1_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_7559, new_AGEMA_signal_7558, add_sub1_1_addc_out[1]}), .b ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, add_sub1_1_addc_out[2]}), .c ({new_AGEMA_signal_8049, new_AGEMA_signal_8048, add_sub1_1_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_6283, new_AGEMA_signal_6282, addc_in[91]}), .b ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, addc_in[90]}), .c ({new_AGEMA_signal_6607, new_AGEMA_signal_6606, add_sub1_1_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, addc_in[89]}), .b ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, addc_in[90]}), .c ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, add_sub1_1_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_6259, new_AGEMA_signal_6258, addc_in[87]}), .b ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, addc_in[86]}), .c ({new_AGEMA_signal_6621, new_AGEMA_signal_6620, add_sub1_1_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_6247, new_AGEMA_signal_6246, addc_in[85]}), .b ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, addc_in[86]}), .c ({new_AGEMA_signal_6623, new_AGEMA_signal_6622, add_sub1_1_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, addc_in[83]}), .b ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, addc_in[82]}), .c ({new_AGEMA_signal_6635, new_AGEMA_signal_6634, add_sub1_1_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_6223, new_AGEMA_signal_6222, addc_in[81]}), .b ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, addc_in[82]}), .c ({new_AGEMA_signal_6637, new_AGEMA_signal_6636, add_sub1_1_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_6211, new_AGEMA_signal_6210, addc_in[79]}), .b ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, addc_in[78]}), .c ({new_AGEMA_signal_6649, new_AGEMA_signal_6648, add_sub1_1_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, addc_in[77]}), .b ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, addc_in[78]}), .c ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, add_sub1_1_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, addc_in[75]}), .b ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, addc_in[74]}), .c ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, add_sub1_1_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, addc_in[73]}), .b ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, addc_in[74]}), .c ({new_AGEMA_signal_6665, new_AGEMA_signal_6664, add_sub1_1_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, addc_in[71]}), .b ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, addc_in[70]}), .c ({new_AGEMA_signal_6677, new_AGEMA_signal_6676, add_sub1_1_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, addc_in[69]}), .b ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, addc_in[70]}), .c ({new_AGEMA_signal_6679, new_AGEMA_signal_6678, add_sub1_1_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, addc_in[67]}), .b ({new_AGEMA_signal_6133, new_AGEMA_signal_6132, addc_in[66]}), .c ({new_AGEMA_signal_6691, new_AGEMA_signal_6690, add_sub1_1_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, addc_in[65]}), .b ({new_AGEMA_signal_6133, new_AGEMA_signal_6132, addc_in[66]}), .c ({new_AGEMA_signal_6693, new_AGEMA_signal_6692, add_sub1_1_subc_rom_sbox_0_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_U8 ( .a ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, add_sub1_2_n8}), .b ({1'b0, 1'b0, add_sub1_2_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_7577, new_AGEMA_signal_7576, add_sub1_2_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_U7 ( .a ({new_AGEMA_signal_6115, new_AGEMA_signal_6114, addc_in[63]}), .b ({1'b0, 1'b0, p256_sel}), .c ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, add_sub1_2_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_U6 ( .a ({new_AGEMA_signal_7053, new_AGEMA_signal_7052, add_sub1_2_n7}), .b ({1'b0, 1'b0, add_sub1_2_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_7579, new_AGEMA_signal_7578, add_sub1_2_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_U5 ( .a ({new_AGEMA_signal_6109, new_AGEMA_signal_6108, addc_in[62]}), .b ({1'b0, 1'b0, add_sub1_2_addc_rom_ic_out[2]}), .c ({new_AGEMA_signal_7053, new_AGEMA_signal_7052, add_sub1_2_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_U4 ( .a ({new_AGEMA_signal_6707, new_AGEMA_signal_6706, add_sub1_2_n6}), .b ({1'b0, 1'b0, add_sub1_2_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_7581, new_AGEMA_signal_7580, add_sub1_2_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_U3 ( .a ({new_AGEMA_signal_6103, new_AGEMA_signal_6102, addc_in[61]}), .b ({1'b0, 1'b0, add_sub1_2_addc_rom_ic_out[1]}), .c ({new_AGEMA_signal_6707, new_AGEMA_signal_6706, add_sub1_2_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_U2 ( .a ({new_AGEMA_signal_7425, new_AGEMA_signal_7424, add_sub1_2_n5}), .b ({1'b0, 1'b0, add_sub1_2_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_7583, new_AGEMA_signal_7582, add_sub1_2_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_U1 ( .a ({new_AGEMA_signal_6097, new_AGEMA_signal_6096, addc_in[60]}), .b ({1'b0, 1'b0, add_sub1_2_addc_rom_ic_out[0]}), .c ({new_AGEMA_signal_7425, new_AGEMA_signal_7424, add_sub1_2_n5}) ) ;
    XOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U4 ( .A (1'b1), .B (p256_sel), .Z (add_sub1_2_addc_rom_ic_out[1]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_2_addc_rom_ic1_ANF_0_n2), .B (1'b0), .ZN (add_sub1_2_addc_rom_ic_out[0]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U2 ( .A (1'b1), .B (add_sub1_2_addc_rom_ic_out[2]), .ZN (add_sub1_2_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_2_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_2_addc_rom_ic_out[2]) ) ;
    AND2_X1 add_sub1_2_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b0), .A2 (1'b1), .ZN (add_sub1_2_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n21), .B (add_sub1_2_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_2_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n19), .B (add_sub1_2_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t5), .B (add_sub1_2_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t7), .B (add_sub1_2_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n17), .B (add_sub1_2_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_2_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t6), .B (add_sub1_2_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n14), .B (add_sub1_2_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_2_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t5), .B (add_sub1_2_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_2_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_2_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n12), .B (add_sub1_2_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_2_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t0), .B (add_sub1_2_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t4), .B (add_sub1_2_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_2_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_2_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_2_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_2_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_7577, new_AGEMA_signal_7576, add_sub1_2_addc_out[3]}), .b ({new_AGEMA_signal_7579, new_AGEMA_signal_7578, add_sub1_2_addc_out[2]}), .c ({new_AGEMA_signal_8089, new_AGEMA_signal_8088, add_sub1_2_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_7581, new_AGEMA_signal_7580, add_sub1_2_addc_out[1]}), .b ({new_AGEMA_signal_7579, new_AGEMA_signal_7578, add_sub1_2_addc_out[2]}), .c ({new_AGEMA_signal_8091, new_AGEMA_signal_8090, add_sub1_2_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, addc_in[59]}), .b ({new_AGEMA_signal_6085, new_AGEMA_signal_6084, addc_in[58]}), .c ({new_AGEMA_signal_6709, new_AGEMA_signal_6708, add_sub1_2_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, addc_in[57]}), .b ({new_AGEMA_signal_6085, new_AGEMA_signal_6084, addc_in[58]}), .c ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, add_sub1_2_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, addc_in[55]}), .b ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, addc_in[54]}), .c ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, add_sub1_2_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, addc_in[53]}), .b ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, addc_in[54]}), .c ({new_AGEMA_signal_6725, new_AGEMA_signal_6724, add_sub1_2_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, addc_in[51]}), .b ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, addc_in[50]}), .c ({new_AGEMA_signal_6737, new_AGEMA_signal_6736, add_sub1_2_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, addc_in[49]}), .b ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, addc_in[50]}), .c ({new_AGEMA_signal_6739, new_AGEMA_signal_6738, add_sub1_2_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, addc_in[47]}), .b ({new_AGEMA_signal_6013, new_AGEMA_signal_6012, addc_in[46]}), .c ({new_AGEMA_signal_6751, new_AGEMA_signal_6750, add_sub1_2_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, addc_in[45]}), .b ({new_AGEMA_signal_6013, new_AGEMA_signal_6012, addc_in[46]}), .c ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, add_sub1_2_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, addc_in[43]}), .b ({new_AGEMA_signal_5989, new_AGEMA_signal_5988, addc_in[42]}), .c ({new_AGEMA_signal_6765, new_AGEMA_signal_6764, add_sub1_2_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, addc_in[41]}), .b ({new_AGEMA_signal_5989, new_AGEMA_signal_5988, addc_in[42]}), .c ({new_AGEMA_signal_6767, new_AGEMA_signal_6766, add_sub1_2_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, addc_in[39]}), .b ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, addc_in[38]}), .c ({new_AGEMA_signal_6779, new_AGEMA_signal_6778, add_sub1_2_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, addc_in[37]}), .b ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, addc_in[38]}), .c ({new_AGEMA_signal_6781, new_AGEMA_signal_6780, add_sub1_2_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, addc_in[35]}), .b ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, addc_in[34]}), .c ({new_AGEMA_signal_6793, new_AGEMA_signal_6792, add_sub1_2_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, addc_in[33]}), .b ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, addc_in[34]}), .c ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, add_sub1_2_subc_rom_sbox_0_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_U8 ( .a ({new_AGEMA_signal_6807, new_AGEMA_signal_6806, add_sub1_3_n8}), .b ({1'b0, 1'b0, add_sub1_3_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_7599, new_AGEMA_signal_7598, add_sub1_3_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_U7 ( .a ({new_AGEMA_signal_5923, new_AGEMA_signal_5922, addc_in[31]}), .b ({1'b0, 1'b0, p256_sel}), .c ({new_AGEMA_signal_6807, new_AGEMA_signal_6806, add_sub1_3_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_U6 ( .a ({new_AGEMA_signal_7125, new_AGEMA_signal_7124, add_sub1_3_n7}), .b ({1'b0, 1'b0, add_sub1_3_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_7601, new_AGEMA_signal_7600, add_sub1_3_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_U5 ( .a ({new_AGEMA_signal_5917, new_AGEMA_signal_5916, addc_in[30]}), .b ({1'b0, 1'b0, add_sub1_3_addc_rom_ic_out_2_}), .c ({new_AGEMA_signal_7125, new_AGEMA_signal_7124, add_sub1_3_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_U4 ( .a ({new_AGEMA_signal_6809, new_AGEMA_signal_6808, add_sub1_3_n6}), .b ({1'b0, 1'b0, add_sub1_3_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_7603, new_AGEMA_signal_7602, add_sub1_3_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_U3 ( .a ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, addc_in[29]}), .b ({1'b0, 1'b0, add_sub1_3_addc_rom_ic_out_1_}), .c ({new_AGEMA_signal_6809, new_AGEMA_signal_6808, add_sub1_3_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_U2 ( .a ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, add_sub1_3_n5}), .b ({1'b0, 1'b0, add_sub1_3_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_7605, new_AGEMA_signal_7604, add_sub1_3_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_U1 ( .a ({new_AGEMA_signal_5905, new_AGEMA_signal_5904, addc_in[28]}), .b ({1'b0, 1'b0, add_sub1_3_addc_rom_ic_out_0_}), .c ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, add_sub1_3_n5}) ) ;
    XOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U4 ( .A (1'b1), .B (p256_sel), .Z (add_sub1_3_addc_rom_ic_out_1_) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_3_addc_rom_ic1_ANF_0_n2), .B (1'b1), .ZN (add_sub1_3_addc_rom_ic_out_0_) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U2 ( .A (1'b1), .B (add_sub1_3_addc_rom_ic_out_2_), .ZN (add_sub1_3_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_3_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_3_addc_rom_ic_out_2_) ) ;
    AND2_X1 add_sub1_3_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b1), .A2 (1'b1), .ZN (add_sub1_3_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n21), .B (add_sub1_3_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_3_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n19), .B (add_sub1_3_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t5), .B (add_sub1_3_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t7), .B (add_sub1_3_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n17), .B (add_sub1_3_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_3_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t6), .B (add_sub1_3_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n14), .B (add_sub1_3_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_3_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t5), .B (add_sub1_3_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_3_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_3_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n12), .B (add_sub1_3_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_3_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t0), .B (add_sub1_3_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t4), .B (add_sub1_3_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_3_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_3_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_3_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_3_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_7599, new_AGEMA_signal_7598, add_sub1_3_addc_out[3]}), .b ({new_AGEMA_signal_7601, new_AGEMA_signal_7600, add_sub1_3_addc_out[2]}), .c ({new_AGEMA_signal_8131, new_AGEMA_signal_8130, add_sub1_3_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_7603, new_AGEMA_signal_7602, add_sub1_3_addc_out[1]}), .b ({new_AGEMA_signal_7601, new_AGEMA_signal_7600, add_sub1_3_addc_out[2]}), .c ({new_AGEMA_signal_8133, new_AGEMA_signal_8132, add_sub1_3_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, addc_in[27]}), .b ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, addc_in[26]}), .c ({new_AGEMA_signal_6811, new_AGEMA_signal_6810, add_sub1_3_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, addc_in[25]}), .b ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, addc_in[26]}), .c ({new_AGEMA_signal_6813, new_AGEMA_signal_6812, add_sub1_3_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, addc_in[23]}), .b ({new_AGEMA_signal_5869, new_AGEMA_signal_5868, addc_in[22]}), .c ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, add_sub1_3_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, addc_in[21]}), .b ({new_AGEMA_signal_5869, new_AGEMA_signal_5868, addc_in[22]}), .c ({new_AGEMA_signal_6827, new_AGEMA_signal_6826, add_sub1_3_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, addc_in[19]}), .b ({new_AGEMA_signal_5845, new_AGEMA_signal_5844, addc_in[18]}), .c ({new_AGEMA_signal_6839, new_AGEMA_signal_6838, add_sub1_3_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, addc_in[17]}), .b ({new_AGEMA_signal_5845, new_AGEMA_signal_5844, addc_in[18]}), .c ({new_AGEMA_signal_6841, new_AGEMA_signal_6840, add_sub1_3_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, addc_in[15]}), .b ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, addc_in[14]}), .c ({new_AGEMA_signal_6853, new_AGEMA_signal_6852, add_sub1_3_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, addc_in[13]}), .b ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, addc_in[14]}), .c ({new_AGEMA_signal_6855, new_AGEMA_signal_6854, add_sub1_3_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, addc_in[11]}), .b ({new_AGEMA_signal_5797, new_AGEMA_signal_5796, addc_in[10]}), .c ({new_AGEMA_signal_6867, new_AGEMA_signal_6866, add_sub1_3_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, addc_in[9]}), .b ({new_AGEMA_signal_5797, new_AGEMA_signal_5796, addc_in[10]}), .c ({new_AGEMA_signal_6869, new_AGEMA_signal_6868, add_sub1_3_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, addc_in[7]}), .b ({new_AGEMA_signal_5773, new_AGEMA_signal_5772, addc_in[6]}), .c ({new_AGEMA_signal_6881, new_AGEMA_signal_6880, add_sub1_3_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, addc_in[5]}), .b ({new_AGEMA_signal_5773, new_AGEMA_signal_5772, addc_in[6]}), .c ({new_AGEMA_signal_6883, new_AGEMA_signal_6882, add_sub1_3_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, addc_in[3]}), .b ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, addc_in[2]}), .c ({new_AGEMA_signal_6895, new_AGEMA_signal_6894, add_sub1_3_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, addc_in[1]}), .b ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, addc_in[2]}), .c ({new_AGEMA_signal_6897, new_AGEMA_signal_6896, add_sub1_3_subc_rom_sbox_0_ANF_2_t5}) ) ;
    //ClockGatingController #(6) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_8619, new_AGEMA_signal_8618, add_sub1_0_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, add_sub1_0_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_8821, new_AGEMA_signal_8820, add_sub1_0_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_8011, new_AGEMA_signal_8010, add_sub1_0_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_8015, new_AGEMA_signal_8014, add_sub1_0_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, add_sub1_0_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_8017, new_AGEMA_signal_8016, add_sub1_0_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_7535, new_AGEMA_signal_7534, add_sub1_0_addc_out[2]}), .c ({new_AGEMA_signal_8619, new_AGEMA_signal_8618, add_sub1_0_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_8005, new_AGEMA_signal_8004, add_sub1_0_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_8621, new_AGEMA_signal_8620, add_sub1_0_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_8825, new_AGEMA_signal_8824, subc_out[124]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_8009, new_AGEMA_signal_8008, add_sub1_0_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_7539, new_AGEMA_signal_7538, add_sub1_0_addc_out[0]}), .c ({new_AGEMA_signal_8621, new_AGEMA_signal_8620, add_sub1_0_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_7537, new_AGEMA_signal_7536, add_sub1_0_addc_out[1]}), .b ({new_AGEMA_signal_7535, new_AGEMA_signal_7534, add_sub1_0_addc_out[2]}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_8009, new_AGEMA_signal_8008, add_sub1_0_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_7537, new_AGEMA_signal_7536, add_sub1_0_addc_out[1]}), .b ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, add_sub1_0_addc_out[3]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_8011, new_AGEMA_signal_8010, add_sub1_0_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_7535, new_AGEMA_signal_7534, add_sub1_0_addc_out[2]}), .b ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, add_sub1_0_addc_out[3]}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_8013, new_AGEMA_signal_8012, add_sub1_0_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_7539, new_AGEMA_signal_7538, add_sub1_0_addc_out[0]}), .b ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, add_sub1_0_addc_out[3]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_8015, new_AGEMA_signal_8014, add_sub1_0_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_7539, new_AGEMA_signal_7538, add_sub1_0_addc_out[0]}), .b ({new_AGEMA_signal_7537, new_AGEMA_signal_7536, add_sub1_0_addc_out[1]}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_8017, new_AGEMA_signal_8016, add_sub1_0_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_6913, new_AGEMA_signal_6912, add_sub1_0_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_6911, new_AGEMA_signal_6910, add_sub1_0_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_7197, new_AGEMA_signal_7196, add_sub1_0_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_6511, new_AGEMA_signal_6510, add_sub1_0_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_6515, new_AGEMA_signal_6514, add_sub1_0_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_6911, new_AGEMA_signal_6910, add_sub1_0_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_6517, new_AGEMA_signal_6516, add_sub1_0_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, addc_in[122]}), .c ({new_AGEMA_signal_6913, new_AGEMA_signal_6912, add_sub1_0_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_6505, new_AGEMA_signal_6504, add_sub1_0_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_6915, new_AGEMA_signal_6914, add_sub1_0_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_7201, new_AGEMA_signal_7200, subc_out[120]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_6509, new_AGEMA_signal_6508, add_sub1_0_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_6457, new_AGEMA_signal_6456, addc_in[120]}), .c ({new_AGEMA_signal_6915, new_AGEMA_signal_6914, add_sub1_0_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6463, new_AGEMA_signal_6462, addc_in[121]}), .b ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, addc_in[122]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_6509, new_AGEMA_signal_6508, add_sub1_0_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6463, new_AGEMA_signal_6462, addc_in[121]}), .b ({new_AGEMA_signal_6475, new_AGEMA_signal_6474, addc_in[123]}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_6511, new_AGEMA_signal_6510, add_sub1_0_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, addc_in[122]}), .b ({new_AGEMA_signal_6475, new_AGEMA_signal_6474, addc_in[123]}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, add_sub1_0_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6457, new_AGEMA_signal_6456, addc_in[120]}), .b ({new_AGEMA_signal_6475, new_AGEMA_signal_6474, addc_in[123]}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_6515, new_AGEMA_signal_6514, add_sub1_0_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6457, new_AGEMA_signal_6456, addc_in[120]}), .b ({new_AGEMA_signal_6463, new_AGEMA_signal_6462, addc_in[121]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_6517, new_AGEMA_signal_6516, add_sub1_0_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_6923, new_AGEMA_signal_6922, add_sub1_0_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_6921, new_AGEMA_signal_6920, add_sub1_0_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_7203, new_AGEMA_signal_7202, add_sub1_0_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_6525, new_AGEMA_signal_6524, add_sub1_0_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_6529, new_AGEMA_signal_6528, add_sub1_0_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_6921, new_AGEMA_signal_6920, add_sub1_0_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, add_sub1_0_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_6445, new_AGEMA_signal_6444, addc_in[118]}), .c ({new_AGEMA_signal_6923, new_AGEMA_signal_6922, add_sub1_0_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, add_sub1_0_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_6925, new_AGEMA_signal_6924, add_sub1_0_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_7207, new_AGEMA_signal_7206, subc_out[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, add_sub1_0_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, addc_in[116]}), .c ({new_AGEMA_signal_6925, new_AGEMA_signal_6924, add_sub1_0_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6439, new_AGEMA_signal_6438, addc_in[117]}), .b ({new_AGEMA_signal_6445, new_AGEMA_signal_6444, addc_in[118]}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, add_sub1_0_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6439, new_AGEMA_signal_6438, addc_in[117]}), .b ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, addc_in[119]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_6525, new_AGEMA_signal_6524, add_sub1_0_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6445, new_AGEMA_signal_6444, addc_in[118]}), .b ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, addc_in[119]}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_6527, new_AGEMA_signal_6526, add_sub1_0_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, addc_in[116]}), .b ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, addc_in[119]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_6529, new_AGEMA_signal_6528, add_sub1_0_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, addc_in[116]}), .b ({new_AGEMA_signal_6439, new_AGEMA_signal_6438, addc_in[117]}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, add_sub1_0_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_6933, new_AGEMA_signal_6932, add_sub1_0_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_6931, new_AGEMA_signal_6930, add_sub1_0_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_7209, new_AGEMA_signal_7208, add_sub1_0_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_6539, new_AGEMA_signal_6538, add_sub1_0_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, add_sub1_0_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_6931, new_AGEMA_signal_6930, add_sub1_0_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_6545, new_AGEMA_signal_6544, add_sub1_0_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_6421, new_AGEMA_signal_6420, addc_in[114]}), .c ({new_AGEMA_signal_6933, new_AGEMA_signal_6932, add_sub1_0_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_6533, new_AGEMA_signal_6532, add_sub1_0_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_6935, new_AGEMA_signal_6934, add_sub1_0_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_7213, new_AGEMA_signal_7212, subc_out[112]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, add_sub1_0_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_6409, new_AGEMA_signal_6408, addc_in[112]}), .c ({new_AGEMA_signal_6935, new_AGEMA_signal_6934, add_sub1_0_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, addc_in[113]}), .b ({new_AGEMA_signal_6421, new_AGEMA_signal_6420, addc_in[114]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, add_sub1_0_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, addc_in[113]}), .b ({new_AGEMA_signal_6427, new_AGEMA_signal_6426, addc_in[115]}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_6539, new_AGEMA_signal_6538, add_sub1_0_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6421, new_AGEMA_signal_6420, addc_in[114]}), .b ({new_AGEMA_signal_6427, new_AGEMA_signal_6426, addc_in[115]}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_6541, new_AGEMA_signal_6540, add_sub1_0_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6409, new_AGEMA_signal_6408, addc_in[112]}), .b ({new_AGEMA_signal_6427, new_AGEMA_signal_6426, addc_in[115]}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, add_sub1_0_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6409, new_AGEMA_signal_6408, addc_in[112]}), .b ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, addc_in[113]}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_6545, new_AGEMA_signal_6544, add_sub1_0_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_6943, new_AGEMA_signal_6942, add_sub1_0_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_6941, new_AGEMA_signal_6940, add_sub1_0_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, add_sub1_0_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_6553, new_AGEMA_signal_6552, add_sub1_0_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_6557, new_AGEMA_signal_6556, add_sub1_0_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_6941, new_AGEMA_signal_6940, add_sub1_0_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_6559, new_AGEMA_signal_6558, add_sub1_0_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, addc_in[110]}), .c ({new_AGEMA_signal_6943, new_AGEMA_signal_6942, add_sub1_0_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_6547, new_AGEMA_signal_6546, add_sub1_0_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_6945, new_AGEMA_signal_6944, add_sub1_0_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_7219, new_AGEMA_signal_7218, subc_out[108]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_6551, new_AGEMA_signal_6550, add_sub1_0_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_6385, new_AGEMA_signal_6384, addc_in[108]}), .c ({new_AGEMA_signal_6945, new_AGEMA_signal_6944, add_sub1_0_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6391, new_AGEMA_signal_6390, addc_in[109]}), .b ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, addc_in[110]}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_6551, new_AGEMA_signal_6550, add_sub1_0_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6391, new_AGEMA_signal_6390, addc_in[109]}), .b ({new_AGEMA_signal_6403, new_AGEMA_signal_6402, addc_in[111]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_6553, new_AGEMA_signal_6552, add_sub1_0_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, addc_in[110]}), .b ({new_AGEMA_signal_6403, new_AGEMA_signal_6402, addc_in[111]}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, add_sub1_0_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6385, new_AGEMA_signal_6384, addc_in[108]}), .b ({new_AGEMA_signal_6403, new_AGEMA_signal_6402, addc_in[111]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_6557, new_AGEMA_signal_6556, add_sub1_0_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6385, new_AGEMA_signal_6384, addc_in[108]}), .b ({new_AGEMA_signal_6391, new_AGEMA_signal_6390, addc_in[109]}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_6559, new_AGEMA_signal_6558, add_sub1_0_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_6953, new_AGEMA_signal_6952, add_sub1_0_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, add_sub1_0_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, add_sub1_0_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, add_sub1_0_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_6571, new_AGEMA_signal_6570, add_sub1_0_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, add_sub1_0_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_6573, new_AGEMA_signal_6572, add_sub1_0_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_6373, new_AGEMA_signal_6372, addc_in[106]}), .c ({new_AGEMA_signal_6953, new_AGEMA_signal_6952, add_sub1_0_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, add_sub1_0_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_6955, new_AGEMA_signal_6954, add_sub1_0_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_7225, new_AGEMA_signal_7224, subc_out[104]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_6565, new_AGEMA_signal_6564, add_sub1_0_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, addc_in[104]}), .c ({new_AGEMA_signal_6955, new_AGEMA_signal_6954, add_sub1_0_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6367, new_AGEMA_signal_6366, addc_in[105]}), .b ({new_AGEMA_signal_6373, new_AGEMA_signal_6372, addc_in[106]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_6565, new_AGEMA_signal_6564, add_sub1_0_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6367, new_AGEMA_signal_6366, addc_in[105]}), .b ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, addc_in[107]}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, add_sub1_0_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6373, new_AGEMA_signal_6372, addc_in[106]}), .b ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, addc_in[107]}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_6569, new_AGEMA_signal_6568, add_sub1_0_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, addc_in[104]}), .b ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, addc_in[107]}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_6571, new_AGEMA_signal_6570, add_sub1_0_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, addc_in[104]}), .b ({new_AGEMA_signal_6367, new_AGEMA_signal_6366, addc_in[105]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_6573, new_AGEMA_signal_6572, add_sub1_0_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_6963, new_AGEMA_signal_6962, add_sub1_0_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_6961, new_AGEMA_signal_6960, add_sub1_0_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_7227, new_AGEMA_signal_7226, add_sub1_0_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_6581, new_AGEMA_signal_6580, add_sub1_0_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, add_sub1_0_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_6961, new_AGEMA_signal_6960, add_sub1_0_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_6587, new_AGEMA_signal_6586, add_sub1_0_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_6349, new_AGEMA_signal_6348, addc_in[102]}), .c ({new_AGEMA_signal_6963, new_AGEMA_signal_6962, add_sub1_0_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_6575, new_AGEMA_signal_6574, add_sub1_0_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_6965, new_AGEMA_signal_6964, add_sub1_0_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_7231, new_AGEMA_signal_7230, subc_out[100]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, add_sub1_0_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_6337, new_AGEMA_signal_6336, addc_in[100]}), .c ({new_AGEMA_signal_6965, new_AGEMA_signal_6964, add_sub1_0_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, addc_in[101]}), .b ({new_AGEMA_signal_6349, new_AGEMA_signal_6348, addc_in[102]}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, add_sub1_0_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, addc_in[101]}), .b ({new_AGEMA_signal_6355, new_AGEMA_signal_6354, addc_in[103]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_6581, new_AGEMA_signal_6580, add_sub1_0_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6349, new_AGEMA_signal_6348, addc_in[102]}), .b ({new_AGEMA_signal_6355, new_AGEMA_signal_6354, addc_in[103]}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_6583, new_AGEMA_signal_6582, add_sub1_0_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6337, new_AGEMA_signal_6336, addc_in[100]}), .b ({new_AGEMA_signal_6355, new_AGEMA_signal_6354, addc_in[103]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, add_sub1_0_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6337, new_AGEMA_signal_6336, addc_in[100]}), .b ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, addc_in[101]}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_6587, new_AGEMA_signal_6586, add_sub1_0_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_6973, new_AGEMA_signal_6972, add_sub1_0_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_6971, new_AGEMA_signal_6970, add_sub1_0_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, add_sub1_0_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_6595, new_AGEMA_signal_6594, add_sub1_0_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_6599, new_AGEMA_signal_6598, add_sub1_0_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_6971, new_AGEMA_signal_6970, add_sub1_0_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_6601, new_AGEMA_signal_6600, add_sub1_0_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, addc_in[98]}), .c ({new_AGEMA_signal_6973, new_AGEMA_signal_6972, add_sub1_0_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_6589, new_AGEMA_signal_6588, add_sub1_0_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_6975, new_AGEMA_signal_6974, add_sub1_0_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_7237, new_AGEMA_signal_7236, subc_out[96]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_6593, new_AGEMA_signal_6592, add_sub1_0_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_6313, new_AGEMA_signal_6312, addc_in[96]}), .c ({new_AGEMA_signal_6975, new_AGEMA_signal_6974, add_sub1_0_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6319, new_AGEMA_signal_6318, addc_in[97]}), .b ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, addc_in[98]}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_6593, new_AGEMA_signal_6592, add_sub1_0_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6319, new_AGEMA_signal_6318, addc_in[97]}), .b ({new_AGEMA_signal_6331, new_AGEMA_signal_6330, addc_in[99]}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_6595, new_AGEMA_signal_6594, add_sub1_0_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, addc_in[98]}), .b ({new_AGEMA_signal_6331, new_AGEMA_signal_6330, addc_in[99]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_6597, new_AGEMA_signal_6596, add_sub1_0_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6313, new_AGEMA_signal_6312, addc_in[96]}), .b ({new_AGEMA_signal_6331, new_AGEMA_signal_6330, addc_in[99]}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_6599, new_AGEMA_signal_6598, add_sub1_0_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6313, new_AGEMA_signal_6312, addc_in[96]}), .b ({new_AGEMA_signal_6319, new_AGEMA_signal_6318, addc_in[97]}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_6601, new_AGEMA_signal_6600, add_sub1_0_subc_rom_sbox_0_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_8643, new_AGEMA_signal_8642, add_sub1_1_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_8641, new_AGEMA_signal_8640, add_sub1_1_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_8827, new_AGEMA_signal_8826, add_sub1_1_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_8053, new_AGEMA_signal_8052, add_sub1_1_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_8057, new_AGEMA_signal_8056, add_sub1_1_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_8641, new_AGEMA_signal_8640, add_sub1_1_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_8059, new_AGEMA_signal_8058, add_sub1_1_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, add_sub1_1_addc_out[2]}), .c ({new_AGEMA_signal_8643, new_AGEMA_signal_8642, add_sub1_1_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_8047, new_AGEMA_signal_8046, add_sub1_1_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_8645, new_AGEMA_signal_8644, add_sub1_1_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_8831, new_AGEMA_signal_8830, subc_out[92]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_8051, new_AGEMA_signal_8050, add_sub1_1_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_7561, new_AGEMA_signal_7560, add_sub1_1_addc_out[0]}), .c ({new_AGEMA_signal_8645, new_AGEMA_signal_8644, add_sub1_1_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_7559, new_AGEMA_signal_7558, add_sub1_1_addc_out[1]}), .b ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, add_sub1_1_addc_out[2]}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_8051, new_AGEMA_signal_8050, add_sub1_1_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_7559, new_AGEMA_signal_7558, add_sub1_1_addc_out[1]}), .b ({new_AGEMA_signal_7555, new_AGEMA_signal_7554, add_sub1_1_addc_out[3]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_8053, new_AGEMA_signal_8052, add_sub1_1_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, add_sub1_1_addc_out[2]}), .b ({new_AGEMA_signal_7555, new_AGEMA_signal_7554, add_sub1_1_addc_out[3]}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_8055, new_AGEMA_signal_8054, add_sub1_1_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_7561, new_AGEMA_signal_7560, add_sub1_1_addc_out[0]}), .b ({new_AGEMA_signal_7555, new_AGEMA_signal_7554, add_sub1_1_addc_out[3]}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_8057, new_AGEMA_signal_8056, add_sub1_1_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_7561, new_AGEMA_signal_7560, add_sub1_1_addc_out[0]}), .b ({new_AGEMA_signal_7559, new_AGEMA_signal_7558, add_sub1_1_addc_out[1]}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_8059, new_AGEMA_signal_8058, add_sub1_1_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_6985, new_AGEMA_signal_6984, add_sub1_1_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_6983, new_AGEMA_signal_6982, add_sub1_1_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, add_sub1_1_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, add_sub1_1_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_6617, new_AGEMA_signal_6616, add_sub1_1_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_6983, new_AGEMA_signal_6982, add_sub1_1_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_6619, new_AGEMA_signal_6618, add_sub1_1_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, addc_in[90]}), .c ({new_AGEMA_signal_6985, new_AGEMA_signal_6984, add_sub1_1_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_6607, new_AGEMA_signal_6606, add_sub1_1_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, add_sub1_1_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_7243, new_AGEMA_signal_7242, subc_out[88]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_6611, new_AGEMA_signal_6610, add_sub1_1_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, addc_in[88]}), .c ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, add_sub1_1_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, addc_in[89]}), .b ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, addc_in[90]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_6611, new_AGEMA_signal_6610, add_sub1_1_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, addc_in[89]}), .b ({new_AGEMA_signal_6283, new_AGEMA_signal_6282, addc_in[91]}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, add_sub1_1_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, addc_in[90]}), .b ({new_AGEMA_signal_6283, new_AGEMA_signal_6282, addc_in[91]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, add_sub1_1_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, addc_in[88]}), .b ({new_AGEMA_signal_6283, new_AGEMA_signal_6282, addc_in[91]}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_6617, new_AGEMA_signal_6616, add_sub1_1_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, addc_in[88]}), .b ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, addc_in[89]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_6619, new_AGEMA_signal_6618, add_sub1_1_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_6995, new_AGEMA_signal_6994, add_sub1_1_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_6993, new_AGEMA_signal_6992, add_sub1_1_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, add_sub1_1_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, add_sub1_1_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, add_sub1_1_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_6993, new_AGEMA_signal_6992, add_sub1_1_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, add_sub1_1_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, addc_in[86]}), .c ({new_AGEMA_signal_6995, new_AGEMA_signal_6994, add_sub1_1_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_6621, new_AGEMA_signal_6620, add_sub1_1_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_6997, new_AGEMA_signal_6996, add_sub1_1_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_7249, new_AGEMA_signal_7248, subc_out[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_6625, new_AGEMA_signal_6624, add_sub1_1_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, addc_in[84]}), .c ({new_AGEMA_signal_6997, new_AGEMA_signal_6996, add_sub1_1_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6247, new_AGEMA_signal_6246, addc_in[85]}), .b ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, addc_in[86]}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_6625, new_AGEMA_signal_6624, add_sub1_1_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6247, new_AGEMA_signal_6246, addc_in[85]}), .b ({new_AGEMA_signal_6259, new_AGEMA_signal_6258, addc_in[87]}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, add_sub1_1_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, addc_in[86]}), .b ({new_AGEMA_signal_6259, new_AGEMA_signal_6258, addc_in[87]}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_6629, new_AGEMA_signal_6628, add_sub1_1_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, addc_in[84]}), .b ({new_AGEMA_signal_6259, new_AGEMA_signal_6258, addc_in[87]}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, add_sub1_1_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, addc_in[84]}), .b ({new_AGEMA_signal_6247, new_AGEMA_signal_6246, addc_in[85]}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, add_sub1_1_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_7005, new_AGEMA_signal_7004, add_sub1_1_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_7003, new_AGEMA_signal_7002, add_sub1_1_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_7251, new_AGEMA_signal_7250, add_sub1_1_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_6641, new_AGEMA_signal_6640, add_sub1_1_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_6645, new_AGEMA_signal_6644, add_sub1_1_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_7003, new_AGEMA_signal_7002, add_sub1_1_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_6647, new_AGEMA_signal_6646, add_sub1_1_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, addc_in[82]}), .c ({new_AGEMA_signal_7005, new_AGEMA_signal_7004, add_sub1_1_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_6635, new_AGEMA_signal_6634, add_sub1_1_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_7007, new_AGEMA_signal_7006, add_sub1_1_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_7255, new_AGEMA_signal_7254, subc_out[80]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, add_sub1_1_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, addc_in[80]}), .c ({new_AGEMA_signal_7007, new_AGEMA_signal_7006, add_sub1_1_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6223, new_AGEMA_signal_6222, addc_in[81]}), .b ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, addc_in[82]}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, add_sub1_1_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6223, new_AGEMA_signal_6222, addc_in[81]}), .b ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, addc_in[83]}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_6641, new_AGEMA_signal_6640, add_sub1_1_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, addc_in[82]}), .b ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, addc_in[83]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_6643, new_AGEMA_signal_6642, add_sub1_1_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, addc_in[80]}), .b ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, addc_in[83]}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_6645, new_AGEMA_signal_6644, add_sub1_1_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, addc_in[80]}), .b ({new_AGEMA_signal_6223, new_AGEMA_signal_6222, addc_in[81]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_6647, new_AGEMA_signal_6646, add_sub1_1_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_7015, new_AGEMA_signal_7014, add_sub1_1_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_7013, new_AGEMA_signal_7012, add_sub1_1_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_7257, new_AGEMA_signal_7256, add_sub1_1_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_6655, new_AGEMA_signal_6654, add_sub1_1_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_6659, new_AGEMA_signal_6658, add_sub1_1_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_7013, new_AGEMA_signal_7012, add_sub1_1_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_6661, new_AGEMA_signal_6660, add_sub1_1_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, addc_in[78]}), .c ({new_AGEMA_signal_7015, new_AGEMA_signal_7014, add_sub1_1_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_6649, new_AGEMA_signal_6648, add_sub1_1_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_7017, new_AGEMA_signal_7016, add_sub1_1_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_7261, new_AGEMA_signal_7260, subc_out[76]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_6653, new_AGEMA_signal_6652, add_sub1_1_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, addc_in[76]}), .c ({new_AGEMA_signal_7017, new_AGEMA_signal_7016, add_sub1_1_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, addc_in[77]}), .b ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, addc_in[78]}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_6653, new_AGEMA_signal_6652, add_sub1_1_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, addc_in[77]}), .b ({new_AGEMA_signal_6211, new_AGEMA_signal_6210, addc_in[79]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_6655, new_AGEMA_signal_6654, add_sub1_1_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, addc_in[78]}), .b ({new_AGEMA_signal_6211, new_AGEMA_signal_6210, addc_in[79]}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, add_sub1_1_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, addc_in[76]}), .b ({new_AGEMA_signal_6211, new_AGEMA_signal_6210, addc_in[79]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_6659, new_AGEMA_signal_6658, add_sub1_1_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, addc_in[76]}), .b ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, addc_in[77]}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_6661, new_AGEMA_signal_6660, add_sub1_1_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_7025, new_AGEMA_signal_7024, add_sub1_1_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_7023, new_AGEMA_signal_7022, add_sub1_1_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, add_sub1_1_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_6669, new_AGEMA_signal_6668, add_sub1_1_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_6673, new_AGEMA_signal_6672, add_sub1_1_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_7023, new_AGEMA_signal_7022, add_sub1_1_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, add_sub1_1_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, addc_in[74]}), .c ({new_AGEMA_signal_7025, new_AGEMA_signal_7024, add_sub1_1_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, add_sub1_1_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_7027, new_AGEMA_signal_7026, add_sub1_1_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_7267, new_AGEMA_signal_7266, subc_out[72]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_6667, new_AGEMA_signal_6666, add_sub1_1_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_6169, new_AGEMA_signal_6168, addc_in[72]}), .c ({new_AGEMA_signal_7027, new_AGEMA_signal_7026, add_sub1_1_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, addc_in[73]}), .b ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, addc_in[74]}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_6667, new_AGEMA_signal_6666, add_sub1_1_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, addc_in[73]}), .b ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, addc_in[75]}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_6669, new_AGEMA_signal_6668, add_sub1_1_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, addc_in[74]}), .b ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, addc_in[75]}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_6671, new_AGEMA_signal_6670, add_sub1_1_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6169, new_AGEMA_signal_6168, addc_in[72]}), .b ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, addc_in[75]}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_6673, new_AGEMA_signal_6672, add_sub1_1_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6169, new_AGEMA_signal_6168, addc_in[72]}), .b ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, addc_in[73]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, add_sub1_1_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_7035, new_AGEMA_signal_7034, add_sub1_1_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_7033, new_AGEMA_signal_7032, add_sub1_1_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_7269, new_AGEMA_signal_7268, add_sub1_1_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_6683, new_AGEMA_signal_6682, add_sub1_1_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, add_sub1_1_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_7033, new_AGEMA_signal_7032, add_sub1_1_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_6689, new_AGEMA_signal_6688, add_sub1_1_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, addc_in[70]}), .c ({new_AGEMA_signal_7035, new_AGEMA_signal_7034, add_sub1_1_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_6677, new_AGEMA_signal_6676, add_sub1_1_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_7037, new_AGEMA_signal_7036, add_sub1_1_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_7273, new_AGEMA_signal_7272, subc_out[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, add_sub1_1_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, addc_in[68]}), .c ({new_AGEMA_signal_7037, new_AGEMA_signal_7036, add_sub1_1_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, addc_in[69]}), .b ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, addc_in[70]}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, add_sub1_1_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, addc_in[69]}), .b ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, addc_in[71]}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_6683, new_AGEMA_signal_6682, add_sub1_1_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6157, new_AGEMA_signal_6156, addc_in[70]}), .b ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, addc_in[71]}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_6685, new_AGEMA_signal_6684, add_sub1_1_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, addc_in[68]}), .b ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, addc_in[71]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, add_sub1_1_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, addc_in[68]}), .b ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, addc_in[69]}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_6689, new_AGEMA_signal_6688, add_sub1_1_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_7045, new_AGEMA_signal_7044, add_sub1_1_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_7043, new_AGEMA_signal_7042, add_sub1_1_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_7275, new_AGEMA_signal_7274, add_sub1_1_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_6697, new_AGEMA_signal_6696, add_sub1_1_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_6701, new_AGEMA_signal_6700, add_sub1_1_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_7043, new_AGEMA_signal_7042, add_sub1_1_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_6703, new_AGEMA_signal_6702, add_sub1_1_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_6133, new_AGEMA_signal_6132, addc_in[66]}), .c ({new_AGEMA_signal_7045, new_AGEMA_signal_7044, add_sub1_1_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_6691, new_AGEMA_signal_6690, add_sub1_1_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_7047, new_AGEMA_signal_7046, add_sub1_1_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_7279, new_AGEMA_signal_7278, subc_out[64]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_6695, new_AGEMA_signal_6694, add_sub1_1_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_6121, new_AGEMA_signal_6120, addc_in[64]}), .c ({new_AGEMA_signal_7047, new_AGEMA_signal_7046, add_sub1_1_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, addc_in[65]}), .b ({new_AGEMA_signal_6133, new_AGEMA_signal_6132, addc_in[66]}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_6695, new_AGEMA_signal_6694, add_sub1_1_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, addc_in[65]}), .b ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, addc_in[67]}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_6697, new_AGEMA_signal_6696, add_sub1_1_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6133, new_AGEMA_signal_6132, addc_in[66]}), .b ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, addc_in[67]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, add_sub1_1_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6121, new_AGEMA_signal_6120, addc_in[64]}), .b ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, addc_in[67]}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_6701, new_AGEMA_signal_6700, add_sub1_1_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6121, new_AGEMA_signal_6120, addc_in[64]}), .b ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, addc_in[65]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_6703, new_AGEMA_signal_6702, add_sub1_1_subc_rom_sbox_0_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_8667, new_AGEMA_signal_8666, add_sub1_2_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_8665, new_AGEMA_signal_8664, add_sub1_2_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_8833, new_AGEMA_signal_8832, add_sub1_2_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_8095, new_AGEMA_signal_8094, add_sub1_2_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_8099, new_AGEMA_signal_8098, add_sub1_2_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_8665, new_AGEMA_signal_8664, add_sub1_2_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_8101, new_AGEMA_signal_8100, add_sub1_2_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_7579, new_AGEMA_signal_7578, add_sub1_2_addc_out[2]}), .c ({new_AGEMA_signal_8667, new_AGEMA_signal_8666, add_sub1_2_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_8089, new_AGEMA_signal_8088, add_sub1_2_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_8669, new_AGEMA_signal_8668, add_sub1_2_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_8837, new_AGEMA_signal_8836, subc_out[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_8093, new_AGEMA_signal_8092, add_sub1_2_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_7583, new_AGEMA_signal_7582, add_sub1_2_addc_out[0]}), .c ({new_AGEMA_signal_8669, new_AGEMA_signal_8668, add_sub1_2_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_7581, new_AGEMA_signal_7580, add_sub1_2_addc_out[1]}), .b ({new_AGEMA_signal_7579, new_AGEMA_signal_7578, add_sub1_2_addc_out[2]}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_8093, new_AGEMA_signal_8092, add_sub1_2_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_7581, new_AGEMA_signal_7580, add_sub1_2_addc_out[1]}), .b ({new_AGEMA_signal_7577, new_AGEMA_signal_7576, add_sub1_2_addc_out[3]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_8095, new_AGEMA_signal_8094, add_sub1_2_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_7579, new_AGEMA_signal_7578, add_sub1_2_addc_out[2]}), .b ({new_AGEMA_signal_7577, new_AGEMA_signal_7576, add_sub1_2_addc_out[3]}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_8097, new_AGEMA_signal_8096, add_sub1_2_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_7583, new_AGEMA_signal_7582, add_sub1_2_addc_out[0]}), .b ({new_AGEMA_signal_7577, new_AGEMA_signal_7576, add_sub1_2_addc_out[3]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_8099, new_AGEMA_signal_8098, add_sub1_2_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_7583, new_AGEMA_signal_7582, add_sub1_2_addc_out[0]}), .b ({new_AGEMA_signal_7581, new_AGEMA_signal_7580, add_sub1_2_addc_out[1]}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_8101, new_AGEMA_signal_8100, add_sub1_2_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_7057, new_AGEMA_signal_7056, add_sub1_2_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_7055, new_AGEMA_signal_7054, add_sub1_2_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_7281, new_AGEMA_signal_7280, add_sub1_2_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_6715, new_AGEMA_signal_6714, add_sub1_2_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_6719, new_AGEMA_signal_6718, add_sub1_2_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_7055, new_AGEMA_signal_7054, add_sub1_2_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_6721, new_AGEMA_signal_6720, add_sub1_2_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_6085, new_AGEMA_signal_6084, addc_in[58]}), .c ({new_AGEMA_signal_7057, new_AGEMA_signal_7056, add_sub1_2_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_6709, new_AGEMA_signal_6708, add_sub1_2_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, add_sub1_2_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_7285, new_AGEMA_signal_7284, subc_out[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_6713, new_AGEMA_signal_6712, add_sub1_2_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, addc_in[56]}), .c ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, add_sub1_2_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, addc_in[57]}), .b ({new_AGEMA_signal_6085, new_AGEMA_signal_6084, addc_in[58]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_6713, new_AGEMA_signal_6712, add_sub1_2_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, addc_in[57]}), .b ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, addc_in[59]}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_6715, new_AGEMA_signal_6714, add_sub1_2_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6085, new_AGEMA_signal_6084, addc_in[58]}), .b ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, addc_in[59]}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_6717, new_AGEMA_signal_6716, add_sub1_2_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, addc_in[56]}), .b ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, addc_in[59]}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_6719, new_AGEMA_signal_6718, add_sub1_2_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, addc_in[56]}), .b ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, addc_in[57]}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_6721, new_AGEMA_signal_6720, add_sub1_2_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_7067, new_AGEMA_signal_7066, add_sub1_2_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, add_sub1_2_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_7287, new_AGEMA_signal_7286, add_sub1_2_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, add_sub1_2_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_6733, new_AGEMA_signal_6732, add_sub1_2_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, add_sub1_2_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, add_sub1_2_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, addc_in[54]}), .c ({new_AGEMA_signal_7067, new_AGEMA_signal_7066, add_sub1_2_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, add_sub1_2_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_7069, new_AGEMA_signal_7068, add_sub1_2_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_7291, new_AGEMA_signal_7290, subc_out[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_6727, new_AGEMA_signal_6726, add_sub1_2_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_6049, new_AGEMA_signal_6048, addc_in[52]}), .c ({new_AGEMA_signal_7069, new_AGEMA_signal_7068, add_sub1_2_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, addc_in[53]}), .b ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, addc_in[54]}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_6727, new_AGEMA_signal_6726, add_sub1_2_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, addc_in[53]}), .b ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, addc_in[55]}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, add_sub1_2_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, addc_in[54]}), .b ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, addc_in[55]}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_6731, new_AGEMA_signal_6730, add_sub1_2_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6049, new_AGEMA_signal_6048, addc_in[52]}), .b ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, addc_in[55]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_6733, new_AGEMA_signal_6732, add_sub1_2_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6049, new_AGEMA_signal_6048, addc_in[52]}), .b ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, addc_in[53]}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, add_sub1_2_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_7077, new_AGEMA_signal_7076, add_sub1_2_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_7075, new_AGEMA_signal_7074, add_sub1_2_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, add_sub1_2_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_6743, new_AGEMA_signal_6742, add_sub1_2_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, add_sub1_2_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_7075, new_AGEMA_signal_7074, add_sub1_2_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_6749, new_AGEMA_signal_6748, add_sub1_2_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, addc_in[50]}), .c ({new_AGEMA_signal_7077, new_AGEMA_signal_7076, add_sub1_2_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_6737, new_AGEMA_signal_6736, add_sub1_2_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_7079, new_AGEMA_signal_7078, add_sub1_2_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_7297, new_AGEMA_signal_7296, subc_out[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, add_sub1_2_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_6025, new_AGEMA_signal_6024, addc_in[48]}), .c ({new_AGEMA_signal_7079, new_AGEMA_signal_7078, add_sub1_2_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, addc_in[49]}), .b ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, addc_in[50]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, add_sub1_2_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, addc_in[49]}), .b ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, addc_in[51]}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_6743, new_AGEMA_signal_6742, add_sub1_2_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, addc_in[50]}), .b ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, addc_in[51]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_6745, new_AGEMA_signal_6744, add_sub1_2_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6025, new_AGEMA_signal_6024, addc_in[48]}), .b ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, addc_in[51]}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, add_sub1_2_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6025, new_AGEMA_signal_6024, addc_in[48]}), .b ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, addc_in[49]}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_6749, new_AGEMA_signal_6748, add_sub1_2_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_7087, new_AGEMA_signal_7086, add_sub1_2_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_7085, new_AGEMA_signal_7084, add_sub1_2_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, add_sub1_2_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_6757, new_AGEMA_signal_6756, add_sub1_2_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_6761, new_AGEMA_signal_6760, add_sub1_2_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_7085, new_AGEMA_signal_7084, add_sub1_2_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_6763, new_AGEMA_signal_6762, add_sub1_2_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_6013, new_AGEMA_signal_6012, addc_in[46]}), .c ({new_AGEMA_signal_7087, new_AGEMA_signal_7086, add_sub1_2_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_6751, new_AGEMA_signal_6750, add_sub1_2_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, add_sub1_2_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_7303, new_AGEMA_signal_7302, subc_out[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_6755, new_AGEMA_signal_6754, add_sub1_2_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_6001, new_AGEMA_signal_6000, addc_in[44]}), .c ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, add_sub1_2_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, addc_in[45]}), .b ({new_AGEMA_signal_6013, new_AGEMA_signal_6012, addc_in[46]}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_6755, new_AGEMA_signal_6754, add_sub1_2_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, addc_in[45]}), .b ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, addc_in[47]}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_6757, new_AGEMA_signal_6756, add_sub1_2_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6013, new_AGEMA_signal_6012, addc_in[46]}), .b ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, addc_in[47]}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, add_sub1_2_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6001, new_AGEMA_signal_6000, addc_in[44]}), .b ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, addc_in[47]}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_6761, new_AGEMA_signal_6760, add_sub1_2_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6001, new_AGEMA_signal_6000, addc_in[44]}), .b ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, addc_in[45]}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_6763, new_AGEMA_signal_6762, add_sub1_2_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_7097, new_AGEMA_signal_7096, add_sub1_2_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_7095, new_AGEMA_signal_7094, add_sub1_2_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_7305, new_AGEMA_signal_7304, add_sub1_2_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, add_sub1_2_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_6775, new_AGEMA_signal_6774, add_sub1_2_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_7095, new_AGEMA_signal_7094, add_sub1_2_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, add_sub1_2_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_5989, new_AGEMA_signal_5988, addc_in[42]}), .c ({new_AGEMA_signal_7097, new_AGEMA_signal_7096, add_sub1_2_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_6765, new_AGEMA_signal_6764, add_sub1_2_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_7099, new_AGEMA_signal_7098, add_sub1_2_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_7309, new_AGEMA_signal_7308, subc_out[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_6769, new_AGEMA_signal_6768, add_sub1_2_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_5977, new_AGEMA_signal_5976, addc_in[40]}), .c ({new_AGEMA_signal_7099, new_AGEMA_signal_7098, add_sub1_2_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, addc_in[41]}), .b ({new_AGEMA_signal_5989, new_AGEMA_signal_5988, addc_in[42]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_6769, new_AGEMA_signal_6768, add_sub1_2_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, addc_in[41]}), .b ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, addc_in[43]}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, add_sub1_2_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5989, new_AGEMA_signal_5988, addc_in[42]}), .b ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, addc_in[43]}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_6773, new_AGEMA_signal_6772, add_sub1_2_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5977, new_AGEMA_signal_5976, addc_in[40]}), .b ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, addc_in[43]}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_6775, new_AGEMA_signal_6774, add_sub1_2_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5977, new_AGEMA_signal_5976, addc_in[40]}), .b ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, addc_in[41]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, add_sub1_2_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, add_sub1_2_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_7105, new_AGEMA_signal_7104, add_sub1_2_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_7311, new_AGEMA_signal_7310, add_sub1_2_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_6785, new_AGEMA_signal_6784, add_sub1_2_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_6789, new_AGEMA_signal_6788, add_sub1_2_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_7105, new_AGEMA_signal_7104, add_sub1_2_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_6791, new_AGEMA_signal_6790, add_sub1_2_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, addc_in[38]}), .c ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, add_sub1_2_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_6779, new_AGEMA_signal_6778, add_sub1_2_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_7109, new_AGEMA_signal_7108, add_sub1_2_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_7315, new_AGEMA_signal_7314, subc_out[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, add_sub1_2_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, addc_in[36]}), .c ({new_AGEMA_signal_7109, new_AGEMA_signal_7108, add_sub1_2_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, addc_in[37]}), .b ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, addc_in[38]}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, add_sub1_2_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, addc_in[37]}), .b ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, addc_in[39]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_6785, new_AGEMA_signal_6784, add_sub1_2_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, addc_in[38]}), .b ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, addc_in[39]}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_6787, new_AGEMA_signal_6786, add_sub1_2_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, addc_in[36]}), .b ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, addc_in[39]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_6789, new_AGEMA_signal_6788, add_sub1_2_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, addc_in[36]}), .b ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, addc_in[37]}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_6791, new_AGEMA_signal_6790, add_sub1_2_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_7117, new_AGEMA_signal_7116, add_sub1_2_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_7115, new_AGEMA_signal_7114, add_sub1_2_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_7317, new_AGEMA_signal_7316, add_sub1_2_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_6799, new_AGEMA_signal_6798, add_sub1_2_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_6803, new_AGEMA_signal_6802, add_sub1_2_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_7115, new_AGEMA_signal_7114, add_sub1_2_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_6805, new_AGEMA_signal_6804, add_sub1_2_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, addc_in[34]}), .c ({new_AGEMA_signal_7117, new_AGEMA_signal_7116, add_sub1_2_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_6793, new_AGEMA_signal_6792, add_sub1_2_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_7119, new_AGEMA_signal_7118, add_sub1_2_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_7321, new_AGEMA_signal_7320, subc_out[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_6797, new_AGEMA_signal_6796, add_sub1_2_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, addc_in[32]}), .c ({new_AGEMA_signal_7119, new_AGEMA_signal_7118, add_sub1_2_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, addc_in[33]}), .b ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, addc_in[34]}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_6797, new_AGEMA_signal_6796, add_sub1_2_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, addc_in[33]}), .b ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, addc_in[35]}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_6799, new_AGEMA_signal_6798, add_sub1_2_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, addc_in[34]}), .b ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, addc_in[35]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_6801, new_AGEMA_signal_6800, add_sub1_2_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, addc_in[32]}), .b ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, addc_in[35]}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_6803, new_AGEMA_signal_6802, add_sub1_2_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, addc_in[32]}), .b ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, addc_in[33]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_6805, new_AGEMA_signal_6804, add_sub1_2_subc_rom_sbox_0_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_8691, new_AGEMA_signal_8690, add_sub1_3_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_8689, new_AGEMA_signal_8688, add_sub1_3_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_8839, new_AGEMA_signal_8838, add_sub1_3_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_8137, new_AGEMA_signal_8136, add_sub1_3_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_8141, new_AGEMA_signal_8140, add_sub1_3_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_8689, new_AGEMA_signal_8688, add_sub1_3_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_8143, new_AGEMA_signal_8142, add_sub1_3_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_7601, new_AGEMA_signal_7600, add_sub1_3_addc_out[2]}), .c ({new_AGEMA_signal_8691, new_AGEMA_signal_8690, add_sub1_3_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_8131, new_AGEMA_signal_8130, add_sub1_3_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_8693, new_AGEMA_signal_8692, add_sub1_3_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_8843, new_AGEMA_signal_8842, subc_out[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_8135, new_AGEMA_signal_8134, add_sub1_3_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_7605, new_AGEMA_signal_7604, add_sub1_3_addc_out[0]}), .c ({new_AGEMA_signal_8693, new_AGEMA_signal_8692, add_sub1_3_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_7603, new_AGEMA_signal_7602, add_sub1_3_addc_out[1]}), .b ({new_AGEMA_signal_7601, new_AGEMA_signal_7600, add_sub1_3_addc_out[2]}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_8135, new_AGEMA_signal_8134, add_sub1_3_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_7603, new_AGEMA_signal_7602, add_sub1_3_addc_out[1]}), .b ({new_AGEMA_signal_7599, new_AGEMA_signal_7598, add_sub1_3_addc_out[3]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_8137, new_AGEMA_signal_8136, add_sub1_3_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_7601, new_AGEMA_signal_7600, add_sub1_3_addc_out[2]}), .b ({new_AGEMA_signal_7599, new_AGEMA_signal_7598, add_sub1_3_addc_out[3]}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_8139, new_AGEMA_signal_8138, add_sub1_3_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_7605, new_AGEMA_signal_7604, add_sub1_3_addc_out[0]}), .b ({new_AGEMA_signal_7599, new_AGEMA_signal_7598, add_sub1_3_addc_out[3]}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_8141, new_AGEMA_signal_8140, add_sub1_3_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_7605, new_AGEMA_signal_7604, add_sub1_3_addc_out[0]}), .b ({new_AGEMA_signal_7603, new_AGEMA_signal_7602, add_sub1_3_addc_out[1]}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_8143, new_AGEMA_signal_8142, add_sub1_3_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_7129, new_AGEMA_signal_7128, add_sub1_3_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_7127, new_AGEMA_signal_7126, add_sub1_3_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_7323, new_AGEMA_signal_7322, add_sub1_3_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_6817, new_AGEMA_signal_6816, add_sub1_3_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_6821, new_AGEMA_signal_6820, add_sub1_3_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_7127, new_AGEMA_signal_7126, add_sub1_3_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_6823, new_AGEMA_signal_6822, add_sub1_3_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, addc_in[26]}), .c ({new_AGEMA_signal_7129, new_AGEMA_signal_7128, add_sub1_3_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_6811, new_AGEMA_signal_6810, add_sub1_3_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_7131, new_AGEMA_signal_7130, add_sub1_3_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_7327, new_AGEMA_signal_7326, subc_out[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_6815, new_AGEMA_signal_6814, add_sub1_3_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_5881, new_AGEMA_signal_5880, addc_in[24]}), .c ({new_AGEMA_signal_7131, new_AGEMA_signal_7130, add_sub1_3_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, addc_in[25]}), .b ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, addc_in[26]}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_6815, new_AGEMA_signal_6814, add_sub1_3_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, addc_in[25]}), .b ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, addc_in[27]}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_6817, new_AGEMA_signal_6816, add_sub1_3_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, addc_in[26]}), .b ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, addc_in[27]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_6819, new_AGEMA_signal_6818, add_sub1_3_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5881, new_AGEMA_signal_5880, addc_in[24]}), .b ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, addc_in[27]}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_6821, new_AGEMA_signal_6820, add_sub1_3_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5881, new_AGEMA_signal_5880, addc_in[24]}), .b ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, addc_in[25]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_6823, new_AGEMA_signal_6822, add_sub1_3_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_7139, new_AGEMA_signal_7138, add_sub1_3_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, add_sub1_3_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_7329, new_AGEMA_signal_7328, add_sub1_3_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, add_sub1_3_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_6835, new_AGEMA_signal_6834, add_sub1_3_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, add_sub1_3_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_6837, new_AGEMA_signal_6836, add_sub1_3_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_5869, new_AGEMA_signal_5868, addc_in[22]}), .c ({new_AGEMA_signal_7139, new_AGEMA_signal_7138, add_sub1_3_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, add_sub1_3_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_7141, new_AGEMA_signal_7140, add_sub1_3_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_7333, new_AGEMA_signal_7332, subc_out[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_6829, new_AGEMA_signal_6828, add_sub1_3_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, addc_in[20]}), .c ({new_AGEMA_signal_7141, new_AGEMA_signal_7140, add_sub1_3_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, addc_in[21]}), .b ({new_AGEMA_signal_5869, new_AGEMA_signal_5868, addc_in[22]}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_6829, new_AGEMA_signal_6828, add_sub1_3_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, addc_in[21]}), .b ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, addc_in[23]}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, add_sub1_3_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5869, new_AGEMA_signal_5868, addc_in[22]}), .b ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, addc_in[23]}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_6833, new_AGEMA_signal_6832, add_sub1_3_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, addc_in[20]}), .b ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, addc_in[23]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_6835, new_AGEMA_signal_6834, add_sub1_3_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, addc_in[20]}), .b ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, addc_in[21]}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_6837, new_AGEMA_signal_6836, add_sub1_3_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_7149, new_AGEMA_signal_7148, add_sub1_3_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_7147, new_AGEMA_signal_7146, add_sub1_3_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_7335, new_AGEMA_signal_7334, add_sub1_3_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_6845, new_AGEMA_signal_6844, add_sub1_3_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, add_sub1_3_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_7147, new_AGEMA_signal_7146, add_sub1_3_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_6851, new_AGEMA_signal_6850, add_sub1_3_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_5845, new_AGEMA_signal_5844, addc_in[18]}), .c ({new_AGEMA_signal_7149, new_AGEMA_signal_7148, add_sub1_3_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_6839, new_AGEMA_signal_6838, add_sub1_3_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_7151, new_AGEMA_signal_7150, add_sub1_3_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_7339, new_AGEMA_signal_7338, subc_out[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, add_sub1_3_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_5833, new_AGEMA_signal_5832, addc_in[16]}), .c ({new_AGEMA_signal_7151, new_AGEMA_signal_7150, add_sub1_3_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, addc_in[17]}), .b ({new_AGEMA_signal_5845, new_AGEMA_signal_5844, addc_in[18]}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, add_sub1_3_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, addc_in[17]}), .b ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, addc_in[19]}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_6845, new_AGEMA_signal_6844, add_sub1_3_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5845, new_AGEMA_signal_5844, addc_in[18]}), .b ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, addc_in[19]}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_6847, new_AGEMA_signal_6846, add_sub1_3_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5833, new_AGEMA_signal_5832, addc_in[16]}), .b ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, addc_in[19]}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, add_sub1_3_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5833, new_AGEMA_signal_5832, addc_in[16]}), .b ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, addc_in[17]}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_6851, new_AGEMA_signal_6850, add_sub1_3_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_7159, new_AGEMA_signal_7158, add_sub1_3_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_7157, new_AGEMA_signal_7156, add_sub1_3_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, add_sub1_3_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_6859, new_AGEMA_signal_6858, add_sub1_3_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_6863, new_AGEMA_signal_6862, add_sub1_3_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_7157, new_AGEMA_signal_7156, add_sub1_3_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_6865, new_AGEMA_signal_6864, add_sub1_3_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, addc_in[14]}), .c ({new_AGEMA_signal_7159, new_AGEMA_signal_7158, add_sub1_3_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_6853, new_AGEMA_signal_6852, add_sub1_3_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, add_sub1_3_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_7345, new_AGEMA_signal_7344, subc_out[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_6857, new_AGEMA_signal_6856, add_sub1_3_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_5809, new_AGEMA_signal_5808, addc_in[12]}), .c ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, add_sub1_3_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, addc_in[13]}), .b ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, addc_in[14]}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_6857, new_AGEMA_signal_6856, add_sub1_3_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, addc_in[13]}), .b ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, addc_in[15]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_6859, new_AGEMA_signal_6858, add_sub1_3_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, addc_in[14]}), .b ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, addc_in[15]}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_6861, new_AGEMA_signal_6860, add_sub1_3_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5809, new_AGEMA_signal_5808, addc_in[12]}), .b ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, addc_in[15]}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_6863, new_AGEMA_signal_6862, add_sub1_3_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5809, new_AGEMA_signal_5808, addc_in[12]}), .b ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, addc_in[13]}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_6865, new_AGEMA_signal_6864, add_sub1_3_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_7169, new_AGEMA_signal_7168, add_sub1_3_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_7167, new_AGEMA_signal_7166, add_sub1_3_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_7347, new_AGEMA_signal_7346, add_sub1_3_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, add_sub1_3_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_6877, new_AGEMA_signal_6876, add_sub1_3_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_7167, new_AGEMA_signal_7166, add_sub1_3_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_6879, new_AGEMA_signal_6878, add_sub1_3_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_5797, new_AGEMA_signal_5796, addc_in[10]}), .c ({new_AGEMA_signal_7169, new_AGEMA_signal_7168, add_sub1_3_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_6867, new_AGEMA_signal_6866, add_sub1_3_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_7171, new_AGEMA_signal_7170, add_sub1_3_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_7351, new_AGEMA_signal_7350, subc_out[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_6871, new_AGEMA_signal_6870, add_sub1_3_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, addc_in[8]}), .c ({new_AGEMA_signal_7171, new_AGEMA_signal_7170, add_sub1_3_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, addc_in[9]}), .b ({new_AGEMA_signal_5797, new_AGEMA_signal_5796, addc_in[10]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_6871, new_AGEMA_signal_6870, add_sub1_3_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, addc_in[9]}), .b ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, addc_in[11]}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, add_sub1_3_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5797, new_AGEMA_signal_5796, addc_in[10]}), .b ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, addc_in[11]}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_6875, new_AGEMA_signal_6874, add_sub1_3_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, addc_in[8]}), .b ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, addc_in[11]}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_6877, new_AGEMA_signal_6876, add_sub1_3_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, addc_in[8]}), .b ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, addc_in[9]}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_6879, new_AGEMA_signal_6878, add_sub1_3_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_7179, new_AGEMA_signal_7178, add_sub1_3_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_7177, new_AGEMA_signal_7176, add_sub1_3_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_7353, new_AGEMA_signal_7352, add_sub1_3_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_6887, new_AGEMA_signal_6886, add_sub1_3_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_6891, new_AGEMA_signal_6890, add_sub1_3_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_7177, new_AGEMA_signal_7176, add_sub1_3_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_6893, new_AGEMA_signal_6892, add_sub1_3_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_5773, new_AGEMA_signal_5772, addc_in[6]}), .c ({new_AGEMA_signal_7179, new_AGEMA_signal_7178, add_sub1_3_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_6881, new_AGEMA_signal_6880, add_sub1_3_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_7181, new_AGEMA_signal_7180, add_sub1_3_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_7357, new_AGEMA_signal_7356, subc_out[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_6885, new_AGEMA_signal_6884, add_sub1_3_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, addc_in[4]}), .c ({new_AGEMA_signal_7181, new_AGEMA_signal_7180, add_sub1_3_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, addc_in[5]}), .b ({new_AGEMA_signal_5773, new_AGEMA_signal_5772, addc_in[6]}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_6885, new_AGEMA_signal_6884, add_sub1_3_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, addc_in[5]}), .b ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, addc_in[7]}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_6887, new_AGEMA_signal_6886, add_sub1_3_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5773, new_AGEMA_signal_5772, addc_in[6]}), .b ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, addc_in[7]}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_6889, new_AGEMA_signal_6888, add_sub1_3_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, addc_in[4]}), .b ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, addc_in[7]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_6891, new_AGEMA_signal_6890, add_sub1_3_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, addc_in[4]}), .b ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, addc_in[5]}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_6893, new_AGEMA_signal_6892, add_sub1_3_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_7189, new_AGEMA_signal_7188, add_sub1_3_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_7187, new_AGEMA_signal_7186, add_sub1_3_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_7359, new_AGEMA_signal_7358, add_sub1_3_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_6901, new_AGEMA_signal_6900, add_sub1_3_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_6905, new_AGEMA_signal_6904, add_sub1_3_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_7187, new_AGEMA_signal_7186, add_sub1_3_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_6907, new_AGEMA_signal_6906, add_sub1_3_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, addc_in[2]}), .c ({new_AGEMA_signal_7189, new_AGEMA_signal_7188, add_sub1_3_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_6895, new_AGEMA_signal_6894, add_sub1_3_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_7191, new_AGEMA_signal_7190, add_sub1_3_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_7363, new_AGEMA_signal_7362, subc_out[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_6899, new_AGEMA_signal_6898, add_sub1_3_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, addc_in[0]}), .c ({new_AGEMA_signal_7191, new_AGEMA_signal_7190, add_sub1_3_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, addc_in[1]}), .b ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, addc_in[2]}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_6899, new_AGEMA_signal_6898, add_sub1_3_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, addc_in[1]}), .b ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, addc_in[3]}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_6901, new_AGEMA_signal_6900, add_sub1_3_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, addc_in[2]}), .b ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, addc_in[3]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, add_sub1_3_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, addc_in[0]}), .b ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, addc_in[3]}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_6905, new_AGEMA_signal_6904, add_sub1_3_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, addc_in[0]}), .b ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, addc_in[1]}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_6907, new_AGEMA_signal_6906, add_sub1_3_subc_rom_sbox_0_ANF_2_t7}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7237, new_AGEMA_signal_7236, subc_out[96]}), .a ({new_AGEMA_signal_7213, new_AGEMA_signal_7212, subc_out[112]}), .c ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7231, new_AGEMA_signal_7230, subc_out[100]}), .a ({new_AGEMA_signal_7207, new_AGEMA_signal_7206, subc_out[116]}), .c ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7225, new_AGEMA_signal_7224, subc_out[104]}), .a ({new_AGEMA_signal_7201, new_AGEMA_signal_7200, subc_out[120]}), .c ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7219, new_AGEMA_signal_7218, subc_out[108]}), .a ({new_AGEMA_signal_8825, new_AGEMA_signal_8824, subc_out[124]}), .c ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7213, new_AGEMA_signal_7212, subc_out[112]}), .a ({new_AGEMA_signal_7237, new_AGEMA_signal_7236, subc_out[96]}), .c ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7207, new_AGEMA_signal_7206, subc_out[116]}), .a ({new_AGEMA_signal_7231, new_AGEMA_signal_7230, subc_out[100]}), .c ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7201, new_AGEMA_signal_7200, subc_out[120]}), .a ({new_AGEMA_signal_7225, new_AGEMA_signal_7224, subc_out[104]}), .c ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8825, new_AGEMA_signal_8824, subc_out[124]}), .a ({new_AGEMA_signal_7219, new_AGEMA_signal_7218, subc_out[108]}), .c ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8831, new_AGEMA_signal_8830, subc_out[92]}), .a ({new_AGEMA_signal_7261, new_AGEMA_signal_7260, subc_out[76]}), .c ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7279, new_AGEMA_signal_7278, subc_out[64]}), .a ({new_AGEMA_signal_7255, new_AGEMA_signal_7254, subc_out[80]}), .c ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7273, new_AGEMA_signal_7272, subc_out[68]}), .a ({new_AGEMA_signal_7249, new_AGEMA_signal_7248, subc_out[84]}), .c ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7267, new_AGEMA_signal_7266, subc_out[72]}), .a ({new_AGEMA_signal_7243, new_AGEMA_signal_7242, subc_out[88]}), .c ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7261, new_AGEMA_signal_7260, subc_out[76]}), .a ({new_AGEMA_signal_8831, new_AGEMA_signal_8830, subc_out[92]}), .c ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7255, new_AGEMA_signal_7254, subc_out[80]}), .a ({new_AGEMA_signal_7279, new_AGEMA_signal_7278, subc_out[64]}), .c ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7249, new_AGEMA_signal_7248, subc_out[84]}), .a ({new_AGEMA_signal_7273, new_AGEMA_signal_7272, subc_out[68]}), .c ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7243, new_AGEMA_signal_7242, subc_out[88]}), .a ({new_AGEMA_signal_7267, new_AGEMA_signal_7266, subc_out[72]}), .c ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7285, new_AGEMA_signal_7284, subc_out[56]}), .a ({new_AGEMA_signal_7309, new_AGEMA_signal_7308, subc_out[40]}), .c ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8837, new_AGEMA_signal_8836, subc_out[60]}), .a ({new_AGEMA_signal_7303, new_AGEMA_signal_7302, subc_out[44]}), .c ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7321, new_AGEMA_signal_7320, subc_out[32]}), .a ({new_AGEMA_signal_7297, new_AGEMA_signal_7296, subc_out[48]}), .c ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7315, new_AGEMA_signal_7314, subc_out[36]}), .a ({new_AGEMA_signal_7291, new_AGEMA_signal_7290, subc_out[52]}), .c ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7309, new_AGEMA_signal_7308, subc_out[40]}), .a ({new_AGEMA_signal_7285, new_AGEMA_signal_7284, subc_out[56]}), .c ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7303, new_AGEMA_signal_7302, subc_out[44]}), .a ({new_AGEMA_signal_8837, new_AGEMA_signal_8836, subc_out[60]}), .c ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7297, new_AGEMA_signal_7296, subc_out[48]}), .a ({new_AGEMA_signal_7321, new_AGEMA_signal_7320, subc_out[32]}), .c ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7291, new_AGEMA_signal_7290, subc_out[52]}), .a ({new_AGEMA_signal_7315, new_AGEMA_signal_7314, subc_out[36]}), .c ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7333, new_AGEMA_signal_7332, subc_out[20]}), .a ({new_AGEMA_signal_7357, new_AGEMA_signal_7356, subc_out[4]}), .c ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7327, new_AGEMA_signal_7326, subc_out[24]}), .a ({new_AGEMA_signal_7351, new_AGEMA_signal_7350, subc_out[8]}), .c ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8843, new_AGEMA_signal_8842, subc_out[28]}), .a ({new_AGEMA_signal_7345, new_AGEMA_signal_7344, subc_out[12]}), .c ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7363, new_AGEMA_signal_7362, subc_out[0]}), .a ({new_AGEMA_signal_7339, new_AGEMA_signal_7338, subc_out[16]}), .c ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7357, new_AGEMA_signal_7356, subc_out[4]}), .a ({new_AGEMA_signal_7333, new_AGEMA_signal_7332, subc_out[20]}), .c ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7351, new_AGEMA_signal_7350, subc_out[8]}), .a ({new_AGEMA_signal_7327, new_AGEMA_signal_7326, subc_out[24]}), .c ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7345, new_AGEMA_signal_7344, subc_out[12]}), .a ({new_AGEMA_signal_8843, new_AGEMA_signal_8842, subc_out[28]}), .c ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7339, new_AGEMA_signal_7338, subc_out[16]}), .a ({new_AGEMA_signal_7363, new_AGEMA_signal_7362, subc_out[0]}), .c ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_10449, new_AGEMA_signal_10448, add_sub1_0_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_8621, new_AGEMA_signal_8620, add_sub1_0_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_11413, new_AGEMA_signal_11412, subc_out[127]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, add_sub1_0_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_8821, new_AGEMA_signal_8820, add_sub1_0_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_9481, new_AGEMA_signal_9480, subc_out[126]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_11415, new_AGEMA_signal_11414, add_sub1_0_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_8013, new_AGEMA_signal_8012, add_sub1_0_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_12365, new_AGEMA_signal_12364, subc_out[125]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_10449, new_AGEMA_signal_10448, add_sub1_0_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_8011, new_AGEMA_signal_8010, add_sub1_0_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_11415, new_AGEMA_signal_11414, add_sub1_0_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, add_sub1_0_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_7537, new_AGEMA_signal_7536, add_sub1_0_addc_out[1]}), .c ({new_AGEMA_signal_10449, new_AGEMA_signal_10448, add_sub1_0_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, add_sub1_0_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, add_sub1_0_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, add_sub1_0_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_8625, new_AGEMA_signal_8624, add_sub1_0_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, add_sub1_0_addc_out[3]}), .c ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, add_sub1_0_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_7539, new_AGEMA_signal_7538, add_sub1_0_addc_out[0]}), .b ({new_AGEMA_signal_8009, new_AGEMA_signal_8008, add_sub1_0_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, add_sub1_0_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_8007, new_AGEMA_signal_8006, add_sub1_0_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_8015, new_AGEMA_signal_8014, add_sub1_0_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_8625, new_AGEMA_signal_8624, add_sub1_0_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_7541, new_AGEMA_signal_7540, add_sub1_0_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6915, new_AGEMA_signal_6914, add_sub1_0_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_8019, new_AGEMA_signal_8018, subc_out[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_7199, new_AGEMA_signal_7198, add_sub1_0_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7197, new_AGEMA_signal_7196, add_sub1_0_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_7367, new_AGEMA_signal_7366, subc_out[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_8021, new_AGEMA_signal_8020, add_sub1_0_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, add_sub1_0_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_8627, new_AGEMA_signal_8626, subc_out[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_7541, new_AGEMA_signal_7540, add_sub1_0_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6511, new_AGEMA_signal_6510, add_sub1_0_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_8021, new_AGEMA_signal_8020, add_sub1_0_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_7369, new_AGEMA_signal_7368, add_sub1_0_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_6463, new_AGEMA_signal_6462, addc_in[121]}), .c ({new_AGEMA_signal_7541, new_AGEMA_signal_7540, add_sub1_0_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_7199, new_AGEMA_signal_7198, add_sub1_0_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_6917, new_AGEMA_signal_6916, add_sub1_0_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_7369, new_AGEMA_signal_7368, add_sub1_0_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_6919, new_AGEMA_signal_6918, add_sub1_0_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_6475, new_AGEMA_signal_6474, addc_in[123]}), .c ({new_AGEMA_signal_7199, new_AGEMA_signal_7198, add_sub1_0_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6457, new_AGEMA_signal_6456, addc_in[120]}), .b ({new_AGEMA_signal_6509, new_AGEMA_signal_6508, add_sub1_0_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_6917, new_AGEMA_signal_6916, add_sub1_0_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, add_sub1_0_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_6515, new_AGEMA_signal_6514, add_sub1_0_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_6919, new_AGEMA_signal_6918, add_sub1_0_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_7543, new_AGEMA_signal_7542, add_sub1_0_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6925, new_AGEMA_signal_6924, add_sub1_0_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_8023, new_AGEMA_signal_8022, subc_out[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_7205, new_AGEMA_signal_7204, add_sub1_0_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7203, new_AGEMA_signal_7202, add_sub1_0_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, subc_out[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_8025, new_AGEMA_signal_8024, add_sub1_0_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_6527, new_AGEMA_signal_6526, add_sub1_0_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, subc_out[117]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_7543, new_AGEMA_signal_7542, add_sub1_0_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6525, new_AGEMA_signal_6524, add_sub1_0_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_8025, new_AGEMA_signal_8024, add_sub1_0_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_7373, new_AGEMA_signal_7372, add_sub1_0_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_6439, new_AGEMA_signal_6438, addc_in[117]}), .c ({new_AGEMA_signal_7543, new_AGEMA_signal_7542, add_sub1_0_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_7205, new_AGEMA_signal_7204, add_sub1_0_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_6927, new_AGEMA_signal_6926, add_sub1_0_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_7373, new_AGEMA_signal_7372, add_sub1_0_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_6929, new_AGEMA_signal_6928, add_sub1_0_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, addc_in[119]}), .c ({new_AGEMA_signal_7205, new_AGEMA_signal_7204, add_sub1_0_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, addc_in[116]}), .b ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, add_sub1_0_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_6927, new_AGEMA_signal_6926, add_sub1_0_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6521, new_AGEMA_signal_6520, add_sub1_0_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_6529, new_AGEMA_signal_6528, add_sub1_0_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_6929, new_AGEMA_signal_6928, add_sub1_0_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_7545, new_AGEMA_signal_7544, add_sub1_0_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6935, new_AGEMA_signal_6934, add_sub1_0_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_8027, new_AGEMA_signal_8026, subc_out[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_7211, new_AGEMA_signal_7210, add_sub1_0_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7209, new_AGEMA_signal_7208, add_sub1_0_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_7375, new_AGEMA_signal_7374, subc_out[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_8029, new_AGEMA_signal_8028, add_sub1_0_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_6541, new_AGEMA_signal_6540, add_sub1_0_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_8631, new_AGEMA_signal_8630, subc_out[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_7545, new_AGEMA_signal_7544, add_sub1_0_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6539, new_AGEMA_signal_6538, add_sub1_0_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_8029, new_AGEMA_signal_8028, add_sub1_0_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, add_sub1_0_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, addc_in[113]}), .c ({new_AGEMA_signal_7545, new_AGEMA_signal_7544, add_sub1_0_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_7211, new_AGEMA_signal_7210, add_sub1_0_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_6937, new_AGEMA_signal_6936, add_sub1_0_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, add_sub1_0_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_6939, new_AGEMA_signal_6938, add_sub1_0_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_6427, new_AGEMA_signal_6426, addc_in[115]}), .c ({new_AGEMA_signal_7211, new_AGEMA_signal_7210, add_sub1_0_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6409, new_AGEMA_signal_6408, addc_in[112]}), .b ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, add_sub1_0_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_6937, new_AGEMA_signal_6936, add_sub1_0_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6535, new_AGEMA_signal_6534, add_sub1_0_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, add_sub1_0_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_6939, new_AGEMA_signal_6938, add_sub1_0_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_7547, new_AGEMA_signal_7546, add_sub1_0_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6945, new_AGEMA_signal_6944, add_sub1_0_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_8031, new_AGEMA_signal_8030, subc_out[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_7217, new_AGEMA_signal_7216, add_sub1_0_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, add_sub1_0_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_7379, new_AGEMA_signal_7378, subc_out[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_8033, new_AGEMA_signal_8032, add_sub1_0_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, add_sub1_0_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_8633, new_AGEMA_signal_8632, subc_out[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_7547, new_AGEMA_signal_7546, add_sub1_0_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6553, new_AGEMA_signal_6552, add_sub1_0_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_8033, new_AGEMA_signal_8032, add_sub1_0_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_7381, new_AGEMA_signal_7380, add_sub1_0_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_6391, new_AGEMA_signal_6390, addc_in[109]}), .c ({new_AGEMA_signal_7547, new_AGEMA_signal_7546, add_sub1_0_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_7217, new_AGEMA_signal_7216, add_sub1_0_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_6947, new_AGEMA_signal_6946, add_sub1_0_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_7381, new_AGEMA_signal_7380, add_sub1_0_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_6949, new_AGEMA_signal_6948, add_sub1_0_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_6403, new_AGEMA_signal_6402, addc_in[111]}), .c ({new_AGEMA_signal_7217, new_AGEMA_signal_7216, add_sub1_0_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6385, new_AGEMA_signal_6384, addc_in[108]}), .b ({new_AGEMA_signal_6551, new_AGEMA_signal_6550, add_sub1_0_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_6947, new_AGEMA_signal_6946, add_sub1_0_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6549, new_AGEMA_signal_6548, add_sub1_0_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_6557, new_AGEMA_signal_6556, add_sub1_0_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_6949, new_AGEMA_signal_6948, add_sub1_0_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_7549, new_AGEMA_signal_7548, add_sub1_0_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6955, new_AGEMA_signal_6954, add_sub1_0_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_8035, new_AGEMA_signal_8034, subc_out[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_7223, new_AGEMA_signal_7222, add_sub1_0_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, add_sub1_0_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_7383, new_AGEMA_signal_7382, subc_out[106]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_8037, new_AGEMA_signal_8036, add_sub1_0_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_6569, new_AGEMA_signal_6568, add_sub1_0_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, subc_out[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_7549, new_AGEMA_signal_7548, add_sub1_0_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, add_sub1_0_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_8037, new_AGEMA_signal_8036, add_sub1_0_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_7385, new_AGEMA_signal_7384, add_sub1_0_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_6367, new_AGEMA_signal_6366, addc_in[105]}), .c ({new_AGEMA_signal_7549, new_AGEMA_signal_7548, add_sub1_0_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_7223, new_AGEMA_signal_7222, add_sub1_0_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_6957, new_AGEMA_signal_6956, add_sub1_0_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_7385, new_AGEMA_signal_7384, add_sub1_0_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_6959, new_AGEMA_signal_6958, add_sub1_0_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, addc_in[107]}), .c ({new_AGEMA_signal_7223, new_AGEMA_signal_7222, add_sub1_0_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, addc_in[104]}), .b ({new_AGEMA_signal_6565, new_AGEMA_signal_6564, add_sub1_0_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_6957, new_AGEMA_signal_6956, add_sub1_0_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6563, new_AGEMA_signal_6562, add_sub1_0_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_6571, new_AGEMA_signal_6570, add_sub1_0_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_6959, new_AGEMA_signal_6958, add_sub1_0_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_7551, new_AGEMA_signal_7550, add_sub1_0_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6965, new_AGEMA_signal_6964, add_sub1_0_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_8039, new_AGEMA_signal_8038, subc_out[103]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_7229, new_AGEMA_signal_7228, add_sub1_0_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7227, new_AGEMA_signal_7226, add_sub1_0_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_7387, new_AGEMA_signal_7386, subc_out[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_8041, new_AGEMA_signal_8040, add_sub1_0_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_6583, new_AGEMA_signal_6582, add_sub1_0_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, subc_out[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_7551, new_AGEMA_signal_7550, add_sub1_0_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6581, new_AGEMA_signal_6580, add_sub1_0_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_8041, new_AGEMA_signal_8040, add_sub1_0_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_7389, new_AGEMA_signal_7388, add_sub1_0_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, addc_in[101]}), .c ({new_AGEMA_signal_7551, new_AGEMA_signal_7550, add_sub1_0_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_7229, new_AGEMA_signal_7228, add_sub1_0_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_6967, new_AGEMA_signal_6966, add_sub1_0_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_7389, new_AGEMA_signal_7388, add_sub1_0_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_6969, new_AGEMA_signal_6968, add_sub1_0_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_6355, new_AGEMA_signal_6354, addc_in[103]}), .c ({new_AGEMA_signal_7229, new_AGEMA_signal_7228, add_sub1_0_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6337, new_AGEMA_signal_6336, addc_in[100]}), .b ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, add_sub1_0_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_6967, new_AGEMA_signal_6966, add_sub1_0_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6577, new_AGEMA_signal_6576, add_sub1_0_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, add_sub1_0_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_6969, new_AGEMA_signal_6968, add_sub1_0_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_7553, new_AGEMA_signal_7552, add_sub1_0_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6975, new_AGEMA_signal_6974, add_sub1_0_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_8043, new_AGEMA_signal_8042, subc_out[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_7235, new_AGEMA_signal_7234, add_sub1_0_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, add_sub1_0_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_7391, new_AGEMA_signal_7390, subc_out[98]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_8045, new_AGEMA_signal_8044, add_sub1_0_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_6597, new_AGEMA_signal_6596, add_sub1_0_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_8639, new_AGEMA_signal_8638, subc_out[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_7553, new_AGEMA_signal_7552, add_sub1_0_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6595, new_AGEMA_signal_6594, add_sub1_0_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_8045, new_AGEMA_signal_8044, add_sub1_0_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_7393, new_AGEMA_signal_7392, add_sub1_0_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_6319, new_AGEMA_signal_6318, addc_in[97]}), .c ({new_AGEMA_signal_7553, new_AGEMA_signal_7552, add_sub1_0_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_7235, new_AGEMA_signal_7234, add_sub1_0_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_6977, new_AGEMA_signal_6976, add_sub1_0_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_7393, new_AGEMA_signal_7392, add_sub1_0_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_6979, new_AGEMA_signal_6978, add_sub1_0_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_6331, new_AGEMA_signal_6330, addc_in[99]}), .c ({new_AGEMA_signal_7235, new_AGEMA_signal_7234, add_sub1_0_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6313, new_AGEMA_signal_6312, addc_in[96]}), .b ({new_AGEMA_signal_6593, new_AGEMA_signal_6592, add_sub1_0_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_6977, new_AGEMA_signal_6976, add_sub1_0_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, add_sub1_0_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_6599, new_AGEMA_signal_6598, add_sub1_0_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_6979, new_AGEMA_signal_6978, add_sub1_0_subc_rom_sbox_0_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_10451, new_AGEMA_signal_10450, add_sub1_1_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_8645, new_AGEMA_signal_8644, add_sub1_1_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_11417, new_AGEMA_signal_11416, subc_out[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_8829, new_AGEMA_signal_8828, add_sub1_1_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_8827, new_AGEMA_signal_8826, add_sub1_1_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_9485, new_AGEMA_signal_9484, subc_out[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_11419, new_AGEMA_signal_11418, add_sub1_1_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_8055, new_AGEMA_signal_8054, add_sub1_1_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_12367, new_AGEMA_signal_12366, subc_out[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_10451, new_AGEMA_signal_10450, add_sub1_1_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_8053, new_AGEMA_signal_8052, add_sub1_1_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_11419, new_AGEMA_signal_11418, add_sub1_1_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_9487, new_AGEMA_signal_9486, add_sub1_1_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_7559, new_AGEMA_signal_7558, add_sub1_1_addc_out[1]}), .c ({new_AGEMA_signal_10451, new_AGEMA_signal_10450, add_sub1_1_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_8829, new_AGEMA_signal_8828, add_sub1_1_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_8647, new_AGEMA_signal_8646, add_sub1_1_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_9487, new_AGEMA_signal_9486, add_sub1_1_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_8649, new_AGEMA_signal_8648, add_sub1_1_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_7555, new_AGEMA_signal_7554, add_sub1_1_addc_out[3]}), .c ({new_AGEMA_signal_8829, new_AGEMA_signal_8828, add_sub1_1_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_7561, new_AGEMA_signal_7560, add_sub1_1_addc_out[0]}), .b ({new_AGEMA_signal_8051, new_AGEMA_signal_8050, add_sub1_1_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_8647, new_AGEMA_signal_8646, add_sub1_1_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_8049, new_AGEMA_signal_8048, add_sub1_1_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_8057, new_AGEMA_signal_8056, add_sub1_1_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_8649, new_AGEMA_signal_8648, add_sub1_1_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_7563, new_AGEMA_signal_7562, add_sub1_1_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, add_sub1_1_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_8061, new_AGEMA_signal_8060, subc_out[91]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_7241, new_AGEMA_signal_7240, add_sub1_1_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, add_sub1_1_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_7397, new_AGEMA_signal_7396, subc_out[90]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_8063, new_AGEMA_signal_8062, add_sub1_1_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, add_sub1_1_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_8651, new_AGEMA_signal_8650, subc_out[89]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_7563, new_AGEMA_signal_7562, add_sub1_1_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, add_sub1_1_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_8063, new_AGEMA_signal_8062, add_sub1_1_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_7399, new_AGEMA_signal_7398, add_sub1_1_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, addc_in[89]}), .c ({new_AGEMA_signal_7563, new_AGEMA_signal_7562, add_sub1_1_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_7241, new_AGEMA_signal_7240, add_sub1_1_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_6989, new_AGEMA_signal_6988, add_sub1_1_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_7399, new_AGEMA_signal_7398, add_sub1_1_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_6991, new_AGEMA_signal_6990, add_sub1_1_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_6283, new_AGEMA_signal_6282, addc_in[91]}), .c ({new_AGEMA_signal_7241, new_AGEMA_signal_7240, add_sub1_1_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, addc_in[88]}), .b ({new_AGEMA_signal_6611, new_AGEMA_signal_6610, add_sub1_1_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_6989, new_AGEMA_signal_6988, add_sub1_1_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, add_sub1_1_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_6617, new_AGEMA_signal_6616, add_sub1_1_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_6991, new_AGEMA_signal_6990, add_sub1_1_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_7565, new_AGEMA_signal_7564, add_sub1_1_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6997, new_AGEMA_signal_6996, add_sub1_1_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_8065, new_AGEMA_signal_8064, subc_out[87]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_7247, new_AGEMA_signal_7246, add_sub1_1_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, add_sub1_1_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, subc_out[86]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_8067, new_AGEMA_signal_8066, add_sub1_1_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_6629, new_AGEMA_signal_6628, add_sub1_1_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_8653, new_AGEMA_signal_8652, subc_out[85]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_7565, new_AGEMA_signal_7564, add_sub1_1_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, add_sub1_1_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_8067, new_AGEMA_signal_8066, add_sub1_1_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_7403, new_AGEMA_signal_7402, add_sub1_1_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_6247, new_AGEMA_signal_6246, addc_in[85]}), .c ({new_AGEMA_signal_7565, new_AGEMA_signal_7564, add_sub1_1_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_7247, new_AGEMA_signal_7246, add_sub1_1_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_6999, new_AGEMA_signal_6998, add_sub1_1_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_7403, new_AGEMA_signal_7402, add_sub1_1_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_7001, new_AGEMA_signal_7000, add_sub1_1_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_6259, new_AGEMA_signal_6258, addc_in[87]}), .c ({new_AGEMA_signal_7247, new_AGEMA_signal_7246, add_sub1_1_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, addc_in[84]}), .b ({new_AGEMA_signal_6625, new_AGEMA_signal_6624, add_sub1_1_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_6999, new_AGEMA_signal_6998, add_sub1_1_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6623, new_AGEMA_signal_6622, add_sub1_1_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, add_sub1_1_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_7001, new_AGEMA_signal_7000, add_sub1_1_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_7567, new_AGEMA_signal_7566, add_sub1_1_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_7007, new_AGEMA_signal_7006, add_sub1_1_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_8069, new_AGEMA_signal_8068, subc_out[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_7253, new_AGEMA_signal_7252, add_sub1_1_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7251, new_AGEMA_signal_7250, add_sub1_1_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_7405, new_AGEMA_signal_7404, subc_out[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_8071, new_AGEMA_signal_8070, add_sub1_1_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_6643, new_AGEMA_signal_6642, add_sub1_1_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, subc_out[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_7567, new_AGEMA_signal_7566, add_sub1_1_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6641, new_AGEMA_signal_6640, add_sub1_1_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_8071, new_AGEMA_signal_8070, add_sub1_1_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_7407, new_AGEMA_signal_7406, add_sub1_1_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_6223, new_AGEMA_signal_6222, addc_in[81]}), .c ({new_AGEMA_signal_7567, new_AGEMA_signal_7566, add_sub1_1_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_7253, new_AGEMA_signal_7252, add_sub1_1_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7009, new_AGEMA_signal_7008, add_sub1_1_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_7407, new_AGEMA_signal_7406, add_sub1_1_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_7011, new_AGEMA_signal_7010, add_sub1_1_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, addc_in[83]}), .c ({new_AGEMA_signal_7253, new_AGEMA_signal_7252, add_sub1_1_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, addc_in[80]}), .b ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, add_sub1_1_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_7009, new_AGEMA_signal_7008, add_sub1_1_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6637, new_AGEMA_signal_6636, add_sub1_1_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_6645, new_AGEMA_signal_6644, add_sub1_1_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_7011, new_AGEMA_signal_7010, add_sub1_1_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_7569, new_AGEMA_signal_7568, add_sub1_1_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_7017, new_AGEMA_signal_7016, add_sub1_1_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_8073, new_AGEMA_signal_8072, subc_out[79]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_7259, new_AGEMA_signal_7258, add_sub1_1_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7257, new_AGEMA_signal_7256, add_sub1_1_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_7409, new_AGEMA_signal_7408, subc_out[78]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_8075, new_AGEMA_signal_8074, add_sub1_1_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, add_sub1_1_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_8657, new_AGEMA_signal_8656, subc_out[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_7569, new_AGEMA_signal_7568, add_sub1_1_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6655, new_AGEMA_signal_6654, add_sub1_1_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_8075, new_AGEMA_signal_8074, add_sub1_1_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_7411, new_AGEMA_signal_7410, add_sub1_1_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, addc_in[77]}), .c ({new_AGEMA_signal_7569, new_AGEMA_signal_7568, add_sub1_1_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_7259, new_AGEMA_signal_7258, add_sub1_1_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7019, new_AGEMA_signal_7018, add_sub1_1_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_7411, new_AGEMA_signal_7410, add_sub1_1_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_7021, new_AGEMA_signal_7020, add_sub1_1_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_6211, new_AGEMA_signal_6210, addc_in[79]}), .c ({new_AGEMA_signal_7259, new_AGEMA_signal_7258, add_sub1_1_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, addc_in[76]}), .b ({new_AGEMA_signal_6653, new_AGEMA_signal_6652, add_sub1_1_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_7019, new_AGEMA_signal_7018, add_sub1_1_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, add_sub1_1_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_6659, new_AGEMA_signal_6658, add_sub1_1_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_7021, new_AGEMA_signal_7020, add_sub1_1_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_7571, new_AGEMA_signal_7570, add_sub1_1_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_7027, new_AGEMA_signal_7026, add_sub1_1_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_8077, new_AGEMA_signal_8076, subc_out[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_7265, new_AGEMA_signal_7264, add_sub1_1_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, add_sub1_1_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_7413, new_AGEMA_signal_7412, subc_out[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_8079, new_AGEMA_signal_8078, add_sub1_1_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_6671, new_AGEMA_signal_6670, add_sub1_1_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_8659, new_AGEMA_signal_8658, subc_out[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_7571, new_AGEMA_signal_7570, add_sub1_1_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6669, new_AGEMA_signal_6668, add_sub1_1_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_8079, new_AGEMA_signal_8078, add_sub1_1_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_7415, new_AGEMA_signal_7414, add_sub1_1_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, addc_in[73]}), .c ({new_AGEMA_signal_7571, new_AGEMA_signal_7570, add_sub1_1_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_7265, new_AGEMA_signal_7264, add_sub1_1_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, add_sub1_1_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_7415, new_AGEMA_signal_7414, add_sub1_1_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_7031, new_AGEMA_signal_7030, add_sub1_1_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, addc_in[75]}), .c ({new_AGEMA_signal_7265, new_AGEMA_signal_7264, add_sub1_1_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6169, new_AGEMA_signal_6168, addc_in[72]}), .b ({new_AGEMA_signal_6667, new_AGEMA_signal_6666, add_sub1_1_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, add_sub1_1_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6665, new_AGEMA_signal_6664, add_sub1_1_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_6673, new_AGEMA_signal_6672, add_sub1_1_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_7031, new_AGEMA_signal_7030, add_sub1_1_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_7573, new_AGEMA_signal_7572, add_sub1_1_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7037, new_AGEMA_signal_7036, add_sub1_1_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_8081, new_AGEMA_signal_8080, subc_out[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_7271, new_AGEMA_signal_7270, add_sub1_1_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7269, new_AGEMA_signal_7268, add_sub1_1_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_7417, new_AGEMA_signal_7416, subc_out[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_8083, new_AGEMA_signal_8082, add_sub1_1_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_6685, new_AGEMA_signal_6684, add_sub1_1_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_8661, new_AGEMA_signal_8660, subc_out[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_7573, new_AGEMA_signal_7572, add_sub1_1_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6683, new_AGEMA_signal_6682, add_sub1_1_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_8083, new_AGEMA_signal_8082, add_sub1_1_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, add_sub1_1_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, addc_in[69]}), .c ({new_AGEMA_signal_7573, new_AGEMA_signal_7572, add_sub1_1_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_7271, new_AGEMA_signal_7270, add_sub1_1_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7039, new_AGEMA_signal_7038, add_sub1_1_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, add_sub1_1_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_7041, new_AGEMA_signal_7040, add_sub1_1_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, addc_in[71]}), .c ({new_AGEMA_signal_7271, new_AGEMA_signal_7270, add_sub1_1_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, addc_in[68]}), .b ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, add_sub1_1_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_7039, new_AGEMA_signal_7038, add_sub1_1_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6679, new_AGEMA_signal_6678, add_sub1_1_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, add_sub1_1_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_7041, new_AGEMA_signal_7040, add_sub1_1_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_7575, new_AGEMA_signal_7574, add_sub1_1_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7047, new_AGEMA_signal_7046, add_sub1_1_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_8085, new_AGEMA_signal_8084, subc_out[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_7277, new_AGEMA_signal_7276, add_sub1_1_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7275, new_AGEMA_signal_7274, add_sub1_1_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_7421, new_AGEMA_signal_7420, subc_out[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_8087, new_AGEMA_signal_8086, add_sub1_1_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, add_sub1_1_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_8663, new_AGEMA_signal_8662, subc_out[65]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_7575, new_AGEMA_signal_7574, add_sub1_1_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6697, new_AGEMA_signal_6696, add_sub1_1_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_8087, new_AGEMA_signal_8086, add_sub1_1_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_7423, new_AGEMA_signal_7422, add_sub1_1_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, addc_in[65]}), .c ({new_AGEMA_signal_7575, new_AGEMA_signal_7574, add_sub1_1_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_7277, new_AGEMA_signal_7276, add_sub1_1_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7049, new_AGEMA_signal_7048, add_sub1_1_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_7423, new_AGEMA_signal_7422, add_sub1_1_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_7051, new_AGEMA_signal_7050, add_sub1_1_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, addc_in[67]}), .c ({new_AGEMA_signal_7277, new_AGEMA_signal_7276, add_sub1_1_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6121, new_AGEMA_signal_6120, addc_in[64]}), .b ({new_AGEMA_signal_6695, new_AGEMA_signal_6694, add_sub1_1_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_7049, new_AGEMA_signal_7048, add_sub1_1_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6693, new_AGEMA_signal_6692, add_sub1_1_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_6701, new_AGEMA_signal_6700, add_sub1_1_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_7051, new_AGEMA_signal_7050, add_sub1_1_subc_rom_sbox_0_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, add_sub1_2_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_8669, new_AGEMA_signal_8668, add_sub1_2_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_11421, new_AGEMA_signal_11420, subc_out[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, add_sub1_2_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_8833, new_AGEMA_signal_8832, add_sub1_2_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, subc_out[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_11423, new_AGEMA_signal_11422, add_sub1_2_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_8097, new_AGEMA_signal_8096, add_sub1_2_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_12369, new_AGEMA_signal_12368, subc_out[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, add_sub1_2_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_8095, new_AGEMA_signal_8094, add_sub1_2_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_11423, new_AGEMA_signal_11422, add_sub1_2_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_9491, new_AGEMA_signal_9490, add_sub1_2_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_7581, new_AGEMA_signal_7580, add_sub1_2_addc_out[1]}), .c ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, add_sub1_2_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, add_sub1_2_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_8671, new_AGEMA_signal_8670, add_sub1_2_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_9491, new_AGEMA_signal_9490, add_sub1_2_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_8673, new_AGEMA_signal_8672, add_sub1_2_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_7577, new_AGEMA_signal_7576, add_sub1_2_addc_out[3]}), .c ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, add_sub1_2_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_7583, new_AGEMA_signal_7582, add_sub1_2_addc_out[0]}), .b ({new_AGEMA_signal_8093, new_AGEMA_signal_8092, add_sub1_2_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_8671, new_AGEMA_signal_8670, add_sub1_2_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_8091, new_AGEMA_signal_8090, add_sub1_2_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_8099, new_AGEMA_signal_8098, add_sub1_2_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({new_AGEMA_signal_8673, new_AGEMA_signal_8672, add_sub1_2_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_7585, new_AGEMA_signal_7584, add_sub1_2_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, add_sub1_2_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_8103, new_AGEMA_signal_8102, subc_out[59]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_7283, new_AGEMA_signal_7282, add_sub1_2_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7281, new_AGEMA_signal_7280, add_sub1_2_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_7427, new_AGEMA_signal_7426, subc_out[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_8105, new_AGEMA_signal_8104, add_sub1_2_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_6717, new_AGEMA_signal_6716, add_sub1_2_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_8675, new_AGEMA_signal_8674, subc_out[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_7585, new_AGEMA_signal_7584, add_sub1_2_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6715, new_AGEMA_signal_6714, add_sub1_2_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_8105, new_AGEMA_signal_8104, add_sub1_2_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_7429, new_AGEMA_signal_7428, add_sub1_2_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, addc_in[57]}), .c ({new_AGEMA_signal_7585, new_AGEMA_signal_7584, add_sub1_2_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_7283, new_AGEMA_signal_7282, add_sub1_2_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7061, new_AGEMA_signal_7060, add_sub1_2_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_7429, new_AGEMA_signal_7428, add_sub1_2_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_7063, new_AGEMA_signal_7062, add_sub1_2_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, addc_in[59]}), .c ({new_AGEMA_signal_7283, new_AGEMA_signal_7282, add_sub1_2_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, addc_in[56]}), .b ({new_AGEMA_signal_6713, new_AGEMA_signal_6712, add_sub1_2_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_7061, new_AGEMA_signal_7060, add_sub1_2_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, add_sub1_2_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_6719, new_AGEMA_signal_6718, add_sub1_2_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({new_AGEMA_signal_7063, new_AGEMA_signal_7062, add_sub1_2_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_7587, new_AGEMA_signal_7586, add_sub1_2_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_7069, new_AGEMA_signal_7068, add_sub1_2_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_8107, new_AGEMA_signal_8106, subc_out[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_7289, new_AGEMA_signal_7288, add_sub1_2_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7287, new_AGEMA_signal_7286, add_sub1_2_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_7431, new_AGEMA_signal_7430, subc_out[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_8109, new_AGEMA_signal_8108, add_sub1_2_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_6731, new_AGEMA_signal_6730, add_sub1_2_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_8677, new_AGEMA_signal_8676, subc_out[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_7587, new_AGEMA_signal_7586, add_sub1_2_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, add_sub1_2_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_8109, new_AGEMA_signal_8108, add_sub1_2_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_7433, new_AGEMA_signal_7432, add_sub1_2_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, addc_in[53]}), .c ({new_AGEMA_signal_7587, new_AGEMA_signal_7586, add_sub1_2_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_7289, new_AGEMA_signal_7288, add_sub1_2_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7071, new_AGEMA_signal_7070, add_sub1_2_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_7433, new_AGEMA_signal_7432, add_sub1_2_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_7073, new_AGEMA_signal_7072, add_sub1_2_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, addc_in[55]}), .c ({new_AGEMA_signal_7289, new_AGEMA_signal_7288, add_sub1_2_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6049, new_AGEMA_signal_6048, addc_in[52]}), .b ({new_AGEMA_signal_6727, new_AGEMA_signal_6726, add_sub1_2_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_7071, new_AGEMA_signal_7070, add_sub1_2_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6725, new_AGEMA_signal_6724, add_sub1_2_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_6733, new_AGEMA_signal_6732, add_sub1_2_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({new_AGEMA_signal_7073, new_AGEMA_signal_7072, add_sub1_2_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_7589, new_AGEMA_signal_7588, add_sub1_2_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_7079, new_AGEMA_signal_7078, add_sub1_2_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_8111, new_AGEMA_signal_8110, subc_out[51]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_7295, new_AGEMA_signal_7294, add_sub1_2_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, add_sub1_2_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_7435, new_AGEMA_signal_7434, subc_out[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_8113, new_AGEMA_signal_8112, add_sub1_2_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_6745, new_AGEMA_signal_6744, add_sub1_2_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, subc_out[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_7589, new_AGEMA_signal_7588, add_sub1_2_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6743, new_AGEMA_signal_6742, add_sub1_2_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_8113, new_AGEMA_signal_8112, add_sub1_2_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_7437, new_AGEMA_signal_7436, add_sub1_2_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, addc_in[49]}), .c ({new_AGEMA_signal_7589, new_AGEMA_signal_7588, add_sub1_2_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_7295, new_AGEMA_signal_7294, add_sub1_2_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7081, new_AGEMA_signal_7080, add_sub1_2_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_7437, new_AGEMA_signal_7436, add_sub1_2_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_7083, new_AGEMA_signal_7082, add_sub1_2_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, addc_in[51]}), .c ({new_AGEMA_signal_7295, new_AGEMA_signal_7294, add_sub1_2_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6025, new_AGEMA_signal_6024, addc_in[48]}), .b ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, add_sub1_2_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_7081, new_AGEMA_signal_7080, add_sub1_2_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6739, new_AGEMA_signal_6738, add_sub1_2_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, add_sub1_2_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({new_AGEMA_signal_7083, new_AGEMA_signal_7082, add_sub1_2_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_7591, new_AGEMA_signal_7590, add_sub1_2_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, add_sub1_2_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_8115, new_AGEMA_signal_8114, subc_out[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_7301, new_AGEMA_signal_7300, add_sub1_2_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, add_sub1_2_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_7439, new_AGEMA_signal_7438, subc_out[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_8117, new_AGEMA_signal_8116, add_sub1_2_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, add_sub1_2_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_8681, new_AGEMA_signal_8680, subc_out[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_7591, new_AGEMA_signal_7590, add_sub1_2_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6757, new_AGEMA_signal_6756, add_sub1_2_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_8117, new_AGEMA_signal_8116, add_sub1_2_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_7441, new_AGEMA_signal_7440, add_sub1_2_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, addc_in[45]}), .c ({new_AGEMA_signal_7591, new_AGEMA_signal_7590, add_sub1_2_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_7301, new_AGEMA_signal_7300, add_sub1_2_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7091, new_AGEMA_signal_7090, add_sub1_2_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_7441, new_AGEMA_signal_7440, add_sub1_2_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_7093, new_AGEMA_signal_7092, add_sub1_2_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, addc_in[47]}), .c ({new_AGEMA_signal_7301, new_AGEMA_signal_7300, add_sub1_2_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6001, new_AGEMA_signal_6000, addc_in[44]}), .b ({new_AGEMA_signal_6755, new_AGEMA_signal_6754, add_sub1_2_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_7091, new_AGEMA_signal_7090, add_sub1_2_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, add_sub1_2_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_6761, new_AGEMA_signal_6760, add_sub1_2_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({new_AGEMA_signal_7093, new_AGEMA_signal_7092, add_sub1_2_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_7593, new_AGEMA_signal_7592, add_sub1_2_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_7099, new_AGEMA_signal_7098, add_sub1_2_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_8119, new_AGEMA_signal_8118, subc_out[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_7307, new_AGEMA_signal_7306, add_sub1_2_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7305, new_AGEMA_signal_7304, add_sub1_2_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_7443, new_AGEMA_signal_7442, subc_out[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_8121, new_AGEMA_signal_8120, add_sub1_2_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_6773, new_AGEMA_signal_6772, add_sub1_2_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_8683, new_AGEMA_signal_8682, subc_out[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_7593, new_AGEMA_signal_7592, add_sub1_2_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, add_sub1_2_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_8121, new_AGEMA_signal_8120, add_sub1_2_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_7445, new_AGEMA_signal_7444, add_sub1_2_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, addc_in[41]}), .c ({new_AGEMA_signal_7593, new_AGEMA_signal_7592, add_sub1_2_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_7307, new_AGEMA_signal_7306, add_sub1_2_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7101, new_AGEMA_signal_7100, add_sub1_2_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_7445, new_AGEMA_signal_7444, add_sub1_2_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_7103, new_AGEMA_signal_7102, add_sub1_2_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, addc_in[43]}), .c ({new_AGEMA_signal_7307, new_AGEMA_signal_7306, add_sub1_2_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5977, new_AGEMA_signal_5976, addc_in[40]}), .b ({new_AGEMA_signal_6769, new_AGEMA_signal_6768, add_sub1_2_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_7101, new_AGEMA_signal_7100, add_sub1_2_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6767, new_AGEMA_signal_6766, add_sub1_2_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_6775, new_AGEMA_signal_6774, add_sub1_2_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({new_AGEMA_signal_7103, new_AGEMA_signal_7102, add_sub1_2_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_7595, new_AGEMA_signal_7594, add_sub1_2_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7109, new_AGEMA_signal_7108, add_sub1_2_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_8123, new_AGEMA_signal_8122, subc_out[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_7313, new_AGEMA_signal_7312, add_sub1_2_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7311, new_AGEMA_signal_7310, add_sub1_2_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_7447, new_AGEMA_signal_7446, subc_out[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_8125, new_AGEMA_signal_8124, add_sub1_2_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_6787, new_AGEMA_signal_6786, add_sub1_2_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_8685, new_AGEMA_signal_8684, subc_out[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_7595, new_AGEMA_signal_7594, add_sub1_2_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6785, new_AGEMA_signal_6784, add_sub1_2_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_8125, new_AGEMA_signal_8124, add_sub1_2_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, add_sub1_2_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, addc_in[37]}), .c ({new_AGEMA_signal_7595, new_AGEMA_signal_7594, add_sub1_2_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_7313, new_AGEMA_signal_7312, add_sub1_2_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7111, new_AGEMA_signal_7110, add_sub1_2_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, add_sub1_2_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_7113, new_AGEMA_signal_7112, add_sub1_2_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, addc_in[39]}), .c ({new_AGEMA_signal_7313, new_AGEMA_signal_7312, add_sub1_2_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, addc_in[36]}), .b ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, add_sub1_2_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_7111, new_AGEMA_signal_7110, add_sub1_2_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6781, new_AGEMA_signal_6780, add_sub1_2_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_6789, new_AGEMA_signal_6788, add_sub1_2_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({new_AGEMA_signal_7113, new_AGEMA_signal_7112, add_sub1_2_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_7597, new_AGEMA_signal_7596, add_sub1_2_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7119, new_AGEMA_signal_7118, add_sub1_2_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_8127, new_AGEMA_signal_8126, subc_out[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_7319, new_AGEMA_signal_7318, add_sub1_2_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7317, new_AGEMA_signal_7316, add_sub1_2_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_7451, new_AGEMA_signal_7450, subc_out[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_8129, new_AGEMA_signal_8128, add_sub1_2_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_6801, new_AGEMA_signal_6800, add_sub1_2_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_8687, new_AGEMA_signal_8686, subc_out[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_7597, new_AGEMA_signal_7596, add_sub1_2_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6799, new_AGEMA_signal_6798, add_sub1_2_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_8129, new_AGEMA_signal_8128, add_sub1_2_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_7453, new_AGEMA_signal_7452, add_sub1_2_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, addc_in[33]}), .c ({new_AGEMA_signal_7597, new_AGEMA_signal_7596, add_sub1_2_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_7319, new_AGEMA_signal_7318, add_sub1_2_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7121, new_AGEMA_signal_7120, add_sub1_2_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_7453, new_AGEMA_signal_7452, add_sub1_2_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_7123, new_AGEMA_signal_7122, add_sub1_2_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, addc_in[35]}), .c ({new_AGEMA_signal_7319, new_AGEMA_signal_7318, add_sub1_2_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, addc_in[32]}), .b ({new_AGEMA_signal_6797, new_AGEMA_signal_6796, add_sub1_2_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_7121, new_AGEMA_signal_7120, add_sub1_2_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, add_sub1_2_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_6803, new_AGEMA_signal_6802, add_sub1_2_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({new_AGEMA_signal_7123, new_AGEMA_signal_7122, add_sub1_2_subc_rom_sbox_0_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_10455, new_AGEMA_signal_10454, add_sub1_3_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_8693, new_AGEMA_signal_8692, add_sub1_3_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_11425, new_AGEMA_signal_11424, subc_out[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_8841, new_AGEMA_signal_8840, add_sub1_3_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_8839, new_AGEMA_signal_8838, add_sub1_3_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_9493, new_AGEMA_signal_9492, subc_out[30]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_11427, new_AGEMA_signal_11426, add_sub1_3_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_8139, new_AGEMA_signal_8138, add_sub1_3_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_12371, new_AGEMA_signal_12370, subc_out[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_10455, new_AGEMA_signal_10454, add_sub1_3_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_8137, new_AGEMA_signal_8136, add_sub1_3_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_11427, new_AGEMA_signal_11426, add_sub1_3_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, add_sub1_3_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_7603, new_AGEMA_signal_7602, add_sub1_3_addc_out[1]}), .c ({new_AGEMA_signal_10455, new_AGEMA_signal_10454, add_sub1_3_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_8841, new_AGEMA_signal_8840, add_sub1_3_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_8695, new_AGEMA_signal_8694, add_sub1_3_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, add_sub1_3_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_8697, new_AGEMA_signal_8696, add_sub1_3_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_7599, new_AGEMA_signal_7598, add_sub1_3_addc_out[3]}), .c ({new_AGEMA_signal_8841, new_AGEMA_signal_8840, add_sub1_3_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_7605, new_AGEMA_signal_7604, add_sub1_3_addc_out[0]}), .b ({new_AGEMA_signal_8135, new_AGEMA_signal_8134, add_sub1_3_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_8695, new_AGEMA_signal_8694, add_sub1_3_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_8133, new_AGEMA_signal_8132, add_sub1_3_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_8141, new_AGEMA_signal_8140, add_sub1_3_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({new_AGEMA_signal_8697, new_AGEMA_signal_8696, add_sub1_3_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_7607, new_AGEMA_signal_7606, add_sub1_3_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_7131, new_AGEMA_signal_7130, add_sub1_3_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_8145, new_AGEMA_signal_8144, subc_out[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_7325, new_AGEMA_signal_7324, add_sub1_3_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7323, new_AGEMA_signal_7322, add_sub1_3_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_7457, new_AGEMA_signal_7456, subc_out[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_8147, new_AGEMA_signal_8146, add_sub1_3_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_6819, new_AGEMA_signal_6818, add_sub1_3_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_8699, new_AGEMA_signal_8698, subc_out[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_7607, new_AGEMA_signal_7606, add_sub1_3_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6817, new_AGEMA_signal_6816, add_sub1_3_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_8147, new_AGEMA_signal_8146, add_sub1_3_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_7459, new_AGEMA_signal_7458, add_sub1_3_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, addc_in[25]}), .c ({new_AGEMA_signal_7607, new_AGEMA_signal_7606, add_sub1_3_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_7325, new_AGEMA_signal_7324, add_sub1_3_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7133, new_AGEMA_signal_7132, add_sub1_3_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_7459, new_AGEMA_signal_7458, add_sub1_3_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_7135, new_AGEMA_signal_7134, add_sub1_3_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, addc_in[27]}), .c ({new_AGEMA_signal_7325, new_AGEMA_signal_7324, add_sub1_3_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5881, new_AGEMA_signal_5880, addc_in[24]}), .b ({new_AGEMA_signal_6815, new_AGEMA_signal_6814, add_sub1_3_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_7133, new_AGEMA_signal_7132, add_sub1_3_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6813, new_AGEMA_signal_6812, add_sub1_3_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_6821, new_AGEMA_signal_6820, add_sub1_3_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({new_AGEMA_signal_7135, new_AGEMA_signal_7134, add_sub1_3_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_7609, new_AGEMA_signal_7608, add_sub1_3_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_7141, new_AGEMA_signal_7140, add_sub1_3_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_8149, new_AGEMA_signal_8148, subc_out[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_7331, new_AGEMA_signal_7330, add_sub1_3_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7329, new_AGEMA_signal_7328, add_sub1_3_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_7461, new_AGEMA_signal_7460, subc_out[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_8151, new_AGEMA_signal_8150, add_sub1_3_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_6833, new_AGEMA_signal_6832, add_sub1_3_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_8701, new_AGEMA_signal_8700, subc_out[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_7609, new_AGEMA_signal_7608, add_sub1_3_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, add_sub1_3_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_8151, new_AGEMA_signal_8150, add_sub1_3_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_7463, new_AGEMA_signal_7462, add_sub1_3_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, addc_in[21]}), .c ({new_AGEMA_signal_7609, new_AGEMA_signal_7608, add_sub1_3_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_7331, new_AGEMA_signal_7330, add_sub1_3_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, add_sub1_3_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_7463, new_AGEMA_signal_7462, add_sub1_3_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_7145, new_AGEMA_signal_7144, add_sub1_3_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, addc_in[23]}), .c ({new_AGEMA_signal_7331, new_AGEMA_signal_7330, add_sub1_3_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, addc_in[20]}), .b ({new_AGEMA_signal_6829, new_AGEMA_signal_6828, add_sub1_3_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, add_sub1_3_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6827, new_AGEMA_signal_6826, add_sub1_3_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_6835, new_AGEMA_signal_6834, add_sub1_3_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({new_AGEMA_signal_7145, new_AGEMA_signal_7144, add_sub1_3_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_7611, new_AGEMA_signal_7610, add_sub1_3_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_7151, new_AGEMA_signal_7150, add_sub1_3_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_8153, new_AGEMA_signal_8152, subc_out[19]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_7337, new_AGEMA_signal_7336, add_sub1_3_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7335, new_AGEMA_signal_7334, add_sub1_3_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_7465, new_AGEMA_signal_7464, subc_out[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_8155, new_AGEMA_signal_8154, add_sub1_3_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_6847, new_AGEMA_signal_6846, add_sub1_3_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, subc_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_7611, new_AGEMA_signal_7610, add_sub1_3_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6845, new_AGEMA_signal_6844, add_sub1_3_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_8155, new_AGEMA_signal_8154, add_sub1_3_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_7467, new_AGEMA_signal_7466, add_sub1_3_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, addc_in[17]}), .c ({new_AGEMA_signal_7611, new_AGEMA_signal_7610, add_sub1_3_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_7337, new_AGEMA_signal_7336, add_sub1_3_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7153, new_AGEMA_signal_7152, add_sub1_3_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_7467, new_AGEMA_signal_7466, add_sub1_3_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_7155, new_AGEMA_signal_7154, add_sub1_3_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, addc_in[19]}), .c ({new_AGEMA_signal_7337, new_AGEMA_signal_7336, add_sub1_3_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5833, new_AGEMA_signal_5832, addc_in[16]}), .b ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, add_sub1_3_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_7153, new_AGEMA_signal_7152, add_sub1_3_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6841, new_AGEMA_signal_6840, add_sub1_3_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, add_sub1_3_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({new_AGEMA_signal_7155, new_AGEMA_signal_7154, add_sub1_3_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_7613, new_AGEMA_signal_7612, add_sub1_3_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, add_sub1_3_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_8157, new_AGEMA_signal_8156, subc_out[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_7343, new_AGEMA_signal_7342, add_sub1_3_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, add_sub1_3_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_7469, new_AGEMA_signal_7468, subc_out[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_8159, new_AGEMA_signal_8158, add_sub1_3_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_6861, new_AGEMA_signal_6860, add_sub1_3_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_8705, new_AGEMA_signal_8704, subc_out[13]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_7613, new_AGEMA_signal_7612, add_sub1_3_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6859, new_AGEMA_signal_6858, add_sub1_3_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_8159, new_AGEMA_signal_8158, add_sub1_3_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_7471, new_AGEMA_signal_7470, add_sub1_3_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, addc_in[13]}), .c ({new_AGEMA_signal_7613, new_AGEMA_signal_7612, add_sub1_3_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_7343, new_AGEMA_signal_7342, add_sub1_3_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7163, new_AGEMA_signal_7162, add_sub1_3_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_7471, new_AGEMA_signal_7470, add_sub1_3_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_7165, new_AGEMA_signal_7164, add_sub1_3_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, addc_in[15]}), .c ({new_AGEMA_signal_7343, new_AGEMA_signal_7342, add_sub1_3_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5809, new_AGEMA_signal_5808, addc_in[12]}), .b ({new_AGEMA_signal_6857, new_AGEMA_signal_6856, add_sub1_3_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_7163, new_AGEMA_signal_7162, add_sub1_3_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6855, new_AGEMA_signal_6854, add_sub1_3_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_6863, new_AGEMA_signal_6862, add_sub1_3_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({new_AGEMA_signal_7165, new_AGEMA_signal_7164, add_sub1_3_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_7615, new_AGEMA_signal_7614, add_sub1_3_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_7171, new_AGEMA_signal_7170, add_sub1_3_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_8161, new_AGEMA_signal_8160, subc_out[11]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_7349, new_AGEMA_signal_7348, add_sub1_3_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7347, new_AGEMA_signal_7346, add_sub1_3_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, subc_out[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_8163, new_AGEMA_signal_8162, add_sub1_3_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_6875, new_AGEMA_signal_6874, add_sub1_3_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_8707, new_AGEMA_signal_8706, subc_out[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_7615, new_AGEMA_signal_7614, add_sub1_3_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, add_sub1_3_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_8163, new_AGEMA_signal_8162, add_sub1_3_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_7475, new_AGEMA_signal_7474, add_sub1_3_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, addc_in[9]}), .c ({new_AGEMA_signal_7615, new_AGEMA_signal_7614, add_sub1_3_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_7349, new_AGEMA_signal_7348, add_sub1_3_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7173, new_AGEMA_signal_7172, add_sub1_3_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_7475, new_AGEMA_signal_7474, add_sub1_3_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_7175, new_AGEMA_signal_7174, add_sub1_3_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, addc_in[11]}), .c ({new_AGEMA_signal_7349, new_AGEMA_signal_7348, add_sub1_3_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, addc_in[8]}), .b ({new_AGEMA_signal_6871, new_AGEMA_signal_6870, add_sub1_3_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_7173, new_AGEMA_signal_7172, add_sub1_3_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6869, new_AGEMA_signal_6868, add_sub1_3_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_6877, new_AGEMA_signal_6876, add_sub1_3_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({new_AGEMA_signal_7175, new_AGEMA_signal_7174, add_sub1_3_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_7617, new_AGEMA_signal_7616, add_sub1_3_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7181, new_AGEMA_signal_7180, add_sub1_3_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_8165, new_AGEMA_signal_8164, subc_out[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_7355, new_AGEMA_signal_7354, add_sub1_3_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7353, new_AGEMA_signal_7352, add_sub1_3_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_7477, new_AGEMA_signal_7476, subc_out[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_8167, new_AGEMA_signal_8166, add_sub1_3_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_6889, new_AGEMA_signal_6888, add_sub1_3_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_8709, new_AGEMA_signal_8708, subc_out[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_7617, new_AGEMA_signal_7616, add_sub1_3_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_6887, new_AGEMA_signal_6886, add_sub1_3_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_8167, new_AGEMA_signal_8166, add_sub1_3_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_7479, new_AGEMA_signal_7478, add_sub1_3_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, addc_in[5]}), .c ({new_AGEMA_signal_7617, new_AGEMA_signal_7616, add_sub1_3_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_7355, new_AGEMA_signal_7354, add_sub1_3_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7183, new_AGEMA_signal_7182, add_sub1_3_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_7479, new_AGEMA_signal_7478, add_sub1_3_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, add_sub1_3_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, addc_in[7]}), .c ({new_AGEMA_signal_7355, new_AGEMA_signal_7354, add_sub1_3_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, addc_in[4]}), .b ({new_AGEMA_signal_6885, new_AGEMA_signal_6884, add_sub1_3_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_7183, new_AGEMA_signal_7182, add_sub1_3_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6883, new_AGEMA_signal_6882, add_sub1_3_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_6891, new_AGEMA_signal_6890, add_sub1_3_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, add_sub1_3_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_7619, new_AGEMA_signal_7618, add_sub1_3_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7191, new_AGEMA_signal_7190, add_sub1_3_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_8169, new_AGEMA_signal_8168, subc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_7361, new_AGEMA_signal_7360, add_sub1_3_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7359, new_AGEMA_signal_7358, add_sub1_3_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_7481, new_AGEMA_signal_7480, subc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_8171, new_AGEMA_signal_8170, add_sub1_3_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, add_sub1_3_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_8711, new_AGEMA_signal_8710, subc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_7619, new_AGEMA_signal_7618, add_sub1_3_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_6901, new_AGEMA_signal_6900, add_sub1_3_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_8171, new_AGEMA_signal_8170, add_sub1_3_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_7483, new_AGEMA_signal_7482, add_sub1_3_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, addc_in[1]}), .c ({new_AGEMA_signal_7619, new_AGEMA_signal_7618, add_sub1_3_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_7361, new_AGEMA_signal_7360, add_sub1_3_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7193, new_AGEMA_signal_7192, add_sub1_3_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_7483, new_AGEMA_signal_7482, add_sub1_3_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_7195, new_AGEMA_signal_7194, add_sub1_3_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, addc_in[3]}), .c ({new_AGEMA_signal_7361, new_AGEMA_signal_7360, add_sub1_3_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, addc_in[0]}), .b ({new_AGEMA_signal_6899, new_AGEMA_signal_6898, add_sub1_3_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_7193, new_AGEMA_signal_7192, add_sub1_3_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6897, new_AGEMA_signal_6896, add_sub1_3_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_6905, new_AGEMA_signal_6904, add_sub1_3_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({new_AGEMA_signal_7195, new_AGEMA_signal_7194, add_sub1_3_subc_rom_sbox_0_ANF_2_t6}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8639, new_AGEMA_signal_8638, subc_out[97]}), .a ({new_AGEMA_signal_8631, new_AGEMA_signal_8630, subc_out[113]}), .c ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7391, new_AGEMA_signal_7390, subc_out[98]}), .a ({new_AGEMA_signal_7375, new_AGEMA_signal_7374, subc_out[114]}), .c ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8043, new_AGEMA_signal_8042, subc_out[99]}), .a ({new_AGEMA_signal_8027, new_AGEMA_signal_8026, subc_out[115]}), .c ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, subc_out[101]}), .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, subc_out[117]}), .c ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7387, new_AGEMA_signal_7386, subc_out[102]}), .a ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, subc_out[118]}), .c ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8039, new_AGEMA_signal_8038, subc_out[103]}), .a ({new_AGEMA_signal_8023, new_AGEMA_signal_8022, subc_out[119]}), .c ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, subc_out[105]}), .a ({new_AGEMA_signal_8627, new_AGEMA_signal_8626, subc_out[121]}), .c ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7383, new_AGEMA_signal_7382, subc_out[106]}), .a ({new_AGEMA_signal_7367, new_AGEMA_signal_7366, subc_out[122]}), .c ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8035, new_AGEMA_signal_8034, subc_out[107]}), .a ({new_AGEMA_signal_8019, new_AGEMA_signal_8018, subc_out[123]}), .c ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8633, new_AGEMA_signal_8632, subc_out[109]}), .a ({new_AGEMA_signal_12365, new_AGEMA_signal_12364, subc_out[125]}), .c ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7379, new_AGEMA_signal_7378, subc_out[110]}), .a ({new_AGEMA_signal_9481, new_AGEMA_signal_9480, subc_out[126]}), .c ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8031, new_AGEMA_signal_8030, subc_out[111]}), .a ({new_AGEMA_signal_11413, new_AGEMA_signal_11412, subc_out[127]}), .c ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8631, new_AGEMA_signal_8630, subc_out[113]}), .a ({new_AGEMA_signal_8639, new_AGEMA_signal_8638, subc_out[97]}), .c ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7375, new_AGEMA_signal_7374, subc_out[114]}), .a ({new_AGEMA_signal_7391, new_AGEMA_signal_7390, subc_out[98]}), .c ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8027, new_AGEMA_signal_8026, subc_out[115]}), .a ({new_AGEMA_signal_8043, new_AGEMA_signal_8042, subc_out[99]}), .c ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, subc_out[117]}), .a ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, subc_out[101]}), .c ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, subc_out[118]}), .a ({new_AGEMA_signal_7387, new_AGEMA_signal_7386, subc_out[102]}), .c ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8023, new_AGEMA_signal_8022, subc_out[119]}), .a ({new_AGEMA_signal_8039, new_AGEMA_signal_8038, subc_out[103]}), .c ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8627, new_AGEMA_signal_8626, subc_out[121]}), .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, subc_out[105]}), .c ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7367, new_AGEMA_signal_7366, subc_out[122]}), .a ({new_AGEMA_signal_7383, new_AGEMA_signal_7382, subc_out[106]}), .c ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8019, new_AGEMA_signal_8018, subc_out[123]}), .a ({new_AGEMA_signal_8035, new_AGEMA_signal_8034, subc_out[107]}), .c ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_12365, new_AGEMA_signal_12364, subc_out[125]}), .a ({new_AGEMA_signal_8633, new_AGEMA_signal_8632, subc_out[109]}), .c ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9481, new_AGEMA_signal_9480, subc_out[126]}), .a ({new_AGEMA_signal_7379, new_AGEMA_signal_7378, subc_out[110]}), .c ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11413, new_AGEMA_signal_11412, subc_out[127]}), .a ({new_AGEMA_signal_8031, new_AGEMA_signal_8030, subc_out[111]}), .c ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_12367, new_AGEMA_signal_12366, subc_out[93]}), .a ({new_AGEMA_signal_8657, new_AGEMA_signal_8656, subc_out[77]}), .c ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9485, new_AGEMA_signal_9484, subc_out[94]}), .a ({new_AGEMA_signal_7409, new_AGEMA_signal_7408, subc_out[78]}), .c ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11417, new_AGEMA_signal_11416, subc_out[95]}), .a ({new_AGEMA_signal_8073, new_AGEMA_signal_8072, subc_out[79]}), .c ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8663, new_AGEMA_signal_8662, subc_out[65]}), .a ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, subc_out[81]}), .c ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7421, new_AGEMA_signal_7420, subc_out[66]}), .a ({new_AGEMA_signal_7405, new_AGEMA_signal_7404, subc_out[82]}), .c ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8085, new_AGEMA_signal_8084, subc_out[67]}), .a ({new_AGEMA_signal_8069, new_AGEMA_signal_8068, subc_out[83]}), .c ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8661, new_AGEMA_signal_8660, subc_out[69]}), .a ({new_AGEMA_signal_8653, new_AGEMA_signal_8652, subc_out[85]}), .c ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7417, new_AGEMA_signal_7416, subc_out[70]}), .a ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, subc_out[86]}), .c ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8081, new_AGEMA_signal_8080, subc_out[71]}), .a ({new_AGEMA_signal_8065, new_AGEMA_signal_8064, subc_out[87]}), .c ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8659, new_AGEMA_signal_8658, subc_out[73]}), .a ({new_AGEMA_signal_8651, new_AGEMA_signal_8650, subc_out[89]}), .c ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7413, new_AGEMA_signal_7412, subc_out[74]}), .a ({new_AGEMA_signal_7397, new_AGEMA_signal_7396, subc_out[90]}), .c ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8077, new_AGEMA_signal_8076, subc_out[75]}), .a ({new_AGEMA_signal_8061, new_AGEMA_signal_8060, subc_out[91]}), .c ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8657, new_AGEMA_signal_8656, subc_out[77]}), .a ({new_AGEMA_signal_12367, new_AGEMA_signal_12366, subc_out[93]}), .c ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7409, new_AGEMA_signal_7408, subc_out[78]}), .a ({new_AGEMA_signal_9485, new_AGEMA_signal_9484, subc_out[94]}), .c ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8073, new_AGEMA_signal_8072, subc_out[79]}), .a ({new_AGEMA_signal_11417, new_AGEMA_signal_11416, subc_out[95]}), .c ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, subc_out[81]}), .a ({new_AGEMA_signal_8663, new_AGEMA_signal_8662, subc_out[65]}), .c ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7405, new_AGEMA_signal_7404, subc_out[82]}), .a ({new_AGEMA_signal_7421, new_AGEMA_signal_7420, subc_out[66]}), .c ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8069, new_AGEMA_signal_8068, subc_out[83]}), .a ({new_AGEMA_signal_8085, new_AGEMA_signal_8084, subc_out[67]}), .c ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8653, new_AGEMA_signal_8652, subc_out[85]}), .a ({new_AGEMA_signal_8661, new_AGEMA_signal_8660, subc_out[69]}), .c ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, subc_out[86]}), .a ({new_AGEMA_signal_7417, new_AGEMA_signal_7416, subc_out[70]}), .c ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8065, new_AGEMA_signal_8064, subc_out[87]}), .a ({new_AGEMA_signal_8081, new_AGEMA_signal_8080, subc_out[71]}), .c ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8651, new_AGEMA_signal_8650, subc_out[89]}), .a ({new_AGEMA_signal_8659, new_AGEMA_signal_8658, subc_out[73]}), .c ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7397, new_AGEMA_signal_7396, subc_out[90]}), .a ({new_AGEMA_signal_7413, new_AGEMA_signal_7412, subc_out[74]}), .c ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8061, new_AGEMA_signal_8060, subc_out[91]}), .a ({new_AGEMA_signal_8077, new_AGEMA_signal_8076, subc_out[75]}), .c ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8675, new_AGEMA_signal_8674, subc_out[57]}), .a ({new_AGEMA_signal_8683, new_AGEMA_signal_8682, subc_out[41]}), .c ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7427, new_AGEMA_signal_7426, subc_out[58]}), .a ({new_AGEMA_signal_7443, new_AGEMA_signal_7442, subc_out[42]}), .c ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8103, new_AGEMA_signal_8102, subc_out[59]}), .a ({new_AGEMA_signal_8119, new_AGEMA_signal_8118, subc_out[43]}), .c ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_12369, new_AGEMA_signal_12368, subc_out[61]}), .a ({new_AGEMA_signal_8681, new_AGEMA_signal_8680, subc_out[45]}), .c ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, subc_out[62]}), .a ({new_AGEMA_signal_7439, new_AGEMA_signal_7438, subc_out[46]}), .c ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11421, new_AGEMA_signal_11420, subc_out[63]}), .a ({new_AGEMA_signal_8115, new_AGEMA_signal_8114, subc_out[47]}), .c ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8687, new_AGEMA_signal_8686, subc_out[33]}), .a ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, subc_out[49]}), .c ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7451, new_AGEMA_signal_7450, subc_out[34]}), .a ({new_AGEMA_signal_7435, new_AGEMA_signal_7434, subc_out[50]}), .c ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8127, new_AGEMA_signal_8126, subc_out[35]}), .a ({new_AGEMA_signal_8111, new_AGEMA_signal_8110, subc_out[51]}), .c ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8685, new_AGEMA_signal_8684, subc_out[37]}), .a ({new_AGEMA_signal_8677, new_AGEMA_signal_8676, subc_out[53]}), .c ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7447, new_AGEMA_signal_7446, subc_out[38]}), .a ({new_AGEMA_signal_7431, new_AGEMA_signal_7430, subc_out[54]}), .c ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8123, new_AGEMA_signal_8122, subc_out[39]}), .a ({new_AGEMA_signal_8107, new_AGEMA_signal_8106, subc_out[55]}), .c ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8683, new_AGEMA_signal_8682, subc_out[41]}), .a ({new_AGEMA_signal_8675, new_AGEMA_signal_8674, subc_out[57]}), .c ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7443, new_AGEMA_signal_7442, subc_out[42]}), .a ({new_AGEMA_signal_7427, new_AGEMA_signal_7426, subc_out[58]}), .c ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8119, new_AGEMA_signal_8118, subc_out[43]}), .a ({new_AGEMA_signal_8103, new_AGEMA_signal_8102, subc_out[59]}), .c ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8681, new_AGEMA_signal_8680, subc_out[45]}), .a ({new_AGEMA_signal_12369, new_AGEMA_signal_12368, subc_out[61]}), .c ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7439, new_AGEMA_signal_7438, subc_out[46]}), .a ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, subc_out[62]}), .c ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8115, new_AGEMA_signal_8114, subc_out[47]}), .a ({new_AGEMA_signal_11421, new_AGEMA_signal_11420, subc_out[63]}), .c ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, subc_out[49]}), .a ({new_AGEMA_signal_8687, new_AGEMA_signal_8686, subc_out[33]}), .c ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7435, new_AGEMA_signal_7434, subc_out[50]}), .a ({new_AGEMA_signal_7451, new_AGEMA_signal_7450, subc_out[34]}), .c ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8111, new_AGEMA_signal_8110, subc_out[51]}), .a ({new_AGEMA_signal_8127, new_AGEMA_signal_8126, subc_out[35]}), .c ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8677, new_AGEMA_signal_8676, subc_out[53]}), .a ({new_AGEMA_signal_8685, new_AGEMA_signal_8684, subc_out[37]}), .c ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7431, new_AGEMA_signal_7430, subc_out[54]}), .a ({new_AGEMA_signal_7447, new_AGEMA_signal_7446, subc_out[38]}), .c ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8107, new_AGEMA_signal_8106, subc_out[55]}), .a ({new_AGEMA_signal_8123, new_AGEMA_signal_8122, subc_out[39]}), .c ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8701, new_AGEMA_signal_8700, subc_out[21]}), .a ({new_AGEMA_signal_8709, new_AGEMA_signal_8708, subc_out[5]}), .c ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7461, new_AGEMA_signal_7460, subc_out[22]}), .a ({new_AGEMA_signal_7477, new_AGEMA_signal_7476, subc_out[6]}), .c ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8149, new_AGEMA_signal_8148, subc_out[23]}), .a ({new_AGEMA_signal_8165, new_AGEMA_signal_8164, subc_out[7]}), .c ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8699, new_AGEMA_signal_8698, subc_out[25]}), .a ({new_AGEMA_signal_8707, new_AGEMA_signal_8706, subc_out[9]}), .c ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7457, new_AGEMA_signal_7456, subc_out[26]}), .a ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, subc_out[10]}), .c ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8145, new_AGEMA_signal_8144, subc_out[27]}), .a ({new_AGEMA_signal_8161, new_AGEMA_signal_8160, subc_out[11]}), .c ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_12371, new_AGEMA_signal_12370, subc_out[29]}), .a ({new_AGEMA_signal_8705, new_AGEMA_signal_8704, subc_out[13]}), .c ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9493, new_AGEMA_signal_9492, subc_out[30]}), .a ({new_AGEMA_signal_7469, new_AGEMA_signal_7468, subc_out[14]}), .c ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11425, new_AGEMA_signal_11424, subc_out[31]}), .a ({new_AGEMA_signal_8157, new_AGEMA_signal_8156, subc_out[15]}), .c ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8711, new_AGEMA_signal_8710, subc_out[1]}), .a ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, subc_out[17]}), .c ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7481, new_AGEMA_signal_7480, subc_out[2]}), .a ({new_AGEMA_signal_7465, new_AGEMA_signal_7464, subc_out[18]}), .c ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8169, new_AGEMA_signal_8168, subc_out[3]}), .a ({new_AGEMA_signal_8153, new_AGEMA_signal_8152, subc_out[19]}), .c ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8709, new_AGEMA_signal_8708, subc_out[5]}), .a ({new_AGEMA_signal_8701, new_AGEMA_signal_8700, subc_out[21]}), .c ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7477, new_AGEMA_signal_7476, subc_out[6]}), .a ({new_AGEMA_signal_7461, new_AGEMA_signal_7460, subc_out[22]}), .c ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8165, new_AGEMA_signal_8164, subc_out[7]}), .a ({new_AGEMA_signal_8149, new_AGEMA_signal_8148, subc_out[23]}), .c ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8707, new_AGEMA_signal_8706, subc_out[9]}), .a ({new_AGEMA_signal_8699, new_AGEMA_signal_8698, subc_out[25]}), .c ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, subc_out[10]}), .a ({new_AGEMA_signal_7457, new_AGEMA_signal_7456, subc_out[26]}), .c ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8161, new_AGEMA_signal_8160, subc_out[11]}), .a ({new_AGEMA_signal_8145, new_AGEMA_signal_8144, subc_out[27]}), .c ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8705, new_AGEMA_signal_8704, subc_out[13]}), .a ({new_AGEMA_signal_12371, new_AGEMA_signal_12370, subc_out[29]}), .c ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7469, new_AGEMA_signal_7468, subc_out[14]}), .a ({new_AGEMA_signal_9493, new_AGEMA_signal_9492, subc_out[30]}), .c ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8157, new_AGEMA_signal_8156, subc_out[15]}), .a ({new_AGEMA_signal_11425, new_AGEMA_signal_11424, subc_out[31]}), .c ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, subc_out[17]}), .a ({new_AGEMA_signal_8711, new_AGEMA_signal_8710, subc_out[1]}), .c ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7465, new_AGEMA_signal_7464, subc_out[18]}), .a ({new_AGEMA_signal_7481, new_AGEMA_signal_7480, subc_out[2]}), .c ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8153, new_AGEMA_signal_8152, subc_out[19]}), .a ({new_AGEMA_signal_8169, new_AGEMA_signal_8168, subc_out[3]}), .c ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U44 ( .a ({new_AGEMA_signal_8919, new_AGEMA_signal_8918, mcs1_mcs_mat1_0_mcs_out[90]}), .b ({new_AGEMA_signal_13527, new_AGEMA_signal_13526, mcs1_mcs_mat1_0_mcs_out[94]}), .c ({new_AGEMA_signal_13995, new_AGEMA_signal_13994, mcs1_mcs_mat1_0_n93}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .c ({new_AGEMA_signal_13029, new_AGEMA_signal_13028, mcs1_mcs_mat1_0_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .b ({new_AGEMA_signal_7669, new_AGEMA_signal_7668, mcs1_mcs_mat1_0_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8173, new_AGEMA_signal_8172, mcs1_mcs_mat1_0_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_7669, new_AGEMA_signal_7668, mcs1_mcs_mat1_0_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_8897, new_AGEMA_signal_8896, mcs1_mcs_mat1_0_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_9517, new_AGEMA_signal_9516, mcs1_mcs_mat1_0_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_7671, new_AGEMA_signal_7670, mcs1_mcs_mat1_0_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_8897, new_AGEMA_signal_8896, mcs1_mcs_mat1_0_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({new_AGEMA_signal_7671, new_AGEMA_signal_7670, mcs1_mcs_mat1_0_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_7673, new_AGEMA_signal_7672, mcs1_mcs_mat1_0_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, mcs1_mcs_mat1_0_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_10481, new_AGEMA_signal_10480, mcs1_mcs_mat1_0_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_8179, new_AGEMA_signal_8178, mcs1_mcs_mat1_0_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_8903, new_AGEMA_signal_8902, mcs1_mcs_mat1_0_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .c ({new_AGEMA_signal_8179, new_AGEMA_signal_8178, mcs1_mcs_mat1_0_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .b ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, mcs1_mcs_mat1_0_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_7673, new_AGEMA_signal_7672, mcs1_mcs_mat1_0_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_13521, new_AGEMA_signal_13520, mcs1_mcs_mat1_0_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_14005, new_AGEMA_signal_14004, mcs1_mcs_mat1_0_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_10487, new_AGEMA_signal_10486, mcs1_mcs_mat1_0_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_13521, new_AGEMA_signal_13520, mcs1_mcs_mat1_0_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({new_AGEMA_signal_10487, new_AGEMA_signal_10486, mcs1_mcs_mat1_0_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_7675, new_AGEMA_signal_7674, mcs1_mcs_mat1_0_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({new_AGEMA_signal_8911, new_AGEMA_signal_8910, mcs1_mcs_mat1_0_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_9533, new_AGEMA_signal_9532, mcs1_mcs_mat1_0_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_7677, new_AGEMA_signal_7676, mcs1_mcs_mat1_0_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_8911, new_AGEMA_signal_8910, mcs1_mcs_mat1_0_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .b ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .c ({new_AGEMA_signal_9535, new_AGEMA_signal_9534, mcs1_mcs_mat1_0_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({new_AGEMA_signal_7677, new_AGEMA_signal_7676, mcs1_mcs_mat1_0_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_7679, new_AGEMA_signal_7678, mcs1_mcs_mat1_0_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_8915, new_AGEMA_signal_8914, mcs1_mcs_mat1_0_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_7679, new_AGEMA_signal_7678, mcs1_mcs_mat1_0_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .c ({new_AGEMA_signal_8187, new_AGEMA_signal_8186, mcs1_mcs_mat1_0_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_7679, new_AGEMA_signal_7678, mcs1_mcs_mat1_0_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_13035, new_AGEMA_signal_13034, mcs1_mcs_mat1_0_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .c ({new_AGEMA_signal_13527, new_AGEMA_signal_13526, mcs1_mcs_mat1_0_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_10501, new_AGEMA_signal_10500, mcs1_mcs_mat1_0_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_13035, new_AGEMA_signal_13034, mcs1_mcs_mat1_0_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_13037, new_AGEMA_signal_13036, mcs1_mcs_mat1_0_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({new_AGEMA_signal_10501, new_AGEMA_signal_10500, mcs1_mcs_mat1_0_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .b ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .c ({new_AGEMA_signal_8919, new_AGEMA_signal_8918, mcs1_mcs_mat1_0_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .b ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_8921, new_AGEMA_signal_8920, mcs1_mcs_mat1_0_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, mcs1_mcs_mat1_0_mcs_out[87]}), .c ({new_AGEMA_signal_10503, new_AGEMA_signal_10502, mcs1_mcs_mat1_0_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .c ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, mcs1_mcs_mat1_0_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .c ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, mcs1_mcs_mat1_0_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_7681, new_AGEMA_signal_7680, mcs1_mcs_mat1_0_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_10513, new_AGEMA_signal_10512, mcs1_mcs_mat1_0_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_11481, new_AGEMA_signal_11480, mcs1_mcs_mat1_0_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({new_AGEMA_signal_10513, new_AGEMA_signal_10512, mcs1_mcs_mat1_0_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_7683, new_AGEMA_signal_7682, mcs1_mcs_mat1_0_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_8193, new_AGEMA_signal_8192, mcs1_mcs_mat1_0_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_7683, new_AGEMA_signal_7682, mcs1_mcs_mat1_0_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({new_AGEMA_signal_7685, new_AGEMA_signal_7684, mcs1_mcs_mat1_0_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_7687, new_AGEMA_signal_7686, mcs1_mcs_mat1_0_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .c ({new_AGEMA_signal_9565, new_AGEMA_signal_9564, mcs1_mcs_mat1_0_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_7687, new_AGEMA_signal_7686, mcs1_mcs_mat1_0_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_14437, new_AGEMA_signal_14436, mcs1_mcs_mat1_0_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_10525, new_AGEMA_signal_10524, mcs1_mcs_mat1_0_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_14925, new_AGEMA_signal_14924, mcs1_mcs_mat1_0_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_14017, new_AGEMA_signal_14016, mcs1_mcs_mat1_0_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_14437, new_AGEMA_signal_14436, mcs1_mcs_mat1_0_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_13537, new_AGEMA_signal_13536, mcs1_mcs_mat1_0_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_14017, new_AGEMA_signal_14016, mcs1_mcs_mat1_0_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_13537, new_AGEMA_signal_13536, mcs1_mcs_mat1_0_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({new_AGEMA_signal_10525, new_AGEMA_signal_10524, mcs1_mcs_mat1_0_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_9571, new_AGEMA_signal_9570, mcs1_mcs_mat1_0_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_8201, new_AGEMA_signal_8200, mcs1_mcs_mat1_0_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_10527, new_AGEMA_signal_10526, mcs1_mcs_mat1_0_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_7689, new_AGEMA_signal_7688, mcs1_mcs_mat1_0_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .c ({new_AGEMA_signal_8201, new_AGEMA_signal_8200, mcs1_mcs_mat1_0_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .c ({new_AGEMA_signal_8203, new_AGEMA_signal_8202, mcs1_mcs_mat1_0_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .c ({new_AGEMA_signal_9571, new_AGEMA_signal_9570, mcs1_mcs_mat1_0_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_7689, new_AGEMA_signal_7688, mcs1_mcs_mat1_0_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, mcs1_mcs_mat1_0_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_7689, new_AGEMA_signal_7688, mcs1_mcs_mat1_0_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .b ({new_AGEMA_signal_7691, new_AGEMA_signal_7690, mcs1_mcs_mat1_0_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_9581, new_AGEMA_signal_9580, mcs1_mcs_mat1_0_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({new_AGEMA_signal_7691, new_AGEMA_signal_7690, mcs1_mcs_mat1_0_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, mcs1_mcs_mat1_0_mcs_out[51]}), .c ({new_AGEMA_signal_10537, new_AGEMA_signal_10536, mcs1_mcs_mat1_0_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .c ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, mcs1_mcs_mat1_0_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_10539, new_AGEMA_signal_10538, mcs1_mcs_mat1_0_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_13047, new_AGEMA_signal_13046, mcs1_mcs_mat1_0_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_10539, new_AGEMA_signal_10538, mcs1_mcs_mat1_0_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_9587, new_AGEMA_signal_9586, mcs1_mcs_mat1_0_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_10543, new_AGEMA_signal_10542, mcs1_mcs_mat1_0_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .b ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_9587, new_AGEMA_signal_9586, mcs1_mcs_mat1_0_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_8937, new_AGEMA_signal_8936, mcs1_mcs_mat1_0_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_9589, new_AGEMA_signal_9588, mcs1_mcs_mat1_0_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .c ({new_AGEMA_signal_8937, new_AGEMA_signal_8936, mcs1_mcs_mat1_0_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({new_AGEMA_signal_7693, new_AGEMA_signal_7692, mcs1_mcs_mat1_0_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({new_AGEMA_signal_7695, new_AGEMA_signal_7694, mcs1_mcs_mat1_0_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_8941, new_AGEMA_signal_8940, mcs1_mcs_mat1_0_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .b ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_9595, new_AGEMA_signal_9594, mcs1_mcs_mat1_0_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_7695, new_AGEMA_signal_7694, mcs1_mcs_mat1_0_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_11519, new_AGEMA_signal_11518, mcs1_mcs_mat1_0_mcs_out[35]}), .b ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_12439, new_AGEMA_signal_12438, mcs1_mcs_mat1_0_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_10555, new_AGEMA_signal_10554, mcs1_mcs_mat1_0_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_7697, new_AGEMA_signal_7696, mcs1_mcs_mat1_0_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_11519, new_AGEMA_signal_11518, mcs1_mcs_mat1_0_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_9599, new_AGEMA_signal_9598, mcs1_mcs_mat1_0_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .c ({new_AGEMA_signal_10555, new_AGEMA_signal_10554, mcs1_mcs_mat1_0_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .c ({new_AGEMA_signal_9599, new_AGEMA_signal_9598, mcs1_mcs_mat1_0_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({new_AGEMA_signal_7697, new_AGEMA_signal_7696, mcs1_mcs_mat1_0_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_10557, new_AGEMA_signal_10556, mcs1_mcs_mat1_0_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_11521, new_AGEMA_signal_11520, mcs1_mcs_mat1_0_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({new_AGEMA_signal_13545, new_AGEMA_signal_13544, mcs1_mcs_mat1_0_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_14023, new_AGEMA_signal_14022, mcs1_mcs_mat1_0_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_10557, new_AGEMA_signal_10556, mcs1_mcs_mat1_0_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_13545, new_AGEMA_signal_13544, mcs1_mcs_mat1_0_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_10557, new_AGEMA_signal_10556, mcs1_mcs_mat1_0_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({new_AGEMA_signal_7699, new_AGEMA_signal_7698, mcs1_mcs_mat1_0_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_7701, new_AGEMA_signal_7700, mcs1_mcs_mat1_0_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_8953, new_AGEMA_signal_8952, mcs1_mcs_mat1_0_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, mcs1_mcs_mat1_0_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_8953, new_AGEMA_signal_8952, mcs1_mcs_mat1_0_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .c ({new_AGEMA_signal_9619, new_AGEMA_signal_9618, mcs1_mcs_mat1_0_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({new_AGEMA_signal_7703, new_AGEMA_signal_7702, mcs1_mcs_mat1_0_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_10577, new_AGEMA_signal_10576, mcs1_mcs_mat1_0_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({new_AGEMA_signal_7705, new_AGEMA_signal_7704, mcs1_mcs_mat1_0_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_7707, new_AGEMA_signal_7706, mcs1_mcs_mat1_0_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_8961, new_AGEMA_signal_8960, mcs1_mcs_mat1_0_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_7707, new_AGEMA_signal_7706, mcs1_mcs_mat1_0_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_8223, new_AGEMA_signal_8222, mcs1_mcs_mat1_0_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_7707, new_AGEMA_signal_7706, mcs1_mcs_mat1_0_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_9631, new_AGEMA_signal_9630, mcs1_mcs_mat1_0_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7709, new_AGEMA_signal_7708, mcs1_mcs_mat1_0_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_10585, new_AGEMA_signal_10584, mcs1_mcs_mat1_0_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_9631, new_AGEMA_signal_9630, mcs1_mcs_mat1_0_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .c ({new_AGEMA_signal_10589, new_AGEMA_signal_10588, mcs1_mcs_mat1_0_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_8965, new_AGEMA_signal_8964, mcs1_mcs_mat1_0_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_9631, new_AGEMA_signal_9630, mcs1_mcs_mat1_0_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_8965, new_AGEMA_signal_8964, mcs1_mcs_mat1_0_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .c ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, mcs1_mcs_mat1_0_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({new_AGEMA_signal_7709, new_AGEMA_signal_7708, mcs1_mcs_mat1_0_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U44 ( .a ({new_AGEMA_signal_8997, new_AGEMA_signal_8996, mcs1_mcs_mat1_1_mcs_out[90]}), .b ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, mcs1_mcs_mat1_1_mcs_out[94]}), .c ({new_AGEMA_signal_10595, new_AGEMA_signal_10594, mcs1_mcs_mat1_1_n93}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .c ({new_AGEMA_signal_8969, new_AGEMA_signal_8968, mcs1_mcs_mat1_1_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .b ({new_AGEMA_signal_7711, new_AGEMA_signal_7710, mcs1_mcs_mat1_1_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8229, new_AGEMA_signal_8228, mcs1_mcs_mat1_1_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_7711, new_AGEMA_signal_7710, mcs1_mcs_mat1_1_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_8975, new_AGEMA_signal_8974, mcs1_mcs_mat1_1_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_9641, new_AGEMA_signal_9640, mcs1_mcs_mat1_1_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_7713, new_AGEMA_signal_7712, mcs1_mcs_mat1_1_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_8975, new_AGEMA_signal_8974, mcs1_mcs_mat1_1_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({new_AGEMA_signal_7713, new_AGEMA_signal_7712, mcs1_mcs_mat1_1_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_10607, new_AGEMA_signal_10606, mcs1_mcs_mat1_1_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_13569, new_AGEMA_signal_13568, mcs1_mcs_mat1_1_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_14043, new_AGEMA_signal_14042, mcs1_mcs_mat1_1_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_11569, new_AGEMA_signal_11568, mcs1_mcs_mat1_1_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_13087, new_AGEMA_signal_13086, mcs1_mcs_mat1_1_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .c ({new_AGEMA_signal_11569, new_AGEMA_signal_11568, mcs1_mcs_mat1_1_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .b ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_13569, new_AGEMA_signal_13568, mcs1_mcs_mat1_1_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_10607, new_AGEMA_signal_10606, mcs1_mcs_mat1_1_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_9647, new_AGEMA_signal_9646, mcs1_mcs_mat1_1_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_10609, new_AGEMA_signal_10608, mcs1_mcs_mat1_1_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_7715, new_AGEMA_signal_7714, mcs1_mcs_mat1_1_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_9647, new_AGEMA_signal_9646, mcs1_mcs_mat1_1_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({new_AGEMA_signal_7715, new_AGEMA_signal_7714, mcs1_mcs_mat1_1_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_7717, new_AGEMA_signal_7716, mcs1_mcs_mat1_1_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({new_AGEMA_signal_8987, new_AGEMA_signal_8986, mcs1_mcs_mat1_1_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_9655, new_AGEMA_signal_9654, mcs1_mcs_mat1_1_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, mcs1_mcs_mat1_1_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_8987, new_AGEMA_signal_8986, mcs1_mcs_mat1_1_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .b ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .c ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, mcs1_mcs_mat1_1_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771]}), .c ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, mcs1_mcs_mat1_1_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_10623, new_AGEMA_signal_10622, mcs1_mcs_mat1_1_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_13091, new_AGEMA_signal_13090, mcs1_mcs_mat1_1_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_10623, new_AGEMA_signal_10622, mcs1_mcs_mat1_1_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .c ({new_AGEMA_signal_11589, new_AGEMA_signal_11588, mcs1_mcs_mat1_1_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_10623, new_AGEMA_signal_10622, mcs1_mcs_mat1_1_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_8991, new_AGEMA_signal_8990, mcs1_mcs_mat1_1_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .c ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, mcs1_mcs_mat1_1_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_7721, new_AGEMA_signal_7720, mcs1_mcs_mat1_1_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_8991, new_AGEMA_signal_8990, mcs1_mcs_mat1_1_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_8993, new_AGEMA_signal_8992, mcs1_mcs_mat1_1_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777]}), .c ({new_AGEMA_signal_7721, new_AGEMA_signal_7720, mcs1_mcs_mat1_1_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .b ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .c ({new_AGEMA_signal_8997, new_AGEMA_signal_8996, mcs1_mcs_mat1_1_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .b ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_8999, new_AGEMA_signal_8998, mcs1_mcs_mat1_1_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, mcs1_mcs_mat1_1_mcs_out[87]}), .c ({new_AGEMA_signal_10627, new_AGEMA_signal_10626, mcs1_mcs_mat1_1_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .c ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, mcs1_mcs_mat1_1_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .c ({new_AGEMA_signal_13579, new_AGEMA_signal_13578, mcs1_mcs_mat1_1_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_10629, new_AGEMA_signal_10628, mcs1_mcs_mat1_1_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_7723, new_AGEMA_signal_7722, mcs1_mcs_mat1_1_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_8243, new_AGEMA_signal_8242, mcs1_mcs_mat1_1_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783]}), .c ({new_AGEMA_signal_7723, new_AGEMA_signal_7722, mcs1_mcs_mat1_1_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_7725, new_AGEMA_signal_7724, mcs1_mcs_mat1_1_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_8247, new_AGEMA_signal_8246, mcs1_mcs_mat1_1_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_7725, new_AGEMA_signal_7724, mcs1_mcs_mat1_1_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789]}), .c ({new_AGEMA_signal_7727, new_AGEMA_signal_7726, mcs1_mcs_mat1_1_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_10641, new_AGEMA_signal_10640, mcs1_mcs_mat1_1_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .c ({new_AGEMA_signal_13583, new_AGEMA_signal_13582, mcs1_mcs_mat1_1_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_10641, new_AGEMA_signal_10640, mcs1_mcs_mat1_1_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_11617, new_AGEMA_signal_11616, mcs1_mcs_mat1_1_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_7729, new_AGEMA_signal_7728, mcs1_mcs_mat1_1_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_12507, new_AGEMA_signal_12506, mcs1_mcs_mat1_1_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_10647, new_AGEMA_signal_10646, mcs1_mcs_mat1_1_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_11617, new_AGEMA_signal_11616, mcs1_mcs_mat1_1_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, mcs1_mcs_mat1_1_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_10647, new_AGEMA_signal_10646, mcs1_mcs_mat1_1_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, mcs1_mcs_mat1_1_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795]}), .c ({new_AGEMA_signal_7729, new_AGEMA_signal_7728, mcs1_mcs_mat1_1_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, mcs1_mcs_mat1_1_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_8255, new_AGEMA_signal_8254, mcs1_mcs_mat1_1_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_10649, new_AGEMA_signal_10648, mcs1_mcs_mat1_1_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_7731, new_AGEMA_signal_7730, mcs1_mcs_mat1_1_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .c ({new_AGEMA_signal_8255, new_AGEMA_signal_8254, mcs1_mcs_mat1_1_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .c ({new_AGEMA_signal_8257, new_AGEMA_signal_8256, mcs1_mcs_mat1_1_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .c ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, mcs1_mcs_mat1_1_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_7731, new_AGEMA_signal_7730, mcs1_mcs_mat1_1_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_9695, new_AGEMA_signal_9694, mcs1_mcs_mat1_1_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_7731, new_AGEMA_signal_7730, mcs1_mcs_mat1_1_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .b ({new_AGEMA_signal_7733, new_AGEMA_signal_7732, mcs1_mcs_mat1_1_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_9703, new_AGEMA_signal_9702, mcs1_mcs_mat1_1_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801]}), .c ({new_AGEMA_signal_7733, new_AGEMA_signal_7732, mcs1_mcs_mat1_1_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({new_AGEMA_signal_13587, new_AGEMA_signal_13586, mcs1_mcs_mat1_1_mcs_out[51]}), .c ({new_AGEMA_signal_14061, new_AGEMA_signal_14060, mcs1_mcs_mat1_1_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .c ({new_AGEMA_signal_13587, new_AGEMA_signal_13586, mcs1_mcs_mat1_1_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_7735, new_AGEMA_signal_7734, mcs1_mcs_mat1_1_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_9015, new_AGEMA_signal_9014, mcs1_mcs_mat1_1_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_7735, new_AGEMA_signal_7734, mcs1_mcs_mat1_1_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, mcs1_mcs_mat1_1_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_10663, new_AGEMA_signal_10662, mcs1_mcs_mat1_1_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .b ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, mcs1_mcs_mat1_1_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_9019, new_AGEMA_signal_9018, mcs1_mcs_mat1_1_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_9713, new_AGEMA_signal_9712, mcs1_mcs_mat1_1_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .c ({new_AGEMA_signal_9019, new_AGEMA_signal_9018, mcs1_mcs_mat1_1_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807]}), .c ({new_AGEMA_signal_7737, new_AGEMA_signal_7736, mcs1_mcs_mat1_1_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({new_AGEMA_signal_7739, new_AGEMA_signal_7738, mcs1_mcs_mat1_1_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9023, new_AGEMA_signal_9022, mcs1_mcs_mat1_1_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .b ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_9719, new_AGEMA_signal_9718, mcs1_mcs_mat1_1_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_7739, new_AGEMA_signal_7738, mcs1_mcs_mat1_1_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_14493, new_AGEMA_signal_14492, mcs1_mcs_mat1_1_mcs_out[35]}), .b ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_14981, new_AGEMA_signal_14980, mcs1_mcs_mat1_1_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_14065, new_AGEMA_signal_14064, mcs1_mcs_mat1_1_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_10673, new_AGEMA_signal_10672, mcs1_mcs_mat1_1_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_14493, new_AGEMA_signal_14492, mcs1_mcs_mat1_1_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_13589, new_AGEMA_signal_13588, mcs1_mcs_mat1_1_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .c ({new_AGEMA_signal_14065, new_AGEMA_signal_14064, mcs1_mcs_mat1_1_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .c ({new_AGEMA_signal_13589, new_AGEMA_signal_13588, mcs1_mcs_mat1_1_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813]}), .c ({new_AGEMA_signal_10673, new_AGEMA_signal_10672, mcs1_mcs_mat1_1_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_7741, new_AGEMA_signal_7740, mcs1_mcs_mat1_1_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_8269, new_AGEMA_signal_8268, mcs1_mcs_mat1_1_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, mcs1_mcs_mat1_1_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_10677, new_AGEMA_signal_10676, mcs1_mcs_mat1_1_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_7741, new_AGEMA_signal_7740, mcs1_mcs_mat1_1_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, mcs1_mcs_mat1_1_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_7741, new_AGEMA_signal_7740, mcs1_mcs_mat1_1_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819]}), .c ({new_AGEMA_signal_7743, new_AGEMA_signal_7742, mcs1_mcs_mat1_1_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_7745, new_AGEMA_signal_7744, mcs1_mcs_mat1_1_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_13103, new_AGEMA_signal_13102, mcs1_mcs_mat1_1_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_13593, new_AGEMA_signal_13592, mcs1_mcs_mat1_1_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_13103, new_AGEMA_signal_13102, mcs1_mcs_mat1_1_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .c ({new_AGEMA_signal_13597, new_AGEMA_signal_13596, mcs1_mcs_mat1_1_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825]}), .c ({new_AGEMA_signal_10693, new_AGEMA_signal_10692, mcs1_mcs_mat1_1_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_7747, new_AGEMA_signal_7746, mcs1_mcs_mat1_1_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831]}), .c ({new_AGEMA_signal_7749, new_AGEMA_signal_7748, mcs1_mcs_mat1_1_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_7751, new_AGEMA_signal_7750, mcs1_mcs_mat1_1_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_9041, new_AGEMA_signal_9040, mcs1_mcs_mat1_1_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_7751, new_AGEMA_signal_7750, mcs1_mcs_mat1_1_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_8281, new_AGEMA_signal_8280, mcs1_mcs_mat1_1_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_7751, new_AGEMA_signal_7750, mcs1_mcs_mat1_1_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_13605, new_AGEMA_signal_13604, mcs1_mcs_mat1_1_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_10707, new_AGEMA_signal_10706, mcs1_mcs_mat1_1_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_14073, new_AGEMA_signal_14072, mcs1_mcs_mat1_1_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_13605, new_AGEMA_signal_13604, mcs1_mcs_mat1_1_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .c ({new_AGEMA_signal_14077, new_AGEMA_signal_14076, mcs1_mcs_mat1_1_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_13111, new_AGEMA_signal_13110, mcs1_mcs_mat1_1_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_13605, new_AGEMA_signal_13604, mcs1_mcs_mat1_1_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_13111, new_AGEMA_signal_13110, mcs1_mcs_mat1_1_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .c ({new_AGEMA_signal_13607, new_AGEMA_signal_13606, mcs1_mcs_mat1_1_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837]}), .c ({new_AGEMA_signal_10707, new_AGEMA_signal_10706, mcs1_mcs_mat1_1_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U44 ( .a ({new_AGEMA_signal_9071, new_AGEMA_signal_9070, mcs1_mcs_mat1_2_mcs_out[90]}), .b ({new_AGEMA_signal_9771, new_AGEMA_signal_9770, mcs1_mcs_mat1_2_mcs_out[94]}), .c ({new_AGEMA_signal_10711, new_AGEMA_signal_10710, mcs1_mcs_mat1_2_n93}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .c ({new_AGEMA_signal_9045, new_AGEMA_signal_9044, mcs1_mcs_mat1_2_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .b ({new_AGEMA_signal_7753, new_AGEMA_signal_7752, mcs1_mcs_mat1_2_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8285, new_AGEMA_signal_8284, mcs1_mcs_mat1_2_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_7753, new_AGEMA_signal_7752, mcs1_mcs_mat1_2_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, mcs1_mcs_mat1_2_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_13619, new_AGEMA_signal_13618, mcs1_mcs_mat1_2_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_10719, new_AGEMA_signal_10718, mcs1_mcs_mat1_2_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, mcs1_mcs_mat1_2_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843]}), .c ({new_AGEMA_signal_10719, new_AGEMA_signal_10718, mcs1_mcs_mat1_2_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_7755, new_AGEMA_signal_7754, mcs1_mcs_mat1_2_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9757, new_AGEMA_signal_9756, mcs1_mcs_mat1_2_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_10721, new_AGEMA_signal_10720, mcs1_mcs_mat1_2_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_8289, new_AGEMA_signal_8288, mcs1_mcs_mat1_2_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_9051, new_AGEMA_signal_9050, mcs1_mcs_mat1_2_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .c ({new_AGEMA_signal_8289, new_AGEMA_signal_8288, mcs1_mcs_mat1_2_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .b ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_9757, new_AGEMA_signal_9756, mcs1_mcs_mat1_2_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_7755, new_AGEMA_signal_7754, mcs1_mcs_mat1_2_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_9761, new_AGEMA_signal_9760, mcs1_mcs_mat1_2_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_10727, new_AGEMA_signal_10726, mcs1_mcs_mat1_2_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_7757, new_AGEMA_signal_7756, mcs1_mcs_mat1_2_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_9761, new_AGEMA_signal_9760, mcs1_mcs_mat1_2_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849]}), .c ({new_AGEMA_signal_7757, new_AGEMA_signal_7756, mcs1_mcs_mat1_2_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_7759, new_AGEMA_signal_7758, mcs1_mcs_mat1_2_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, mcs1_mcs_mat1_2_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_13625, new_AGEMA_signal_13624, mcs1_mcs_mat1_2_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_10735, new_AGEMA_signal_10734, mcs1_mcs_mat1_2_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, mcs1_mcs_mat1_2_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .b ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .c ({new_AGEMA_signal_13627, new_AGEMA_signal_13626, mcs1_mcs_mat1_2_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855]}), .c ({new_AGEMA_signal_10735, new_AGEMA_signal_10734, mcs1_mcs_mat1_2_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_7761, new_AGEMA_signal_7760, mcs1_mcs_mat1_2_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_9061, new_AGEMA_signal_9060, mcs1_mcs_mat1_2_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_7761, new_AGEMA_signal_7760, mcs1_mcs_mat1_2_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .c ({new_AGEMA_signal_8297, new_AGEMA_signal_8296, mcs1_mcs_mat1_2_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_7761, new_AGEMA_signal_7760, mcs1_mcs_mat1_2_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_9065, new_AGEMA_signal_9064, mcs1_mcs_mat1_2_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .c ({new_AGEMA_signal_9771, new_AGEMA_signal_9770, mcs1_mcs_mat1_2_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_7763, new_AGEMA_signal_7762, mcs1_mcs_mat1_2_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_9065, new_AGEMA_signal_9064, mcs1_mcs_mat1_2_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_9067, new_AGEMA_signal_9066, mcs1_mcs_mat1_2_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861]}), .c ({new_AGEMA_signal_7763, new_AGEMA_signal_7762, mcs1_mcs_mat1_2_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .b ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .c ({new_AGEMA_signal_9071, new_AGEMA_signal_9070, mcs1_mcs_mat1_2_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .b ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_9073, new_AGEMA_signal_9072, mcs1_mcs_mat1_2_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({new_AGEMA_signal_13635, new_AGEMA_signal_13634, mcs1_mcs_mat1_2_mcs_out[87]}), .c ({new_AGEMA_signal_14101, new_AGEMA_signal_14100, mcs1_mcs_mat1_2_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .c ({new_AGEMA_signal_13635, new_AGEMA_signal_13634, mcs1_mcs_mat1_2_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .c ({new_AGEMA_signal_9781, new_AGEMA_signal_9780, mcs1_mcs_mat1_2_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_7765, new_AGEMA_signal_7764, mcs1_mcs_mat1_2_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_7767, new_AGEMA_signal_7766, mcs1_mcs_mat1_2_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_8305, new_AGEMA_signal_8304, mcs1_mcs_mat1_2_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867]}), .c ({new_AGEMA_signal_7767, new_AGEMA_signal_7766, mcs1_mcs_mat1_2_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_7769, new_AGEMA_signal_7768, mcs1_mcs_mat1_2_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_8309, new_AGEMA_signal_8308, mcs1_mcs_mat1_2_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_7769, new_AGEMA_signal_7768, mcs1_mcs_mat1_2_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873]}), .c ({new_AGEMA_signal_10755, new_AGEMA_signal_10754, mcs1_mcs_mat1_2_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_7771, new_AGEMA_signal_7770, mcs1_mcs_mat1_2_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .c ({new_AGEMA_signal_9795, new_AGEMA_signal_9794, mcs1_mcs_mat1_2_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_7771, new_AGEMA_signal_7770, mcs1_mcs_mat1_2_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_11727, new_AGEMA_signal_11726, mcs1_mcs_mat1_2_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_7773, new_AGEMA_signal_7772, mcs1_mcs_mat1_2_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_12589, new_AGEMA_signal_12588, mcs1_mcs_mat1_2_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_10763, new_AGEMA_signal_10762, mcs1_mcs_mat1_2_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_11727, new_AGEMA_signal_11726, mcs1_mcs_mat1_2_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_9799, new_AGEMA_signal_9798, mcs1_mcs_mat1_2_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_10763, new_AGEMA_signal_10762, mcs1_mcs_mat1_2_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_9799, new_AGEMA_signal_9798, mcs1_mcs_mat1_2_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879]}), .c ({new_AGEMA_signal_7773, new_AGEMA_signal_7772, mcs1_mcs_mat1_2_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_9805, new_AGEMA_signal_9804, mcs1_mcs_mat1_2_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_8317, new_AGEMA_signal_8316, mcs1_mcs_mat1_2_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_10765, new_AGEMA_signal_10764, mcs1_mcs_mat1_2_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_7775, new_AGEMA_signal_7774, mcs1_mcs_mat1_2_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .c ({new_AGEMA_signal_8317, new_AGEMA_signal_8316, mcs1_mcs_mat1_2_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .c ({new_AGEMA_signal_8319, new_AGEMA_signal_8318, mcs1_mcs_mat1_2_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .c ({new_AGEMA_signal_9805, new_AGEMA_signal_9804, mcs1_mcs_mat1_2_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_7775, new_AGEMA_signal_7774, mcs1_mcs_mat1_2_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_9807, new_AGEMA_signal_9806, mcs1_mcs_mat1_2_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_7775, new_AGEMA_signal_7774, mcs1_mcs_mat1_2_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .b ({new_AGEMA_signal_10771, new_AGEMA_signal_10770, mcs1_mcs_mat1_2_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_13647, new_AGEMA_signal_13646, mcs1_mcs_mat1_2_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885]}), .c ({new_AGEMA_signal_10771, new_AGEMA_signal_10770, mcs1_mcs_mat1_2_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({new_AGEMA_signal_9811, new_AGEMA_signal_9810, mcs1_mcs_mat1_2_mcs_out[51]}), .c ({new_AGEMA_signal_10773, new_AGEMA_signal_10772, mcs1_mcs_mat1_2_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .c ({new_AGEMA_signal_9811, new_AGEMA_signal_9810, mcs1_mcs_mat1_2_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_7777, new_AGEMA_signal_7776, mcs1_mcs_mat1_2_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_9087, new_AGEMA_signal_9086, mcs1_mcs_mat1_2_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_7777, new_AGEMA_signal_7776, mcs1_mcs_mat1_2_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_9817, new_AGEMA_signal_9816, mcs1_mcs_mat1_2_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_10779, new_AGEMA_signal_10778, mcs1_mcs_mat1_2_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .b ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_9817, new_AGEMA_signal_9816, mcs1_mcs_mat1_2_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_9091, new_AGEMA_signal_9090, mcs1_mcs_mat1_2_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_9819, new_AGEMA_signal_9818, mcs1_mcs_mat1_2_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .c ({new_AGEMA_signal_9091, new_AGEMA_signal_9090, mcs1_mcs_mat1_2_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891]}), .c ({new_AGEMA_signal_7779, new_AGEMA_signal_7778, mcs1_mcs_mat1_2_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({new_AGEMA_signal_10785, new_AGEMA_signal_10784, mcs1_mcs_mat1_2_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_13165, new_AGEMA_signal_13164, mcs1_mcs_mat1_2_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .b ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_13653, new_AGEMA_signal_13652, mcs1_mcs_mat1_2_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_10785, new_AGEMA_signal_10784, mcs1_mcs_mat1_2_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_11743, new_AGEMA_signal_11742, mcs1_mcs_mat1_2_mcs_out[35]}), .b ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_12595, new_AGEMA_signal_12594, mcs1_mcs_mat1_2_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_10789, new_AGEMA_signal_10788, mcs1_mcs_mat1_2_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_7781, new_AGEMA_signal_7780, mcs1_mcs_mat1_2_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_11743, new_AGEMA_signal_11742, mcs1_mcs_mat1_2_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_9823, new_AGEMA_signal_9822, mcs1_mcs_mat1_2_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .c ({new_AGEMA_signal_10789, new_AGEMA_signal_10788, mcs1_mcs_mat1_2_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .c ({new_AGEMA_signal_9823, new_AGEMA_signal_9822, mcs1_mcs_mat1_2_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897]}), .c ({new_AGEMA_signal_7781, new_AGEMA_signal_7780, mcs1_mcs_mat1_2_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_7783, new_AGEMA_signal_7782, mcs1_mcs_mat1_2_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_8329, new_AGEMA_signal_8328, mcs1_mcs_mat1_2_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({new_AGEMA_signal_9827, new_AGEMA_signal_9826, mcs1_mcs_mat1_2_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_10793, new_AGEMA_signal_10792, mcs1_mcs_mat1_2_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_7783, new_AGEMA_signal_7782, mcs1_mcs_mat1_2_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_9827, new_AGEMA_signal_9826, mcs1_mcs_mat1_2_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_7783, new_AGEMA_signal_7782, mcs1_mcs_mat1_2_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903]}), .c ({new_AGEMA_signal_7785, new_AGEMA_signal_7784, mcs1_mcs_mat1_2_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_10803, new_AGEMA_signal_10802, mcs1_mcs_mat1_2_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_9101, new_AGEMA_signal_9100, mcs1_mcs_mat1_2_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_9839, new_AGEMA_signal_9838, mcs1_mcs_mat1_2_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_9101, new_AGEMA_signal_9100, mcs1_mcs_mat1_2_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .c ({new_AGEMA_signal_9843, new_AGEMA_signal_9842, mcs1_mcs_mat1_2_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909]}), .c ({new_AGEMA_signal_7787, new_AGEMA_signal_7786, mcs1_mcs_mat1_2_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_7789, new_AGEMA_signal_7788, mcs1_mcs_mat1_2_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915]}), .c ({new_AGEMA_signal_7791, new_AGEMA_signal_7790, mcs1_mcs_mat1_2_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_10821, new_AGEMA_signal_10820, mcs1_mcs_mat1_2_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_13177, new_AGEMA_signal_13176, mcs1_mcs_mat1_2_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_10821, new_AGEMA_signal_10820, mcs1_mcs_mat1_2_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_11771, new_AGEMA_signal_11770, mcs1_mcs_mat1_2_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_10821, new_AGEMA_signal_10820, mcs1_mcs_mat1_2_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_9857, new_AGEMA_signal_9856, mcs1_mcs_mat1_2_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7793, new_AGEMA_signal_7792, mcs1_mcs_mat1_2_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_10823, new_AGEMA_signal_10822, mcs1_mcs_mat1_2_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_9857, new_AGEMA_signal_9856, mcs1_mcs_mat1_2_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .c ({new_AGEMA_signal_10827, new_AGEMA_signal_10826, mcs1_mcs_mat1_2_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_9111, new_AGEMA_signal_9110, mcs1_mcs_mat1_2_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_9857, new_AGEMA_signal_9856, mcs1_mcs_mat1_2_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_9111, new_AGEMA_signal_9110, mcs1_mcs_mat1_2_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .c ({new_AGEMA_signal_9859, new_AGEMA_signal_9858, mcs1_mcs_mat1_2_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921]}), .c ({new_AGEMA_signal_7793, new_AGEMA_signal_7792, mcs1_mcs_mat1_2_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U44 ( .a ({new_AGEMA_signal_13223, new_AGEMA_signal_13222, mcs1_mcs_mat1_3_mcs_out[90]}), .b ({new_AGEMA_signal_9889, new_AGEMA_signal_9888, mcs1_mcs_mat1_3_mcs_out[94]}), .c ({new_AGEMA_signal_13671, new_AGEMA_signal_13670, mcs1_mcs_mat1_3_n93}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .c ({new_AGEMA_signal_9115, new_AGEMA_signal_9114, mcs1_mcs_mat1_3_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .b ({new_AGEMA_signal_10831, new_AGEMA_signal_10830, mcs1_mcs_mat1_3_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, mcs1_mcs_mat1_3_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_10831, new_AGEMA_signal_10830, mcs1_mcs_mat1_3_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_9117, new_AGEMA_signal_9116, mcs1_mcs_mat1_3_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_9863, new_AGEMA_signal_9862, mcs1_mcs_mat1_3_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_7795, new_AGEMA_signal_7794, mcs1_mcs_mat1_3_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_9117, new_AGEMA_signal_9116, mcs1_mcs_mat1_3_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927]}), .c ({new_AGEMA_signal_7795, new_AGEMA_signal_7794, mcs1_mcs_mat1_3_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_7797, new_AGEMA_signal_7796, mcs1_mcs_mat1_3_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9871, new_AGEMA_signal_9870, mcs1_mcs_mat1_3_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_10837, new_AGEMA_signal_10836, mcs1_mcs_mat1_3_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_8345, new_AGEMA_signal_8344, mcs1_mcs_mat1_3_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_9123, new_AGEMA_signal_9122, mcs1_mcs_mat1_3_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .c ({new_AGEMA_signal_8345, new_AGEMA_signal_8344, mcs1_mcs_mat1_3_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .b ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_9871, new_AGEMA_signal_9870, mcs1_mcs_mat1_3_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_7797, new_AGEMA_signal_7796, mcs1_mcs_mat1_3_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_9875, new_AGEMA_signal_9874, mcs1_mcs_mat1_3_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_10843, new_AGEMA_signal_10842, mcs1_mcs_mat1_3_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_7799, new_AGEMA_signal_7798, mcs1_mcs_mat1_3_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_9875, new_AGEMA_signal_9874, mcs1_mcs_mat1_3_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933]}), .c ({new_AGEMA_signal_7799, new_AGEMA_signal_7798, mcs1_mcs_mat1_3_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_10847, new_AGEMA_signal_10846, mcs1_mcs_mat1_3_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({new_AGEMA_signal_9129, new_AGEMA_signal_9128, mcs1_mcs_mat1_3_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_9879, new_AGEMA_signal_9878, mcs1_mcs_mat1_3_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_7801, new_AGEMA_signal_7800, mcs1_mcs_mat1_3_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_9129, new_AGEMA_signal_9128, mcs1_mcs_mat1_3_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .b ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .c ({new_AGEMA_signal_9881, new_AGEMA_signal_9880, mcs1_mcs_mat1_3_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939]}), .c ({new_AGEMA_signal_7801, new_AGEMA_signal_7800, mcs1_mcs_mat1_3_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_7803, new_AGEMA_signal_7802, mcs1_mcs_mat1_3_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_9133, new_AGEMA_signal_9132, mcs1_mcs_mat1_3_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_7803, new_AGEMA_signal_7802, mcs1_mcs_mat1_3_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .c ({new_AGEMA_signal_8353, new_AGEMA_signal_8352, mcs1_mcs_mat1_3_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_7803, new_AGEMA_signal_7802, mcs1_mcs_mat1_3_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_9137, new_AGEMA_signal_9136, mcs1_mcs_mat1_3_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .c ({new_AGEMA_signal_9889, new_AGEMA_signal_9888, mcs1_mcs_mat1_3_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_7805, new_AGEMA_signal_7804, mcs1_mcs_mat1_3_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_9137, new_AGEMA_signal_9136, mcs1_mcs_mat1_3_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_9139, new_AGEMA_signal_9138, mcs1_mcs_mat1_3_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945]}), .c ({new_AGEMA_signal_7805, new_AGEMA_signal_7804, mcs1_mcs_mat1_3_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .b ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .c ({new_AGEMA_signal_13223, new_AGEMA_signal_13222, mcs1_mcs_mat1_3_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .b ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_13225, new_AGEMA_signal_13224, mcs1_mcs_mat1_3_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({new_AGEMA_signal_9895, new_AGEMA_signal_9894, mcs1_mcs_mat1_3_mcs_out[87]}), .c ({new_AGEMA_signal_10859, new_AGEMA_signal_10858, mcs1_mcs_mat1_3_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .c ({new_AGEMA_signal_9895, new_AGEMA_signal_9894, mcs1_mcs_mat1_3_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .c ({new_AGEMA_signal_9901, new_AGEMA_signal_9900, mcs1_mcs_mat1_3_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_7807, new_AGEMA_signal_7806, mcs1_mcs_mat1_3_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_7809, new_AGEMA_signal_7808, mcs1_mcs_mat1_3_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_8361, new_AGEMA_signal_8360, mcs1_mcs_mat1_3_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951]}), .c ({new_AGEMA_signal_7809, new_AGEMA_signal_7808, mcs1_mcs_mat1_3_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_10871, new_AGEMA_signal_10870, mcs1_mcs_mat1_3_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_11829, new_AGEMA_signal_11828, mcs1_mcs_mat1_3_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_10871, new_AGEMA_signal_10870, mcs1_mcs_mat1_3_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957]}), .c ({new_AGEMA_signal_7811, new_AGEMA_signal_7810, mcs1_mcs_mat1_3_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_7813, new_AGEMA_signal_7812, mcs1_mcs_mat1_3_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .c ({new_AGEMA_signal_9915, new_AGEMA_signal_9914, mcs1_mcs_mat1_3_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_7813, new_AGEMA_signal_7812, mcs1_mcs_mat1_3_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_11845, new_AGEMA_signal_11844, mcs1_mcs_mat1_3_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_7815, new_AGEMA_signal_7814, mcs1_mcs_mat1_3_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_12653, new_AGEMA_signal_12652, mcs1_mcs_mat1_3_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_10883, new_AGEMA_signal_10882, mcs1_mcs_mat1_3_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_11845, new_AGEMA_signal_11844, mcs1_mcs_mat1_3_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_9919, new_AGEMA_signal_9918, mcs1_mcs_mat1_3_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_10883, new_AGEMA_signal_10882, mcs1_mcs_mat1_3_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_9919, new_AGEMA_signal_9918, mcs1_mcs_mat1_3_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963]}), .c ({new_AGEMA_signal_7815, new_AGEMA_signal_7814, mcs1_mcs_mat1_3_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_13699, new_AGEMA_signal_13698, mcs1_mcs_mat1_3_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, mcs1_mcs_mat1_3_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_14151, new_AGEMA_signal_14150, mcs1_mcs_mat1_3_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_10885, new_AGEMA_signal_10884, mcs1_mcs_mat1_3_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .c ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, mcs1_mcs_mat1_3_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .c ({new_AGEMA_signal_11849, new_AGEMA_signal_11848, mcs1_mcs_mat1_3_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .c ({new_AGEMA_signal_13699, new_AGEMA_signal_13698, mcs1_mcs_mat1_3_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_10885, new_AGEMA_signal_10884, mcs1_mcs_mat1_3_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_13701, new_AGEMA_signal_13700, mcs1_mcs_mat1_3_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_10885, new_AGEMA_signal_10884, mcs1_mcs_mat1_3_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .b ({new_AGEMA_signal_7817, new_AGEMA_signal_7816, mcs1_mcs_mat1_3_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_9927, new_AGEMA_signal_9926, mcs1_mcs_mat1_3_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969]}), .c ({new_AGEMA_signal_7817, new_AGEMA_signal_7816, mcs1_mcs_mat1_3_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({new_AGEMA_signal_9931, new_AGEMA_signal_9930, mcs1_mcs_mat1_3_mcs_out[51]}), .c ({new_AGEMA_signal_10891, new_AGEMA_signal_10890, mcs1_mcs_mat1_3_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .c ({new_AGEMA_signal_9931, new_AGEMA_signal_9930, mcs1_mcs_mat1_3_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_7819, new_AGEMA_signal_7818, mcs1_mcs_mat1_3_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_9157, new_AGEMA_signal_9156, mcs1_mcs_mat1_3_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_7819, new_AGEMA_signal_7818, mcs1_mcs_mat1_3_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_13705, new_AGEMA_signal_13704, mcs1_mcs_mat1_3_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_14159, new_AGEMA_signal_14158, mcs1_mcs_mat1_3_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .b ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_13705, new_AGEMA_signal_13704, mcs1_mcs_mat1_3_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_13235, new_AGEMA_signal_13234, mcs1_mcs_mat1_3_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_13707, new_AGEMA_signal_13706, mcs1_mcs_mat1_3_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .c ({new_AGEMA_signal_13235, new_AGEMA_signal_13234, mcs1_mcs_mat1_3_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975]}), .c ({new_AGEMA_signal_10895, new_AGEMA_signal_10894, mcs1_mcs_mat1_3_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({new_AGEMA_signal_7821, new_AGEMA_signal_7820, mcs1_mcs_mat1_3_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9161, new_AGEMA_signal_9160, mcs1_mcs_mat1_3_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .b ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_9939, new_AGEMA_signal_9938, mcs1_mcs_mat1_3_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_7821, new_AGEMA_signal_7820, mcs1_mcs_mat1_3_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_11865, new_AGEMA_signal_11864, mcs1_mcs_mat1_3_mcs_out[35]}), .b ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_12665, new_AGEMA_signal_12664, mcs1_mcs_mat1_3_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_10903, new_AGEMA_signal_10902, mcs1_mcs_mat1_3_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_7823, new_AGEMA_signal_7822, mcs1_mcs_mat1_3_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_11865, new_AGEMA_signal_11864, mcs1_mcs_mat1_3_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_9943, new_AGEMA_signal_9942, mcs1_mcs_mat1_3_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .c ({new_AGEMA_signal_10903, new_AGEMA_signal_10902, mcs1_mcs_mat1_3_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .c ({new_AGEMA_signal_9943, new_AGEMA_signal_9942, mcs1_mcs_mat1_3_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981]}), .c ({new_AGEMA_signal_7823, new_AGEMA_signal_7822, mcs1_mcs_mat1_3_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_7825, new_AGEMA_signal_7824, mcs1_mcs_mat1_3_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_8379, new_AGEMA_signal_8378, mcs1_mcs_mat1_3_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({new_AGEMA_signal_9947, new_AGEMA_signal_9946, mcs1_mcs_mat1_3_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_10907, new_AGEMA_signal_10906, mcs1_mcs_mat1_3_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_7825, new_AGEMA_signal_7824, mcs1_mcs_mat1_3_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_9947, new_AGEMA_signal_9946, mcs1_mcs_mat1_3_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_7825, new_AGEMA_signal_7824, mcs1_mcs_mat1_3_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987]}), .c ({new_AGEMA_signal_10911, new_AGEMA_signal_10910, mcs1_mcs_mat1_3_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_7827, new_AGEMA_signal_7826, mcs1_mcs_mat1_3_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_9173, new_AGEMA_signal_9172, mcs1_mcs_mat1_3_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_9959, new_AGEMA_signal_9958, mcs1_mcs_mat1_3_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_9173, new_AGEMA_signal_9172, mcs1_mcs_mat1_3_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .c ({new_AGEMA_signal_9963, new_AGEMA_signal_9962, mcs1_mcs_mat1_3_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993]}), .c ({new_AGEMA_signal_7829, new_AGEMA_signal_7828, mcs1_mcs_mat1_3_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_7831, new_AGEMA_signal_7830, mcs1_mcs_mat1_3_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999]}), .c ({new_AGEMA_signal_10931, new_AGEMA_signal_10930, mcs1_mcs_mat1_3_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_7833, new_AGEMA_signal_7832, mcs1_mcs_mat1_3_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_9179, new_AGEMA_signal_9178, mcs1_mcs_mat1_3_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_7833, new_AGEMA_signal_7832, mcs1_mcs_mat1_3_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, mcs1_mcs_mat1_3_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_7833, new_AGEMA_signal_7832, mcs1_mcs_mat1_3_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, mcs1_mcs_mat1_3_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7835, new_AGEMA_signal_7834, mcs1_mcs_mat1_3_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_10935, new_AGEMA_signal_10934, mcs1_mcs_mat1_3_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, mcs1_mcs_mat1_3_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .c ({new_AGEMA_signal_10939, new_AGEMA_signal_10938, mcs1_mcs_mat1_3_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_9183, new_AGEMA_signal_9182, mcs1_mcs_mat1_3_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, mcs1_mcs_mat1_3_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_9183, new_AGEMA_signal_9182, mcs1_mcs_mat1_3_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .c ({new_AGEMA_signal_9977, new_AGEMA_signal_9976, mcs1_mcs_mat1_3_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005]}), .c ({new_AGEMA_signal_7835, new_AGEMA_signal_7834, mcs1_mcs_mat1_3_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U44 ( .a ({new_AGEMA_signal_9213, new_AGEMA_signal_9212, mcs1_mcs_mat1_4_mcs_out[90]}), .b ({new_AGEMA_signal_13745, new_AGEMA_signal_13744, mcs1_mcs_mat1_4_mcs_out[94]}), .c ({new_AGEMA_signal_14181, new_AGEMA_signal_14180, mcs1_mcs_mat1_4_n93}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .c ({new_AGEMA_signal_13283, new_AGEMA_signal_13282, mcs1_mcs_mat1_4_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .b ({new_AGEMA_signal_7837, new_AGEMA_signal_7836, mcs1_mcs_mat1_4_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, mcs1_mcs_mat1_4_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_7837, new_AGEMA_signal_7836, mcs1_mcs_mat1_4_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_9191, new_AGEMA_signal_9190, mcs1_mcs_mat1_4_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_9985, new_AGEMA_signal_9984, mcs1_mcs_mat1_4_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_7839, new_AGEMA_signal_7838, mcs1_mcs_mat1_4_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_9191, new_AGEMA_signal_9190, mcs1_mcs_mat1_4_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011]}), .c ({new_AGEMA_signal_7839, new_AGEMA_signal_7838, mcs1_mcs_mat1_4_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_7841, new_AGEMA_signal_7840, mcs1_mcs_mat1_4_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, mcs1_mcs_mat1_4_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_10951, new_AGEMA_signal_10950, mcs1_mcs_mat1_4_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, mcs1_mcs_mat1_4_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_9197, new_AGEMA_signal_9196, mcs1_mcs_mat1_4_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .c ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, mcs1_mcs_mat1_4_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .b ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, mcs1_mcs_mat1_4_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_7841, new_AGEMA_signal_7840, mcs1_mcs_mat1_4_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_13739, new_AGEMA_signal_13738, mcs1_mcs_mat1_4_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_14191, new_AGEMA_signal_14190, mcs1_mcs_mat1_4_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_10957, new_AGEMA_signal_10956, mcs1_mcs_mat1_4_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_13739, new_AGEMA_signal_13738, mcs1_mcs_mat1_4_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017]}), .c ({new_AGEMA_signal_10957, new_AGEMA_signal_10956, mcs1_mcs_mat1_4_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_7843, new_AGEMA_signal_7842, mcs1_mcs_mat1_4_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({new_AGEMA_signal_9205, new_AGEMA_signal_9204, mcs1_mcs_mat1_4_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_10001, new_AGEMA_signal_10000, mcs1_mcs_mat1_4_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_7845, new_AGEMA_signal_7844, mcs1_mcs_mat1_4_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_9205, new_AGEMA_signal_9204, mcs1_mcs_mat1_4_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .b ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .c ({new_AGEMA_signal_10003, new_AGEMA_signal_10002, mcs1_mcs_mat1_4_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023]}), .c ({new_AGEMA_signal_7845, new_AGEMA_signal_7844, mcs1_mcs_mat1_4_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_7847, new_AGEMA_signal_7846, mcs1_mcs_mat1_4_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_9209, new_AGEMA_signal_9208, mcs1_mcs_mat1_4_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_7847, new_AGEMA_signal_7846, mcs1_mcs_mat1_4_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .c ({new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_4_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_7847, new_AGEMA_signal_7846, mcs1_mcs_mat1_4_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_13289, new_AGEMA_signal_13288, mcs1_mcs_mat1_4_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .c ({new_AGEMA_signal_13745, new_AGEMA_signal_13744, mcs1_mcs_mat1_4_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_10971, new_AGEMA_signal_10970, mcs1_mcs_mat1_4_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_13289, new_AGEMA_signal_13288, mcs1_mcs_mat1_4_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_13291, new_AGEMA_signal_13290, mcs1_mcs_mat1_4_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029]}), .c ({new_AGEMA_signal_10971, new_AGEMA_signal_10970, mcs1_mcs_mat1_4_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .b ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .c ({new_AGEMA_signal_9213, new_AGEMA_signal_9212, mcs1_mcs_mat1_4_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .b ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_9215, new_AGEMA_signal_9214, mcs1_mcs_mat1_4_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, mcs1_mcs_mat1_4_mcs_out[87]}), .c ({new_AGEMA_signal_10973, new_AGEMA_signal_10972, mcs1_mcs_mat1_4_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .c ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, mcs1_mcs_mat1_4_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .c ({new_AGEMA_signal_10017, new_AGEMA_signal_10016, mcs1_mcs_mat1_4_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_7849, new_AGEMA_signal_7848, mcs1_mcs_mat1_4_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_10983, new_AGEMA_signal_10982, mcs1_mcs_mat1_4_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_11949, new_AGEMA_signal_11948, mcs1_mcs_mat1_4_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035]}), .c ({new_AGEMA_signal_10983, new_AGEMA_signal_10982, mcs1_mcs_mat1_4_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_7851, new_AGEMA_signal_7850, mcs1_mcs_mat1_4_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_4_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_7851, new_AGEMA_signal_7850, mcs1_mcs_mat1_4_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041]}), .c ({new_AGEMA_signal_7853, new_AGEMA_signal_7852, mcs1_mcs_mat1_4_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_7855, new_AGEMA_signal_7854, mcs1_mcs_mat1_4_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .c ({new_AGEMA_signal_10033, new_AGEMA_signal_10032, mcs1_mcs_mat1_4_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_7855, new_AGEMA_signal_7854, mcs1_mcs_mat1_4_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_14635, new_AGEMA_signal_14634, mcs1_mcs_mat1_4_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_10995, new_AGEMA_signal_10994, mcs1_mcs_mat1_4_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_15115, new_AGEMA_signal_15114, mcs1_mcs_mat1_4_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_14203, new_AGEMA_signal_14202, mcs1_mcs_mat1_4_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_14635, new_AGEMA_signal_14634, mcs1_mcs_mat1_4_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_13755, new_AGEMA_signal_13754, mcs1_mcs_mat1_4_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_14203, new_AGEMA_signal_14202, mcs1_mcs_mat1_4_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_13755, new_AGEMA_signal_13754, mcs1_mcs_mat1_4_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047]}), .c ({new_AGEMA_signal_10995, new_AGEMA_signal_10994, mcs1_mcs_mat1_4_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_10039, new_AGEMA_signal_10038, mcs1_mcs_mat1_4_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_8423, new_AGEMA_signal_8422, mcs1_mcs_mat1_4_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_10997, new_AGEMA_signal_10996, mcs1_mcs_mat1_4_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_7857, new_AGEMA_signal_7856, mcs1_mcs_mat1_4_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .c ({new_AGEMA_signal_8423, new_AGEMA_signal_8422, mcs1_mcs_mat1_4_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .c ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, mcs1_mcs_mat1_4_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .c ({new_AGEMA_signal_10039, new_AGEMA_signal_10038, mcs1_mcs_mat1_4_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_7857, new_AGEMA_signal_7856, mcs1_mcs_mat1_4_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_10041, new_AGEMA_signal_10040, mcs1_mcs_mat1_4_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_7857, new_AGEMA_signal_7856, mcs1_mcs_mat1_4_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .b ({new_AGEMA_signal_7859, new_AGEMA_signal_7858, mcs1_mcs_mat1_4_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_10049, new_AGEMA_signal_10048, mcs1_mcs_mat1_4_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053]}), .c ({new_AGEMA_signal_7859, new_AGEMA_signal_7858, mcs1_mcs_mat1_4_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({new_AGEMA_signal_10053, new_AGEMA_signal_10052, mcs1_mcs_mat1_4_mcs_out[51]}), .c ({new_AGEMA_signal_11007, new_AGEMA_signal_11006, mcs1_mcs_mat1_4_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .c ({new_AGEMA_signal_10053, new_AGEMA_signal_10052, mcs1_mcs_mat1_4_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_11009, new_AGEMA_signal_11008, mcs1_mcs_mat1_4_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_13301, new_AGEMA_signal_13300, mcs1_mcs_mat1_4_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_11009, new_AGEMA_signal_11008, mcs1_mcs_mat1_4_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_10055, new_AGEMA_signal_10054, mcs1_mcs_mat1_4_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_11013, new_AGEMA_signal_11012, mcs1_mcs_mat1_4_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .b ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_10055, new_AGEMA_signal_10054, mcs1_mcs_mat1_4_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_9231, new_AGEMA_signal_9230, mcs1_mcs_mat1_4_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_10057, new_AGEMA_signal_10056, mcs1_mcs_mat1_4_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .c ({new_AGEMA_signal_9231, new_AGEMA_signal_9230, mcs1_mcs_mat1_4_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059]}), .c ({new_AGEMA_signal_7861, new_AGEMA_signal_7860, mcs1_mcs_mat1_4_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({new_AGEMA_signal_7863, new_AGEMA_signal_7862, mcs1_mcs_mat1_4_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9235, new_AGEMA_signal_9234, mcs1_mcs_mat1_4_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .b ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_10063, new_AGEMA_signal_10062, mcs1_mcs_mat1_4_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_7863, new_AGEMA_signal_7862, mcs1_mcs_mat1_4_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_11987, new_AGEMA_signal_11986, mcs1_mcs_mat1_4_mcs_out[35]}), .b ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_12733, new_AGEMA_signal_12732, mcs1_mcs_mat1_4_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_11025, new_AGEMA_signal_11024, mcs1_mcs_mat1_4_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_7865, new_AGEMA_signal_7864, mcs1_mcs_mat1_4_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_11987, new_AGEMA_signal_11986, mcs1_mcs_mat1_4_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_10067, new_AGEMA_signal_10066, mcs1_mcs_mat1_4_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .c ({new_AGEMA_signal_11025, new_AGEMA_signal_11024, mcs1_mcs_mat1_4_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .c ({new_AGEMA_signal_10067, new_AGEMA_signal_10066, mcs1_mcs_mat1_4_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065]}), .c ({new_AGEMA_signal_7865, new_AGEMA_signal_7864, mcs1_mcs_mat1_4_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_11027, new_AGEMA_signal_11026, mcs1_mcs_mat1_4_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_11989, new_AGEMA_signal_11988, mcs1_mcs_mat1_4_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({new_AGEMA_signal_13763, new_AGEMA_signal_13762, mcs1_mcs_mat1_4_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_14209, new_AGEMA_signal_14208, mcs1_mcs_mat1_4_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_11027, new_AGEMA_signal_11026, mcs1_mcs_mat1_4_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_13763, new_AGEMA_signal_13762, mcs1_mcs_mat1_4_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_11027, new_AGEMA_signal_11026, mcs1_mcs_mat1_4_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071]}), .c ({new_AGEMA_signal_7867, new_AGEMA_signal_7866, mcs1_mcs_mat1_4_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_7869, new_AGEMA_signal_7868, mcs1_mcs_mat1_4_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_9247, new_AGEMA_signal_9246, mcs1_mcs_mat1_4_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_10083, new_AGEMA_signal_10082, mcs1_mcs_mat1_4_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_9247, new_AGEMA_signal_9246, mcs1_mcs_mat1_4_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .c ({new_AGEMA_signal_10087, new_AGEMA_signal_10086, mcs1_mcs_mat1_4_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077]}), .c ({new_AGEMA_signal_7871, new_AGEMA_signal_7870, mcs1_mcs_mat1_4_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_11047, new_AGEMA_signal_11046, mcs1_mcs_mat1_4_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083]}), .c ({new_AGEMA_signal_7873, new_AGEMA_signal_7872, mcs1_mcs_mat1_4_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_7875, new_AGEMA_signal_7874, mcs1_mcs_mat1_4_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_9255, new_AGEMA_signal_9254, mcs1_mcs_mat1_4_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_7875, new_AGEMA_signal_7874, mcs1_mcs_mat1_4_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_8445, new_AGEMA_signal_8444, mcs1_mcs_mat1_4_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_7875, new_AGEMA_signal_7874, mcs1_mcs_mat1_4_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_10099, new_AGEMA_signal_10098, mcs1_mcs_mat1_4_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7877, new_AGEMA_signal_7876, mcs1_mcs_mat1_4_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_11055, new_AGEMA_signal_11054, mcs1_mcs_mat1_4_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_10099, new_AGEMA_signal_10098, mcs1_mcs_mat1_4_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .c ({new_AGEMA_signal_11059, new_AGEMA_signal_11058, mcs1_mcs_mat1_4_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_9259, new_AGEMA_signal_9258, mcs1_mcs_mat1_4_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_10099, new_AGEMA_signal_10098, mcs1_mcs_mat1_4_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_9259, new_AGEMA_signal_9258, mcs1_mcs_mat1_4_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .c ({new_AGEMA_signal_10101, new_AGEMA_signal_10100, mcs1_mcs_mat1_4_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089]}), .c ({new_AGEMA_signal_7877, new_AGEMA_signal_7876, mcs1_mcs_mat1_4_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U44 ( .a ({new_AGEMA_signal_9291, new_AGEMA_signal_9290, mcs1_mcs_mat1_5_mcs_out[90]}), .b ({new_AGEMA_signal_10131, new_AGEMA_signal_10130, mcs1_mcs_mat1_5_mcs_out[94]}), .c ({new_AGEMA_signal_11065, new_AGEMA_signal_11064, mcs1_mcs_mat1_5_n93}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .c ({new_AGEMA_signal_9263, new_AGEMA_signal_9262, mcs1_mcs_mat1_5_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .b ({new_AGEMA_signal_7879, new_AGEMA_signal_7878, mcs1_mcs_mat1_5_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8451, new_AGEMA_signal_8450, mcs1_mcs_mat1_5_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_7879, new_AGEMA_signal_7878, mcs1_mcs_mat1_5_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_9269, new_AGEMA_signal_9268, mcs1_mcs_mat1_5_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_10109, new_AGEMA_signal_10108, mcs1_mcs_mat1_5_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_7881, new_AGEMA_signal_7880, mcs1_mcs_mat1_5_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_9269, new_AGEMA_signal_9268, mcs1_mcs_mat1_5_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095]}), .c ({new_AGEMA_signal_7881, new_AGEMA_signal_7880, mcs1_mcs_mat1_5_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_11077, new_AGEMA_signal_11076, mcs1_mcs_mat1_5_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_13787, new_AGEMA_signal_13786, mcs1_mcs_mat1_5_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_14229, new_AGEMA_signal_14228, mcs1_mcs_mat1_5_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_12037, new_AGEMA_signal_12036, mcs1_mcs_mat1_5_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, mcs1_mcs_mat1_5_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .c ({new_AGEMA_signal_12037, new_AGEMA_signal_12036, mcs1_mcs_mat1_5_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .b ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_13787, new_AGEMA_signal_13786, mcs1_mcs_mat1_5_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_11077, new_AGEMA_signal_11076, mcs1_mcs_mat1_5_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_10115, new_AGEMA_signal_10114, mcs1_mcs_mat1_5_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_11079, new_AGEMA_signal_11078, mcs1_mcs_mat1_5_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_7883, new_AGEMA_signal_7882, mcs1_mcs_mat1_5_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_10115, new_AGEMA_signal_10114, mcs1_mcs_mat1_5_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101]}), .c ({new_AGEMA_signal_7883, new_AGEMA_signal_7882, mcs1_mcs_mat1_5_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_7885, new_AGEMA_signal_7884, mcs1_mcs_mat1_5_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({new_AGEMA_signal_9281, new_AGEMA_signal_9280, mcs1_mcs_mat1_5_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_10123, new_AGEMA_signal_10122, mcs1_mcs_mat1_5_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_7887, new_AGEMA_signal_7886, mcs1_mcs_mat1_5_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_9281, new_AGEMA_signal_9280, mcs1_mcs_mat1_5_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .b ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .c ({new_AGEMA_signal_10125, new_AGEMA_signal_10124, mcs1_mcs_mat1_5_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107]}), .c ({new_AGEMA_signal_7887, new_AGEMA_signal_7886, mcs1_mcs_mat1_5_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_11093, new_AGEMA_signal_11092, mcs1_mcs_mat1_5_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_13345, new_AGEMA_signal_13344, mcs1_mcs_mat1_5_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_11093, new_AGEMA_signal_11092, mcs1_mcs_mat1_5_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .c ({new_AGEMA_signal_12057, new_AGEMA_signal_12056, mcs1_mcs_mat1_5_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_11093, new_AGEMA_signal_11092, mcs1_mcs_mat1_5_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_9285, new_AGEMA_signal_9284, mcs1_mcs_mat1_5_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .c ({new_AGEMA_signal_10131, new_AGEMA_signal_10130, mcs1_mcs_mat1_5_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_7889, new_AGEMA_signal_7888, mcs1_mcs_mat1_5_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_9285, new_AGEMA_signal_9284, mcs1_mcs_mat1_5_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_9287, new_AGEMA_signal_9286, mcs1_mcs_mat1_5_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113]}), .c ({new_AGEMA_signal_7889, new_AGEMA_signal_7888, mcs1_mcs_mat1_5_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .b ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .c ({new_AGEMA_signal_9291, new_AGEMA_signal_9290, mcs1_mcs_mat1_5_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .b ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_9293, new_AGEMA_signal_9292, mcs1_mcs_mat1_5_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({new_AGEMA_signal_10137, new_AGEMA_signal_10136, mcs1_mcs_mat1_5_mcs_out[87]}), .c ({new_AGEMA_signal_11097, new_AGEMA_signal_11096, mcs1_mcs_mat1_5_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .c ({new_AGEMA_signal_10137, new_AGEMA_signal_10136, mcs1_mcs_mat1_5_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .c ({new_AGEMA_signal_13797, new_AGEMA_signal_13796, mcs1_mcs_mat1_5_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_11099, new_AGEMA_signal_11098, mcs1_mcs_mat1_5_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_7891, new_AGEMA_signal_7890, mcs1_mcs_mat1_5_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_8465, new_AGEMA_signal_8464, mcs1_mcs_mat1_5_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119]}), .c ({new_AGEMA_signal_7891, new_AGEMA_signal_7890, mcs1_mcs_mat1_5_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_7893, new_AGEMA_signal_7892, mcs1_mcs_mat1_5_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, mcs1_mcs_mat1_5_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_7893, new_AGEMA_signal_7892, mcs1_mcs_mat1_5_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125]}), .c ({new_AGEMA_signal_7895, new_AGEMA_signal_7894, mcs1_mcs_mat1_5_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_11111, new_AGEMA_signal_11110, mcs1_mcs_mat1_5_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .c ({new_AGEMA_signal_13801, new_AGEMA_signal_13800, mcs1_mcs_mat1_5_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_11111, new_AGEMA_signal_11110, mcs1_mcs_mat1_5_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_12085, new_AGEMA_signal_12084, mcs1_mcs_mat1_5_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_7897, new_AGEMA_signal_7896, mcs1_mcs_mat1_5_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_12801, new_AGEMA_signal_12800, mcs1_mcs_mat1_5_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_11117, new_AGEMA_signal_11116, mcs1_mcs_mat1_5_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_12085, new_AGEMA_signal_12084, mcs1_mcs_mat1_5_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, mcs1_mcs_mat1_5_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_11117, new_AGEMA_signal_11116, mcs1_mcs_mat1_5_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, mcs1_mcs_mat1_5_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131]}), .c ({new_AGEMA_signal_7897, new_AGEMA_signal_7896, mcs1_mcs_mat1_5_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_10161, new_AGEMA_signal_10160, mcs1_mcs_mat1_5_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_8477, new_AGEMA_signal_8476, mcs1_mcs_mat1_5_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_11119, new_AGEMA_signal_11118, mcs1_mcs_mat1_5_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_7899, new_AGEMA_signal_7898, mcs1_mcs_mat1_5_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .c ({new_AGEMA_signal_8477, new_AGEMA_signal_8476, mcs1_mcs_mat1_5_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .c ({new_AGEMA_signal_8479, new_AGEMA_signal_8478, mcs1_mcs_mat1_5_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .c ({new_AGEMA_signal_10161, new_AGEMA_signal_10160, mcs1_mcs_mat1_5_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_7899, new_AGEMA_signal_7898, mcs1_mcs_mat1_5_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_10163, new_AGEMA_signal_10162, mcs1_mcs_mat1_5_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_7899, new_AGEMA_signal_7898, mcs1_mcs_mat1_5_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .b ({new_AGEMA_signal_7901, new_AGEMA_signal_7900, mcs1_mcs_mat1_5_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_10171, new_AGEMA_signal_10170, mcs1_mcs_mat1_5_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137]}), .c ({new_AGEMA_signal_7901, new_AGEMA_signal_7900, mcs1_mcs_mat1_5_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({new_AGEMA_signal_13805, new_AGEMA_signal_13804, mcs1_mcs_mat1_5_mcs_out[51]}), .c ({new_AGEMA_signal_14247, new_AGEMA_signal_14246, mcs1_mcs_mat1_5_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .c ({new_AGEMA_signal_13805, new_AGEMA_signal_13804, mcs1_mcs_mat1_5_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_7903, new_AGEMA_signal_7902, mcs1_mcs_mat1_5_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_9309, new_AGEMA_signal_9308, mcs1_mcs_mat1_5_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_7903, new_AGEMA_signal_7902, mcs1_mcs_mat1_5_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_10179, new_AGEMA_signal_10178, mcs1_mcs_mat1_5_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_11133, new_AGEMA_signal_11132, mcs1_mcs_mat1_5_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .b ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_10179, new_AGEMA_signal_10178, mcs1_mcs_mat1_5_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_9313, new_AGEMA_signal_9312, mcs1_mcs_mat1_5_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_10181, new_AGEMA_signal_10180, mcs1_mcs_mat1_5_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .c ({new_AGEMA_signal_9313, new_AGEMA_signal_9312, mcs1_mcs_mat1_5_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143]}), .c ({new_AGEMA_signal_7905, new_AGEMA_signal_7904, mcs1_mcs_mat1_5_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({new_AGEMA_signal_7907, new_AGEMA_signal_7906, mcs1_mcs_mat1_5_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9317, new_AGEMA_signal_9316, mcs1_mcs_mat1_5_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_10187, new_AGEMA_signal_10186, mcs1_mcs_mat1_5_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_7907, new_AGEMA_signal_7906, mcs1_mcs_mat1_5_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_14691, new_AGEMA_signal_14690, mcs1_mcs_mat1_5_mcs_out[35]}), .b ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_15171, new_AGEMA_signal_15170, mcs1_mcs_mat1_5_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_14251, new_AGEMA_signal_14250, mcs1_mcs_mat1_5_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_11143, new_AGEMA_signal_11142, mcs1_mcs_mat1_5_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_14691, new_AGEMA_signal_14690, mcs1_mcs_mat1_5_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_13807, new_AGEMA_signal_13806, mcs1_mcs_mat1_5_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .c ({new_AGEMA_signal_14251, new_AGEMA_signal_14250, mcs1_mcs_mat1_5_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .c ({new_AGEMA_signal_13807, new_AGEMA_signal_13806, mcs1_mcs_mat1_5_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149]}), .c ({new_AGEMA_signal_11143, new_AGEMA_signal_11142, mcs1_mcs_mat1_5_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_7909, new_AGEMA_signal_7908, mcs1_mcs_mat1_5_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_8491, new_AGEMA_signal_8490, mcs1_mcs_mat1_5_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, mcs1_mcs_mat1_5_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_11147, new_AGEMA_signal_11146, mcs1_mcs_mat1_5_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_7909, new_AGEMA_signal_7908, mcs1_mcs_mat1_5_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, mcs1_mcs_mat1_5_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_7909, new_AGEMA_signal_7908, mcs1_mcs_mat1_5_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155]}), .c ({new_AGEMA_signal_7911, new_AGEMA_signal_7910, mcs1_mcs_mat1_5_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_7913, new_AGEMA_signal_7912, mcs1_mcs_mat1_5_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_13357, new_AGEMA_signal_13356, mcs1_mcs_mat1_5_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_13811, new_AGEMA_signal_13810, mcs1_mcs_mat1_5_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_13357, new_AGEMA_signal_13356, mcs1_mcs_mat1_5_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .c ({new_AGEMA_signal_13815, new_AGEMA_signal_13814, mcs1_mcs_mat1_5_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161]}), .c ({new_AGEMA_signal_11163, new_AGEMA_signal_11162, mcs1_mcs_mat1_5_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_7915, new_AGEMA_signal_7914, mcs1_mcs_mat1_5_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167]}), .c ({new_AGEMA_signal_7917, new_AGEMA_signal_7916, mcs1_mcs_mat1_5_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_7919, new_AGEMA_signal_7918, mcs1_mcs_mat1_5_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_9335, new_AGEMA_signal_9334, mcs1_mcs_mat1_5_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_7919, new_AGEMA_signal_7918, mcs1_mcs_mat1_5_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_8503, new_AGEMA_signal_8502, mcs1_mcs_mat1_5_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_7919, new_AGEMA_signal_7918, mcs1_mcs_mat1_5_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_13823, new_AGEMA_signal_13822, mcs1_mcs_mat1_5_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_11177, new_AGEMA_signal_11176, mcs1_mcs_mat1_5_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_14259, new_AGEMA_signal_14258, mcs1_mcs_mat1_5_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_13823, new_AGEMA_signal_13822, mcs1_mcs_mat1_5_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .c ({new_AGEMA_signal_14263, new_AGEMA_signal_14262, mcs1_mcs_mat1_5_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, mcs1_mcs_mat1_5_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_13823, new_AGEMA_signal_13822, mcs1_mcs_mat1_5_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, mcs1_mcs_mat1_5_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .c ({new_AGEMA_signal_13825, new_AGEMA_signal_13824, mcs1_mcs_mat1_5_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173]}), .c ({new_AGEMA_signal_11177, new_AGEMA_signal_11176, mcs1_mcs_mat1_5_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U44 ( .a ({new_AGEMA_signal_9365, new_AGEMA_signal_9364, mcs1_mcs_mat1_6_mcs_out[90]}), .b ({new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_6_mcs_out[94]}), .c ({new_AGEMA_signal_11181, new_AGEMA_signal_11180, mcs1_mcs_mat1_6_n93}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .c ({new_AGEMA_signal_9339, new_AGEMA_signal_9338, mcs1_mcs_mat1_6_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .b ({new_AGEMA_signal_7921, new_AGEMA_signal_7920, mcs1_mcs_mat1_6_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_8507, new_AGEMA_signal_8506, mcs1_mcs_mat1_6_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_7921, new_AGEMA_signal_7920, mcs1_mcs_mat1_6_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_13397, new_AGEMA_signal_13396, mcs1_mcs_mat1_6_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_13837, new_AGEMA_signal_13836, mcs1_mcs_mat1_6_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_11189, new_AGEMA_signal_11188, mcs1_mcs_mat1_6_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_13397, new_AGEMA_signal_13396, mcs1_mcs_mat1_6_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179]}), .c ({new_AGEMA_signal_11189, new_AGEMA_signal_11188, mcs1_mcs_mat1_6_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_7923, new_AGEMA_signal_7922, mcs1_mcs_mat1_6_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, mcs1_mcs_mat1_6_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_11191, new_AGEMA_signal_11190, mcs1_mcs_mat1_6_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_8511, new_AGEMA_signal_8510, mcs1_mcs_mat1_6_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_9345, new_AGEMA_signal_9344, mcs1_mcs_mat1_6_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .c ({new_AGEMA_signal_8511, new_AGEMA_signal_8510, mcs1_mcs_mat1_6_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, mcs1_mcs_mat1_6_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_7923, new_AGEMA_signal_7922, mcs1_mcs_mat1_6_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_10229, new_AGEMA_signal_10228, mcs1_mcs_mat1_6_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_11197, new_AGEMA_signal_11196, mcs1_mcs_mat1_6_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_7925, new_AGEMA_signal_7924, mcs1_mcs_mat1_6_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_10229, new_AGEMA_signal_10228, mcs1_mcs_mat1_6_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185]}), .c ({new_AGEMA_signal_7925, new_AGEMA_signal_7924, mcs1_mcs_mat1_6_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_7927, new_AGEMA_signal_7926, mcs1_mcs_mat1_6_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({new_AGEMA_signal_13403, new_AGEMA_signal_13402, mcs1_mcs_mat1_6_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_13843, new_AGEMA_signal_13842, mcs1_mcs_mat1_6_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_11205, new_AGEMA_signal_11204, mcs1_mcs_mat1_6_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_13403, new_AGEMA_signal_13402, mcs1_mcs_mat1_6_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .c ({new_AGEMA_signal_13845, new_AGEMA_signal_13844, mcs1_mcs_mat1_6_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191]}), .c ({new_AGEMA_signal_11205, new_AGEMA_signal_11204, mcs1_mcs_mat1_6_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_7929, new_AGEMA_signal_7928, mcs1_mcs_mat1_6_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_9355, new_AGEMA_signal_9354, mcs1_mcs_mat1_6_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_7929, new_AGEMA_signal_7928, mcs1_mcs_mat1_6_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .c ({new_AGEMA_signal_8519, new_AGEMA_signal_8518, mcs1_mcs_mat1_6_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_7929, new_AGEMA_signal_7928, mcs1_mcs_mat1_6_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_9359, new_AGEMA_signal_9358, mcs1_mcs_mat1_6_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .c ({new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_6_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_7931, new_AGEMA_signal_7930, mcs1_mcs_mat1_6_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_9359, new_AGEMA_signal_9358, mcs1_mcs_mat1_6_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_9361, new_AGEMA_signal_9360, mcs1_mcs_mat1_6_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197]}), .c ({new_AGEMA_signal_7931, new_AGEMA_signal_7930, mcs1_mcs_mat1_6_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .b ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .c ({new_AGEMA_signal_9365, new_AGEMA_signal_9364, mcs1_mcs_mat1_6_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .b ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_9367, new_AGEMA_signal_9366, mcs1_mcs_mat1_6_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({new_AGEMA_signal_13853, new_AGEMA_signal_13852, mcs1_mcs_mat1_6_mcs_out[87]}), .c ({new_AGEMA_signal_14287, new_AGEMA_signal_14286, mcs1_mcs_mat1_6_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .c ({new_AGEMA_signal_13853, new_AGEMA_signal_13852, mcs1_mcs_mat1_6_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .c ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, mcs1_mcs_mat1_6_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_7933, new_AGEMA_signal_7932, mcs1_mcs_mat1_6_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, mcs1_mcs_mat1_6_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_8527, new_AGEMA_signal_8526, mcs1_mcs_mat1_6_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203]}), .c ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, mcs1_mcs_mat1_6_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_7937, new_AGEMA_signal_7936, mcs1_mcs_mat1_6_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_8531, new_AGEMA_signal_8530, mcs1_mcs_mat1_6_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_7937, new_AGEMA_signal_7936, mcs1_mcs_mat1_6_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209]}), .c ({new_AGEMA_signal_11225, new_AGEMA_signal_11224, mcs1_mcs_mat1_6_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_7939, new_AGEMA_signal_7938, mcs1_mcs_mat1_6_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .c ({new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_6_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_7939, new_AGEMA_signal_7938, mcs1_mcs_mat1_6_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_12195, new_AGEMA_signal_12194, mcs1_mcs_mat1_6_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_7941, new_AGEMA_signal_7940, mcs1_mcs_mat1_6_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_12883, new_AGEMA_signal_12882, mcs1_mcs_mat1_6_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_11233, new_AGEMA_signal_11232, mcs1_mcs_mat1_6_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_12195, new_AGEMA_signal_12194, mcs1_mcs_mat1_6_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, mcs1_mcs_mat1_6_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_11233, new_AGEMA_signal_11232, mcs1_mcs_mat1_6_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, mcs1_mcs_mat1_6_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215]}), .c ({new_AGEMA_signal_7941, new_AGEMA_signal_7940, mcs1_mcs_mat1_6_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, mcs1_mcs_mat1_6_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_8539, new_AGEMA_signal_8538, mcs1_mcs_mat1_6_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_11235, new_AGEMA_signal_11234, mcs1_mcs_mat1_6_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_7943, new_AGEMA_signal_7942, mcs1_mcs_mat1_6_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .c ({new_AGEMA_signal_8539, new_AGEMA_signal_8538, mcs1_mcs_mat1_6_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .c ({new_AGEMA_signal_8541, new_AGEMA_signal_8540, mcs1_mcs_mat1_6_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .c ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, mcs1_mcs_mat1_6_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_7943, new_AGEMA_signal_7942, mcs1_mcs_mat1_6_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_10275, new_AGEMA_signal_10274, mcs1_mcs_mat1_6_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_7943, new_AGEMA_signal_7942, mcs1_mcs_mat1_6_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .b ({new_AGEMA_signal_11241, new_AGEMA_signal_11240, mcs1_mcs_mat1_6_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_13865, new_AGEMA_signal_13864, mcs1_mcs_mat1_6_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221]}), .c ({new_AGEMA_signal_11241, new_AGEMA_signal_11240, mcs1_mcs_mat1_6_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({new_AGEMA_signal_10279, new_AGEMA_signal_10278, mcs1_mcs_mat1_6_mcs_out[51]}), .c ({new_AGEMA_signal_11243, new_AGEMA_signal_11242, mcs1_mcs_mat1_6_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .c ({new_AGEMA_signal_10279, new_AGEMA_signal_10278, mcs1_mcs_mat1_6_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_7945, new_AGEMA_signal_7944, mcs1_mcs_mat1_6_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_9381, new_AGEMA_signal_9380, mcs1_mcs_mat1_6_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_7945, new_AGEMA_signal_7944, mcs1_mcs_mat1_6_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_10285, new_AGEMA_signal_10284, mcs1_mcs_mat1_6_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_11249, new_AGEMA_signal_11248, mcs1_mcs_mat1_6_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .b ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_10285, new_AGEMA_signal_10284, mcs1_mcs_mat1_6_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_9385, new_AGEMA_signal_9384, mcs1_mcs_mat1_6_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_10287, new_AGEMA_signal_10286, mcs1_mcs_mat1_6_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .c ({new_AGEMA_signal_9385, new_AGEMA_signal_9384, mcs1_mcs_mat1_6_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227]}), .c ({new_AGEMA_signal_7947, new_AGEMA_signal_7946, mcs1_mcs_mat1_6_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({new_AGEMA_signal_11255, new_AGEMA_signal_11254, mcs1_mcs_mat1_6_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_13419, new_AGEMA_signal_13418, mcs1_mcs_mat1_6_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .b ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_13871, new_AGEMA_signal_13870, mcs1_mcs_mat1_6_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_11255, new_AGEMA_signal_11254, mcs1_mcs_mat1_6_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_12211, new_AGEMA_signal_12210, mcs1_mcs_mat1_6_mcs_out[35]}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_12889, new_AGEMA_signal_12888, mcs1_mcs_mat1_6_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_11259, new_AGEMA_signal_11258, mcs1_mcs_mat1_6_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_7949, new_AGEMA_signal_7948, mcs1_mcs_mat1_6_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_12211, new_AGEMA_signal_12210, mcs1_mcs_mat1_6_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_10291, new_AGEMA_signal_10290, mcs1_mcs_mat1_6_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .c ({new_AGEMA_signal_11259, new_AGEMA_signal_11258, mcs1_mcs_mat1_6_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .c ({new_AGEMA_signal_10291, new_AGEMA_signal_10290, mcs1_mcs_mat1_6_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233]}), .c ({new_AGEMA_signal_7949, new_AGEMA_signal_7948, mcs1_mcs_mat1_6_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_7951, new_AGEMA_signal_7950, mcs1_mcs_mat1_6_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_8551, new_AGEMA_signal_8550, mcs1_mcs_mat1_6_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({new_AGEMA_signal_10295, new_AGEMA_signal_10294, mcs1_mcs_mat1_6_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_11263, new_AGEMA_signal_11262, mcs1_mcs_mat1_6_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_7951, new_AGEMA_signal_7950, mcs1_mcs_mat1_6_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_10295, new_AGEMA_signal_10294, mcs1_mcs_mat1_6_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_7951, new_AGEMA_signal_7950, mcs1_mcs_mat1_6_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239]}), .c ({new_AGEMA_signal_7953, new_AGEMA_signal_7952, mcs1_mcs_mat1_6_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_11273, new_AGEMA_signal_11272, mcs1_mcs_mat1_6_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_9395, new_AGEMA_signal_9394, mcs1_mcs_mat1_6_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_10307, new_AGEMA_signal_10306, mcs1_mcs_mat1_6_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_9395, new_AGEMA_signal_9394, mcs1_mcs_mat1_6_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .c ({new_AGEMA_signal_10311, new_AGEMA_signal_10310, mcs1_mcs_mat1_6_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245]}), .c ({new_AGEMA_signal_7955, new_AGEMA_signal_7954, mcs1_mcs_mat1_6_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_7957, new_AGEMA_signal_7956, mcs1_mcs_mat1_6_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251]}), .c ({new_AGEMA_signal_7959, new_AGEMA_signal_7958, mcs1_mcs_mat1_6_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_11291, new_AGEMA_signal_11290, mcs1_mcs_mat1_6_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_13431, new_AGEMA_signal_13430, mcs1_mcs_mat1_6_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_11291, new_AGEMA_signal_11290, mcs1_mcs_mat1_6_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_12239, new_AGEMA_signal_12238, mcs1_mcs_mat1_6_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_11291, new_AGEMA_signal_11290, mcs1_mcs_mat1_6_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_10325, new_AGEMA_signal_10324, mcs1_mcs_mat1_6_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_7961, new_AGEMA_signal_7960, mcs1_mcs_mat1_6_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_11293, new_AGEMA_signal_11292, mcs1_mcs_mat1_6_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_10325, new_AGEMA_signal_10324, mcs1_mcs_mat1_6_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .c ({new_AGEMA_signal_11297, new_AGEMA_signal_11296, mcs1_mcs_mat1_6_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_9405, new_AGEMA_signal_9404, mcs1_mcs_mat1_6_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_10325, new_AGEMA_signal_10324, mcs1_mcs_mat1_6_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_9405, new_AGEMA_signal_9404, mcs1_mcs_mat1_6_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .c ({new_AGEMA_signal_10327, new_AGEMA_signal_10326, mcs1_mcs_mat1_6_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257]}), .c ({new_AGEMA_signal_7961, new_AGEMA_signal_7960, mcs1_mcs_mat1_6_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U44 ( .a ({new_AGEMA_signal_13477, new_AGEMA_signal_13476, mcs1_mcs_mat1_7_mcs_out[90]}), .b ({new_AGEMA_signal_10357, new_AGEMA_signal_10356, mcs1_mcs_mat1_7_mcs_out[94]}), .c ({new_AGEMA_signal_13889, new_AGEMA_signal_13888, mcs1_mcs_mat1_7_n93}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .c ({new_AGEMA_signal_9409, new_AGEMA_signal_9408, mcs1_mcs_mat1_7_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .b ({new_AGEMA_signal_11301, new_AGEMA_signal_11300, mcs1_mcs_mat1_7_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_12261, new_AGEMA_signal_12260, mcs1_mcs_mat1_7_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_11301, new_AGEMA_signal_11300, mcs1_mcs_mat1_7_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_9411, new_AGEMA_signal_9410, mcs1_mcs_mat1_7_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_10331, new_AGEMA_signal_10330, mcs1_mcs_mat1_7_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_7963, new_AGEMA_signal_7962, mcs1_mcs_mat1_7_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_9411, new_AGEMA_signal_9410, mcs1_mcs_mat1_7_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263]}), .c ({new_AGEMA_signal_7963, new_AGEMA_signal_7962, mcs1_mcs_mat1_7_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_7965, new_AGEMA_signal_7964, mcs1_mcs_mat1_7_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_10339, new_AGEMA_signal_10338, mcs1_mcs_mat1_7_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_11307, new_AGEMA_signal_11306, mcs1_mcs_mat1_7_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_8567, new_AGEMA_signal_8566, mcs1_mcs_mat1_7_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_9417, new_AGEMA_signal_9416, mcs1_mcs_mat1_7_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .c ({new_AGEMA_signal_8567, new_AGEMA_signal_8566, mcs1_mcs_mat1_7_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .b ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_10339, new_AGEMA_signal_10338, mcs1_mcs_mat1_7_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_7965, new_AGEMA_signal_7964, mcs1_mcs_mat1_7_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_10343, new_AGEMA_signal_10342, mcs1_mcs_mat1_7_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_11313, new_AGEMA_signal_11312, mcs1_mcs_mat1_7_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_7967, new_AGEMA_signal_7966, mcs1_mcs_mat1_7_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_10343, new_AGEMA_signal_10342, mcs1_mcs_mat1_7_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269]}), .c ({new_AGEMA_signal_7967, new_AGEMA_signal_7966, mcs1_mcs_mat1_7_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_11317, new_AGEMA_signal_11316, mcs1_mcs_mat1_7_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({new_AGEMA_signal_9423, new_AGEMA_signal_9422, mcs1_mcs_mat1_7_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_10347, new_AGEMA_signal_10346, mcs1_mcs_mat1_7_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_7969, new_AGEMA_signal_7968, mcs1_mcs_mat1_7_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_9423, new_AGEMA_signal_9422, mcs1_mcs_mat1_7_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .b ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .c ({new_AGEMA_signal_10349, new_AGEMA_signal_10348, mcs1_mcs_mat1_7_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275]}), .c ({new_AGEMA_signal_7969, new_AGEMA_signal_7968, mcs1_mcs_mat1_7_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_7971, new_AGEMA_signal_7970, mcs1_mcs_mat1_7_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_9427, new_AGEMA_signal_9426, mcs1_mcs_mat1_7_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_7971, new_AGEMA_signal_7970, mcs1_mcs_mat1_7_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .c ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, mcs1_mcs_mat1_7_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_7971, new_AGEMA_signal_7970, mcs1_mcs_mat1_7_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_9431, new_AGEMA_signal_9430, mcs1_mcs_mat1_7_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .c ({new_AGEMA_signal_10357, new_AGEMA_signal_10356, mcs1_mcs_mat1_7_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_7973, new_AGEMA_signal_7972, mcs1_mcs_mat1_7_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_9431, new_AGEMA_signal_9430, mcs1_mcs_mat1_7_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_9433, new_AGEMA_signal_9432, mcs1_mcs_mat1_7_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281]}), .c ({new_AGEMA_signal_7973, new_AGEMA_signal_7972, mcs1_mcs_mat1_7_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .b ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .c ({new_AGEMA_signal_13477, new_AGEMA_signal_13476, mcs1_mcs_mat1_7_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .b ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_13479, new_AGEMA_signal_13478, mcs1_mcs_mat1_7_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({new_AGEMA_signal_10363, new_AGEMA_signal_10362, mcs1_mcs_mat1_7_mcs_out[87]}), .c ({new_AGEMA_signal_11329, new_AGEMA_signal_11328, mcs1_mcs_mat1_7_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .c ({new_AGEMA_signal_10363, new_AGEMA_signal_10362, mcs1_mcs_mat1_7_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .c ({new_AGEMA_signal_10369, new_AGEMA_signal_10368, mcs1_mcs_mat1_7_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_7975, new_AGEMA_signal_7974, mcs1_mcs_mat1_7_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_7977, new_AGEMA_signal_7976, mcs1_mcs_mat1_7_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_7_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287]}), .c ({new_AGEMA_signal_7977, new_AGEMA_signal_7976, mcs1_mcs_mat1_7_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_11341, new_AGEMA_signal_11340, mcs1_mcs_mat1_7_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_12297, new_AGEMA_signal_12296, mcs1_mcs_mat1_7_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_11341, new_AGEMA_signal_11340, mcs1_mcs_mat1_7_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293]}), .c ({new_AGEMA_signal_7979, new_AGEMA_signal_7978, mcs1_mcs_mat1_7_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_7981, new_AGEMA_signal_7980, mcs1_mcs_mat1_7_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .c ({new_AGEMA_signal_10383, new_AGEMA_signal_10382, mcs1_mcs_mat1_7_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_7981, new_AGEMA_signal_7980, mcs1_mcs_mat1_7_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_12313, new_AGEMA_signal_12312, mcs1_mcs_mat1_7_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_7983, new_AGEMA_signal_7982, mcs1_mcs_mat1_7_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_12947, new_AGEMA_signal_12946, mcs1_mcs_mat1_7_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_11353, new_AGEMA_signal_11352, mcs1_mcs_mat1_7_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_12313, new_AGEMA_signal_12312, mcs1_mcs_mat1_7_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_10387, new_AGEMA_signal_10386, mcs1_mcs_mat1_7_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_11353, new_AGEMA_signal_11352, mcs1_mcs_mat1_7_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_10387, new_AGEMA_signal_10386, mcs1_mcs_mat1_7_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299]}), .c ({new_AGEMA_signal_7983, new_AGEMA_signal_7982, mcs1_mcs_mat1_7_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_13917, new_AGEMA_signal_13916, mcs1_mcs_mat1_7_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_12315, new_AGEMA_signal_12314, mcs1_mcs_mat1_7_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_14337, new_AGEMA_signal_14336, mcs1_mcs_mat1_7_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_11355, new_AGEMA_signal_11354, mcs1_mcs_mat1_7_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .c ({new_AGEMA_signal_12315, new_AGEMA_signal_12314, mcs1_mcs_mat1_7_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .c ({new_AGEMA_signal_12317, new_AGEMA_signal_12316, mcs1_mcs_mat1_7_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .c ({new_AGEMA_signal_13917, new_AGEMA_signal_13916, mcs1_mcs_mat1_7_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_11355, new_AGEMA_signal_11354, mcs1_mcs_mat1_7_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_13919, new_AGEMA_signal_13918, mcs1_mcs_mat1_7_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_11355, new_AGEMA_signal_11354, mcs1_mcs_mat1_7_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .b ({new_AGEMA_signal_7985, new_AGEMA_signal_7984, mcs1_mcs_mat1_7_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_10395, new_AGEMA_signal_10394, mcs1_mcs_mat1_7_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305]}), .c ({new_AGEMA_signal_7985, new_AGEMA_signal_7984, mcs1_mcs_mat1_7_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({new_AGEMA_signal_10399, new_AGEMA_signal_10398, mcs1_mcs_mat1_7_mcs_out[51]}), .c ({new_AGEMA_signal_11361, new_AGEMA_signal_11360, mcs1_mcs_mat1_7_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .c ({new_AGEMA_signal_10399, new_AGEMA_signal_10398, mcs1_mcs_mat1_7_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_7987, new_AGEMA_signal_7986, mcs1_mcs_mat1_7_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_9451, new_AGEMA_signal_9450, mcs1_mcs_mat1_7_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_7987, new_AGEMA_signal_7986, mcs1_mcs_mat1_7_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_13923, new_AGEMA_signal_13922, mcs1_mcs_mat1_7_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_14345, new_AGEMA_signal_14344, mcs1_mcs_mat1_7_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .b ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_13923, new_AGEMA_signal_13922, mcs1_mcs_mat1_7_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_13489, new_AGEMA_signal_13488, mcs1_mcs_mat1_7_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_13925, new_AGEMA_signal_13924, mcs1_mcs_mat1_7_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .c ({new_AGEMA_signal_13489, new_AGEMA_signal_13488, mcs1_mcs_mat1_7_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311]}), .c ({new_AGEMA_signal_11365, new_AGEMA_signal_11364, mcs1_mcs_mat1_7_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({new_AGEMA_signal_7989, new_AGEMA_signal_7988, mcs1_mcs_mat1_7_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_9455, new_AGEMA_signal_9454, mcs1_mcs_mat1_7_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .b ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_7_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_7989, new_AGEMA_signal_7988, mcs1_mcs_mat1_7_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_12333, new_AGEMA_signal_12332, mcs1_mcs_mat1_7_mcs_out[35]}), .b ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_12959, new_AGEMA_signal_12958, mcs1_mcs_mat1_7_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_11373, new_AGEMA_signal_11372, mcs1_mcs_mat1_7_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_7991, new_AGEMA_signal_7990, mcs1_mcs_mat1_7_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_12333, new_AGEMA_signal_12332, mcs1_mcs_mat1_7_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, mcs1_mcs_mat1_7_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .c ({new_AGEMA_signal_11373, new_AGEMA_signal_11372, mcs1_mcs_mat1_7_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .c ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, mcs1_mcs_mat1_7_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317]}), .c ({new_AGEMA_signal_7991, new_AGEMA_signal_7990, mcs1_mcs_mat1_7_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_7993, new_AGEMA_signal_7992, mcs1_mcs_mat1_7_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_8601, new_AGEMA_signal_8600, mcs1_mcs_mat1_7_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({new_AGEMA_signal_10415, new_AGEMA_signal_10414, mcs1_mcs_mat1_7_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_11377, new_AGEMA_signal_11376, mcs1_mcs_mat1_7_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_7993, new_AGEMA_signal_7992, mcs1_mcs_mat1_7_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_10415, new_AGEMA_signal_10414, mcs1_mcs_mat1_7_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_7993, new_AGEMA_signal_7992, mcs1_mcs_mat1_7_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323]}), .c ({new_AGEMA_signal_11381, new_AGEMA_signal_11380, mcs1_mcs_mat1_7_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_7995, new_AGEMA_signal_7994, mcs1_mcs_mat1_7_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_9467, new_AGEMA_signal_9466, mcs1_mcs_mat1_7_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_10427, new_AGEMA_signal_10426, mcs1_mcs_mat1_7_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_9467, new_AGEMA_signal_9466, mcs1_mcs_mat1_7_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .c ({new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_7_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329]}), .c ({new_AGEMA_signal_7997, new_AGEMA_signal_7996, mcs1_mcs_mat1_7_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_7999, new_AGEMA_signal_7998, mcs1_mcs_mat1_7_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335]}), .c ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, mcs1_mcs_mat1_7_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_8001, new_AGEMA_signal_8000, mcs1_mcs_mat1_7_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_9473, new_AGEMA_signal_9472, mcs1_mcs_mat1_7_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_8001, new_AGEMA_signal_8000, mcs1_mcs_mat1_7_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, mcs1_mcs_mat1_7_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_8001, new_AGEMA_signal_8000, mcs1_mcs_mat1_7_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_10443, new_AGEMA_signal_10442, mcs1_mcs_mat1_7_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8003, new_AGEMA_signal_8002, mcs1_mcs_mat1_7_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_11405, new_AGEMA_signal_11404, mcs1_mcs_mat1_7_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_10443, new_AGEMA_signal_10442, mcs1_mcs_mat1_7_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .c ({new_AGEMA_signal_11409, new_AGEMA_signal_11408, mcs1_mcs_mat1_7_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_9477, new_AGEMA_signal_9476, mcs1_mcs_mat1_7_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_10443, new_AGEMA_signal_10442, mcs1_mcs_mat1_7_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_9477, new_AGEMA_signal_9476, mcs1_mcs_mat1_7_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .c ({new_AGEMA_signal_10445, new_AGEMA_signal_10444, mcs1_mcs_mat1_7_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341]}), .c ({new_AGEMA_signal_8003, new_AGEMA_signal_8002, mcs1_mcs_mat1_7_mcs_rom0_31_x0x4}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) U515 ( .a ({new_AGEMA_signal_16141, new_AGEMA_signal_16140, mcs_out[128]}), .b ({w0_s2[0], w0_s1[0], w0_s0[0]}), .c ({new_AGEMA_signal_16181, new_AGEMA_signal_16180, y0_1[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U516 ( .a ({new_AGEMA_signal_15187, new_AGEMA_signal_15186, mcs_out[228]}), .b ({w0_s2[100], w0_s1[100], w0_s0[100]}), .c ({new_AGEMA_signal_15297, new_AGEMA_signal_15296, y0_1[100]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U517 ( .a ({new_AGEMA_signal_15701, new_AGEMA_signal_15700, mcs_out[229]}), .b ({w0_s2[101], w0_s1[101], w0_s0[101]}), .c ({new_AGEMA_signal_15797, new_AGEMA_signal_15796, y0_1[101]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U518 ( .a ({new_AGEMA_signal_16117, new_AGEMA_signal_16116, mcs_out[230]}), .b ({w0_s2[102], w0_s1[102], w0_s0[102]}), .c ({new_AGEMA_signal_16183, new_AGEMA_signal_16182, y0_1[102]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U519 ( .a ({new_AGEMA_signal_16115, new_AGEMA_signal_16114, mcs_out[231]}), .b ({w0_s2[103], w0_s1[103], w0_s0[103]}), .c ({new_AGEMA_signal_16185, new_AGEMA_signal_16184, y0_1[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U520 ( .a ({new_AGEMA_signal_16099, new_AGEMA_signal_16098, mcs_out[232]}), .b ({w0_s2[104], w0_s1[104], w0_s0[104]}), .c ({new_AGEMA_signal_16187, new_AGEMA_signal_16186, y0_1[104]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U521 ( .a ({new_AGEMA_signal_14661, new_AGEMA_signal_14660, mcs_out[233]}), .b ({w0_s2[105], w0_s1[105], w0_s0[105]}), .c ({new_AGEMA_signal_14825, new_AGEMA_signal_14824, y0_1[105]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U522 ( .a ({new_AGEMA_signal_15137, new_AGEMA_signal_15136, mcs_out[234]}), .b ({w0_s2[106], w0_s1[106], w0_s0[106]}), .c ({new_AGEMA_signal_15299, new_AGEMA_signal_15298, y0_1[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U523 ( .a ({new_AGEMA_signal_15665, new_AGEMA_signal_15664, mcs_out[235]}), .b ({w0_s2[107], w0_s1[107], w0_s0[107]}), .c ({new_AGEMA_signal_15799, new_AGEMA_signal_15798, y0_1[107]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U524 ( .a ({new_AGEMA_signal_13731, new_AGEMA_signal_13730, mcs_out[236]}), .b ({w0_s2[108], w0_s1[108], w0_s0[108]}), .c ({new_AGEMA_signal_13945, new_AGEMA_signal_13944, y0_1[108]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U525 ( .a ({new_AGEMA_signal_14179, new_AGEMA_signal_14178, mcs_out[237]}), .b ({w0_s2[109], w0_s1[109], w0_s0[109]}), .c ({new_AGEMA_signal_14361, new_AGEMA_signal_14360, y0_1[109]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U526 ( .a ({new_AGEMA_signal_15677, new_AGEMA_signal_15676, mcs_out[138]}), .b ({w0_s2[10], w0_s1[10], w0_s0[10]}), .c ({new_AGEMA_signal_15801, new_AGEMA_signal_15800, y0_1[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U527 ( .a ({new_AGEMA_signal_14177, new_AGEMA_signal_14176, mcs_out[238]}), .b ({w0_s2[110], w0_s1[110], w0_s0[110]}), .c ({new_AGEMA_signal_14363, new_AGEMA_signal_14362, y0_1[110]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U528 ( .a ({new_AGEMA_signal_13725, new_AGEMA_signal_13724, mcs_out[239]}), .b ({w0_s2[111], w0_s1[111], w0_s0[111]}), .c ({new_AGEMA_signal_13947, new_AGEMA_signal_13946, y0_1[111]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U529 ( .a ({new_AGEMA_signal_15601, new_AGEMA_signal_15600, mcs_out[240]}), .b ({w0_s2[112], w0_s1[112], w0_s0[112]}), .c ({new_AGEMA_signal_15803, new_AGEMA_signal_15802, y0_1[112]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U530 ( .a ({new_AGEMA_signal_16061, new_AGEMA_signal_16060, mcs_out[241]}), .b ({w0_s2[113], w0_s1[113], w0_s0[113]}), .c ({new_AGEMA_signal_16189, new_AGEMA_signal_16188, y0_1[113]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U531 ( .a ({new_AGEMA_signal_14559, new_AGEMA_signal_14558, mcs_out[242]}), .b ({w0_s2[114], w0_s1[114], w0_s0[114]}), .c ({new_AGEMA_signal_14827, new_AGEMA_signal_14826, y0_1[114]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U532 ( .a ({new_AGEMA_signal_16059, new_AGEMA_signal_16058, mcs_out[243]}), .b ({w0_s2[115], w0_s1[115], w0_s0[115]}), .c ({new_AGEMA_signal_16191, new_AGEMA_signal_16190, y0_1[115]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U533 ( .a ({new_AGEMA_signal_14997, new_AGEMA_signal_14996, mcs_out[244]}), .b ({w0_s2[116], w0_s1[116], w0_s0[116]}), .c ({new_AGEMA_signal_15301, new_AGEMA_signal_15300, y0_1[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U534 ( .a ({new_AGEMA_signal_15563, new_AGEMA_signal_15562, mcs_out[245]}), .b ({w0_s2[117], w0_s1[117], w0_s0[117]}), .c ({new_AGEMA_signal_15805, new_AGEMA_signal_15804, y0_1[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U535 ( .a ({new_AGEMA_signal_16043, new_AGEMA_signal_16042, mcs_out[246]}), .b ({w0_s2[118], w0_s1[118], w0_s0[118]}), .c ({new_AGEMA_signal_16193, new_AGEMA_signal_16192, y0_1[118]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U536 ( .a ({new_AGEMA_signal_16041, new_AGEMA_signal_16040, mcs_out[247]}), .b ({w0_s2[119], w0_s1[119], w0_s0[119]}), .c ({new_AGEMA_signal_16195, new_AGEMA_signal_16194, y0_1[119]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U537 ( .a ({new_AGEMA_signal_16103, new_AGEMA_signal_16102, mcs_out[139]}), .b ({w0_s2[11], w0_s1[11], w0_s0[11]}), .c ({new_AGEMA_signal_16197, new_AGEMA_signal_16196, y0_1[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U538 ( .a ({new_AGEMA_signal_16025, new_AGEMA_signal_16024, mcs_out[248]}), .b ({w0_s2[120], w0_s1[120], w0_s0[120]}), .c ({new_AGEMA_signal_16199, new_AGEMA_signal_16198, y0_1[120]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U539 ( .a ({new_AGEMA_signal_14463, new_AGEMA_signal_14462, mcs_out[249]}), .b ({w0_s2[121], w0_s1[121], w0_s0[121]}), .c ({new_AGEMA_signal_14829, new_AGEMA_signal_14828, y0_1[121]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U540 ( .a ({new_AGEMA_signal_14947, new_AGEMA_signal_14946, mcs_out[250]}), .b ({w0_s2[122], w0_s1[122], w0_s0[122]}), .c ({new_AGEMA_signal_15303, new_AGEMA_signal_15302, y0_1[122]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U541 ( .a ({new_AGEMA_signal_15527, new_AGEMA_signal_15526, mcs_out[251]}), .b ({w0_s2[123], w0_s1[123], w0_s0[123]}), .c ({new_AGEMA_signal_15807, new_AGEMA_signal_15806, y0_1[123]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U542 ( .a ({new_AGEMA_signal_13513, new_AGEMA_signal_13512, mcs_out[252]}), .b ({w0_s2[124], w0_s1[124], w0_s0[124]}), .c ({new_AGEMA_signal_13949, new_AGEMA_signal_13948, y0_1[124]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U543 ( .a ({new_AGEMA_signal_13993, new_AGEMA_signal_13992, mcs_out[253]}), .b ({w0_s2[125], w0_s1[125], w0_s0[125]}), .c ({new_AGEMA_signal_14365, new_AGEMA_signal_14364, y0_1[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U544 ( .a ({new_AGEMA_signal_13991, new_AGEMA_signal_13990, mcs_out[254]}), .b ({w0_s2[126], w0_s1[126], w0_s0[126]}), .c ({new_AGEMA_signal_14367, new_AGEMA_signal_14366, y0_1[126]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U545 ( .a ({new_AGEMA_signal_13507, new_AGEMA_signal_13506, mcs_out[255]}), .b ({w0_s2[127], w0_s1[127], w0_s0[127]}), .c ({new_AGEMA_signal_13951, new_AGEMA_signal_13950, y0_1[127]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U546 ( .a ({new_AGEMA_signal_16089, new_AGEMA_signal_16088, mcs_out[140]}), .b ({w0_s2[12], w0_s1[12], w0_s0[12]}), .c ({new_AGEMA_signal_16201, new_AGEMA_signal_16200, y0_1[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U547 ( .a ({new_AGEMA_signal_14615, new_AGEMA_signal_14614, mcs_out[141]}), .b ({w0_s2[13], w0_s1[13], w0_s0[13]}), .c ({new_AGEMA_signal_14831, new_AGEMA_signal_14830, y0_1[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U548 ( .a ({new_AGEMA_signal_13733, new_AGEMA_signal_13732, mcs_out[142]}), .b ({w0_s2[14], w0_s1[14], w0_s0[14]}), .c ({new_AGEMA_signal_13953, new_AGEMA_signal_13952, y0_1[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U549 ( .a ({new_AGEMA_signal_15647, new_AGEMA_signal_15646, mcs_out[143]}), .b ({w0_s2[15], w0_s1[15], w0_s0[15]}), .c ({new_AGEMA_signal_15809, new_AGEMA_signal_15808, y0_1[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U550 ( .a ({new_AGEMA_signal_16067, new_AGEMA_signal_16066, mcs_out[144]}), .b ({w0_s2[16], w0_s1[16], w0_s0[16]}), .c ({new_AGEMA_signal_16203, new_AGEMA_signal_16202, y0_1[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U551 ( .a ({new_AGEMA_signal_15057, new_AGEMA_signal_15056, mcs_out[145]}), .b ({w0_s2[17], w0_s1[17], w0_s0[17]}), .c ({new_AGEMA_signal_15305, new_AGEMA_signal_15304, y0_1[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U552 ( .a ({new_AGEMA_signal_16065, new_AGEMA_signal_16064, mcs_out[146]}), .b ({w0_s2[18], w0_s1[18], w0_s0[18]}), .c ({new_AGEMA_signal_16205, new_AGEMA_signal_16204, y0_1[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U553 ( .a ({new_AGEMA_signal_14563, new_AGEMA_signal_14562, mcs_out[147]}), .b ({w0_s2[19], w0_s1[19], w0_s0[19]}), .c ({new_AGEMA_signal_14833, new_AGEMA_signal_14832, y0_1[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U554 ( .a ({new_AGEMA_signal_15247, new_AGEMA_signal_15246, mcs_out[129]}), .b ({w0_s2[1], w0_s1[1], w0_s0[1]}), .c ({new_AGEMA_signal_15307, new_AGEMA_signal_15306, y0_1[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U555 ( .a ({new_AGEMA_signal_15575, new_AGEMA_signal_15574, mcs_out[148]}), .b ({w0_s2[20], w0_s1[20], w0_s0[20]}), .c ({new_AGEMA_signal_15811, new_AGEMA_signal_15810, y0_1[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U556 ( .a ({new_AGEMA_signal_16047, new_AGEMA_signal_16046, mcs_out[149]}), .b ({w0_s2[21], w0_s1[21], w0_s0[21]}), .c ({new_AGEMA_signal_16207, new_AGEMA_signal_16206, y0_1[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U557 ( .a ({new_AGEMA_signal_16045, new_AGEMA_signal_16044, mcs_out[150]}), .b ({w0_s2[22], w0_s1[22], w0_s0[22]}), .c ({new_AGEMA_signal_16209, new_AGEMA_signal_16208, y0_1[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U558 ( .a ({new_AGEMA_signal_15569, new_AGEMA_signal_15568, mcs_out[151]}), .b ({w0_s2[23], w0_s1[23], w0_s0[23]}), .c ({new_AGEMA_signal_15813, new_AGEMA_signal_15812, y0_1[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U559 ( .a ({new_AGEMA_signal_16365, new_AGEMA_signal_16364, mcs_out[152]}), .b ({w0_s2[24], w0_s1[24], w0_s0[24]}), .c ({new_AGEMA_signal_16437, new_AGEMA_signal_16436, y0_1[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U560 ( .a ({new_AGEMA_signal_14473, new_AGEMA_signal_14472, mcs_out[153]}), .b ({w0_s2[25], w0_s1[25], w0_s0[25]}), .c ({new_AGEMA_signal_14835, new_AGEMA_signal_14834, y0_1[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U561 ( .a ({new_AGEMA_signal_15539, new_AGEMA_signal_15538, mcs_out[154]}), .b ({w0_s2[26], w0_s1[26], w0_s0[26]}), .c ({new_AGEMA_signal_15815, new_AGEMA_signal_15814, y0_1[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U562 ( .a ({new_AGEMA_signal_16029, new_AGEMA_signal_16028, mcs_out[155]}), .b ({w0_s2[27], w0_s1[27], w0_s0[27]}), .c ({new_AGEMA_signal_16211, new_AGEMA_signal_16210, y0_1[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U563 ( .a ({new_AGEMA_signal_16015, new_AGEMA_signal_16014, mcs_out[156]}), .b ({w0_s2[28], w0_s1[28], w0_s0[28]}), .c ({new_AGEMA_signal_16213, new_AGEMA_signal_16212, y0_1[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U564 ( .a ({new_AGEMA_signal_14417, new_AGEMA_signal_14416, mcs_out[157]}), .b ({w0_s2[29], w0_s1[29], w0_s0[29]}), .c ({new_AGEMA_signal_14837, new_AGEMA_signal_14836, y0_1[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U565 ( .a ({new_AGEMA_signal_16139, new_AGEMA_signal_16138, mcs_out[130]}), .b ({w0_s2[2], w0_s1[2], w0_s0[2]}), .c ({new_AGEMA_signal_16215, new_AGEMA_signal_16214, y0_1[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U566 ( .a ({new_AGEMA_signal_13515, new_AGEMA_signal_13514, mcs_out[158]}), .b ({w0_s2[30], w0_s1[30], w0_s0[30]}), .c ({new_AGEMA_signal_13955, new_AGEMA_signal_13954, y0_1[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U567 ( .a ({new_AGEMA_signal_15509, new_AGEMA_signal_15508, mcs_out[159]}), .b ({w0_s2[31], w0_s1[31], w0_s0[31]}), .c ({new_AGEMA_signal_15817, new_AGEMA_signal_15816, y0_1[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U568 ( .a ({new_AGEMA_signal_13893, new_AGEMA_signal_13892, mcs_out[160]}), .b ({w0_s2[32], w0_s1[32], w0_s0[32]}), .c ({new_AGEMA_signal_13957, new_AGEMA_signal_13956, y0_1[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U569 ( .a ({new_AGEMA_signal_14319, new_AGEMA_signal_14318, mcs_out[161]}), .b ({w0_s2[33], w0_s1[33], w0_s0[33]}), .c ({new_AGEMA_signal_14369, new_AGEMA_signal_14368, y0_1[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U570 ( .a ({new_AGEMA_signal_14317, new_AGEMA_signal_14316, mcs_out[162]}), .b ({w0_s2[34], w0_s1[34], w0_s0[34]}), .c ({new_AGEMA_signal_14371, new_AGEMA_signal_14370, y0_1[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U571 ( .a ({new_AGEMA_signal_14315, new_AGEMA_signal_14314, mcs_out[163]}), .b ({w0_s2[35], w0_s1[35], w0_s0[35]}), .c ({new_AGEMA_signal_14373, new_AGEMA_signal_14372, y0_1[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U572 ( .a ({new_AGEMA_signal_15195, new_AGEMA_signal_15194, mcs_out[164]}), .b ({w0_s2[36], w0_s1[36], w0_s0[36]}), .c ({new_AGEMA_signal_15309, new_AGEMA_signal_15308, y0_1[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U573 ( .a ({new_AGEMA_signal_13831, new_AGEMA_signal_13830, mcs_out[165]}), .b ({w0_s2[37], w0_s1[37], w0_s0[37]}), .c ({new_AGEMA_signal_13959, new_AGEMA_signal_13958, y0_1[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U574 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, mcs_out[166]}), .b ({w0_s2[38], w0_s1[38], w0_s0[38]}), .c ({new_AGEMA_signal_12977, new_AGEMA_signal_12976, y0_1[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U575 ( .a ({new_AGEMA_signal_14715, new_AGEMA_signal_14714, mcs_out[167]}), .b ({w0_s2[39], w0_s1[39], w0_s0[39]}), .c ({new_AGEMA_signal_14839, new_AGEMA_signal_14838, y0_1[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U576 ( .a ({new_AGEMA_signal_14761, new_AGEMA_signal_14760, mcs_out[131]}), .b ({w0_s2[3], w0_s1[3], w0_s0[3]}), .c ({new_AGEMA_signal_14841, new_AGEMA_signal_14840, y0_1[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U577 ( .a ({new_AGEMA_signal_15671, new_AGEMA_signal_15670, mcs_out[168]}), .b ({w0_s2[40], w0_s1[40], w0_s0[40]}), .c ({new_AGEMA_signal_15819, new_AGEMA_signal_15818, y0_1[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U578 ( .a ({new_AGEMA_signal_15147, new_AGEMA_signal_15146, mcs_out[169]}), .b ({w0_s2[41], w0_s1[41], w0_s0[41]}), .c ({new_AGEMA_signal_15311, new_AGEMA_signal_15310, y0_1[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U579 ( .a ({new_AGEMA_signal_15145, new_AGEMA_signal_15144, mcs_out[170]}), .b ({w0_s2[42], w0_s1[42], w0_s0[42]}), .c ({new_AGEMA_signal_15313, new_AGEMA_signal_15312, y0_1[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U580 ( .a ({new_AGEMA_signal_15143, new_AGEMA_signal_15142, mcs_out[171]}), .b ({w0_s2[43], w0_s1[43], w0_s0[43]}), .c ({new_AGEMA_signal_15315, new_AGEMA_signal_15314, y0_1[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U581 ( .a ({new_AGEMA_signal_16087, new_AGEMA_signal_16086, mcs_out[172]}), .b ({w0_s2[44], w0_s1[44], w0_s0[44]}), .c ({new_AGEMA_signal_16217, new_AGEMA_signal_16216, y0_1[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U582 ( .a ({new_AGEMA_signal_14613, new_AGEMA_signal_14612, mcs_out[173]}), .b ({w0_s2[45], w0_s1[45], w0_s0[45]}), .c ({new_AGEMA_signal_14843, new_AGEMA_signal_14842, y0_1[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U583 ( .a ({new_AGEMA_signal_14611, new_AGEMA_signal_14610, mcs_out[174]}), .b ({w0_s2[46], w0_s1[46], w0_s0[46]}), .c ({new_AGEMA_signal_14845, new_AGEMA_signal_14844, y0_1[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U584 ( .a ({new_AGEMA_signal_15641, new_AGEMA_signal_15640, mcs_out[175]}), .b ({w0_s2[47], w0_s1[47], w0_s0[47]}), .c ({new_AGEMA_signal_15821, new_AGEMA_signal_15820, y0_1[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U585 ( .a ({new_AGEMA_signal_13675, new_AGEMA_signal_13674, mcs_out[176]}), .b ({w0_s2[48], w0_s1[48], w0_s0[48]}), .c ({new_AGEMA_signal_13961, new_AGEMA_signal_13960, y0_1[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U586 ( .a ({new_AGEMA_signal_14133, new_AGEMA_signal_14132, mcs_out[177]}), .b ({w0_s2[49], w0_s1[49], w0_s0[49]}), .c ({new_AGEMA_signal_14375, new_AGEMA_signal_14374, y0_1[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U587 ( .a ({new_AGEMA_signal_15713, new_AGEMA_signal_15712, mcs_out[132]}), .b ({w0_s2[4], w0_s1[4], w0_s0[4]}), .c ({new_AGEMA_signal_15823, new_AGEMA_signal_15822, y0_1[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U588 ( .a ({new_AGEMA_signal_14131, new_AGEMA_signal_14130, mcs_out[178]}), .b ({w0_s2[50], w0_s1[50], w0_s0[50]}), .c ({new_AGEMA_signal_14377, new_AGEMA_signal_14376, y0_1[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U589 ( .a ({new_AGEMA_signal_14129, new_AGEMA_signal_14128, mcs_out[179]}), .b ({w0_s2[51], w0_s1[51], w0_s0[51]}), .c ({new_AGEMA_signal_14379, new_AGEMA_signal_14378, y0_1[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U590 ( .a ({new_AGEMA_signal_15005, new_AGEMA_signal_15004, mcs_out[180]}), .b ({w0_s2[52], w0_s1[52], w0_s0[52]}), .c ({new_AGEMA_signal_15317, new_AGEMA_signal_15316, y0_1[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U591 ( .a ({new_AGEMA_signal_13613, new_AGEMA_signal_13612, mcs_out[181]}), .b ({w0_s2[53], w0_s1[53], w0_s0[53]}), .c ({new_AGEMA_signal_13963, new_AGEMA_signal_13962, y0_1[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U592 ( .a ({new_AGEMA_signal_12547, new_AGEMA_signal_12546, mcs_out[182]}), .b ({w0_s2[54], w0_s1[54], w0_s0[54]}), .c ({new_AGEMA_signal_12979, new_AGEMA_signal_12978, y0_1[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U593 ( .a ({new_AGEMA_signal_14517, new_AGEMA_signal_14516, mcs_out[183]}), .b ({w0_s2[55], w0_s1[55], w0_s0[55]}), .c ({new_AGEMA_signal_14847, new_AGEMA_signal_14846, y0_1[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U594 ( .a ({new_AGEMA_signal_15533, new_AGEMA_signal_15532, mcs_out[184]}), .b ({w0_s2[56], w0_s1[56], w0_s0[56]}), .c ({new_AGEMA_signal_15825, new_AGEMA_signal_15824, y0_1[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U595 ( .a ({new_AGEMA_signal_14957, new_AGEMA_signal_14956, mcs_out[185]}), .b ({w0_s2[57], w0_s1[57], w0_s0[57]}), .c ({new_AGEMA_signal_15319, new_AGEMA_signal_15318, y0_1[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U596 ( .a ({new_AGEMA_signal_14955, new_AGEMA_signal_14954, mcs_out[186]}), .b ({w0_s2[58], w0_s1[58], w0_s0[58]}), .c ({new_AGEMA_signal_15321, new_AGEMA_signal_15320, y0_1[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U597 ( .a ({new_AGEMA_signal_14953, new_AGEMA_signal_14952, mcs_out[187]}), .b ({w0_s2[59], w0_s1[59], w0_s0[59]}), .c ({new_AGEMA_signal_15323, new_AGEMA_signal_15322, y0_1[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U598 ( .a ({new_AGEMA_signal_16121, new_AGEMA_signal_16120, mcs_out[133]}), .b ({w0_s2[5], w0_s1[5], w0_s0[5]}), .c ({new_AGEMA_signal_16219, new_AGEMA_signal_16218, y0_1[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U599 ( .a ({new_AGEMA_signal_16013, new_AGEMA_signal_16012, mcs_out[188]}), .b ({w0_s2[60], w0_s1[60], w0_s0[60]}), .c ({new_AGEMA_signal_16221, new_AGEMA_signal_16220, y0_1[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U600 ( .a ({new_AGEMA_signal_14415, new_AGEMA_signal_14414, mcs_out[189]}), .b ({w0_s2[61], w0_s1[61], w0_s0[61]}), .c ({new_AGEMA_signal_14849, new_AGEMA_signal_14848, y0_1[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U601 ( .a ({new_AGEMA_signal_14413, new_AGEMA_signal_14412, mcs_out[190]}), .b ({w0_s2[62], w0_s1[62], w0_s0[62]}), .c ({new_AGEMA_signal_14851, new_AGEMA_signal_14850, y0_1[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U602 ( .a ({new_AGEMA_signal_15503, new_AGEMA_signal_15502, mcs_out[191]}), .b ({w0_s2[63], w0_s1[63], w0_s0[63]}), .c ({new_AGEMA_signal_15827, new_AGEMA_signal_15826, y0_1[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U603 ( .a ({new_AGEMA_signal_16137, new_AGEMA_signal_16136, mcs_out[192]}), .b ({w0_s2[64], w0_s1[64], w0_s0[64]}), .c ({new_AGEMA_signal_16223, new_AGEMA_signal_16222, y0_1[64]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U604 ( .a ({new_AGEMA_signal_15745, new_AGEMA_signal_15744, mcs_out[193]}), .b ({w0_s2[65], w0_s1[65], w0_s0[65]}), .c ({new_AGEMA_signal_15829, new_AGEMA_signal_15828, y0_1[65]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U605 ( .a ({new_AGEMA_signal_15743, new_AGEMA_signal_15742, mcs_out[194]}), .b ({w0_s2[66], w0_s1[66], w0_s0[66]}), .c ({new_AGEMA_signal_15831, new_AGEMA_signal_15830, y0_1[66]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U606 ( .a ({new_AGEMA_signal_15741, new_AGEMA_signal_15740, mcs_out[195]}), .b ({w0_s2[67], w0_s1[67], w0_s0[67]}), .c ({new_AGEMA_signal_15833, new_AGEMA_signal_15832, y0_1[67]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U607 ( .a ({new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs_out[196]}), .b ({w0_s2[68], w0_s1[68], w0_s0[68]}), .c ({new_AGEMA_signal_15835, new_AGEMA_signal_15834, y0_1[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U608 ( .a ({new_AGEMA_signal_15191, new_AGEMA_signal_15190, mcs_out[197]}), .b ({w0_s2[69], w0_s1[69], w0_s0[69]}), .c ({new_AGEMA_signal_15325, new_AGEMA_signal_15324, y0_1[69]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U609 ( .a ({new_AGEMA_signal_16119, new_AGEMA_signal_16118, mcs_out[134]}), .b ({w0_s2[6], w0_s1[6], w0_s0[6]}), .c ({new_AGEMA_signal_16225, new_AGEMA_signal_16224, y0_1[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U610 ( .a ({new_AGEMA_signal_14711, new_AGEMA_signal_14710, mcs_out[198]}), .b ({w0_s2[70], w0_s1[70], w0_s0[70]}), .c ({new_AGEMA_signal_14853, new_AGEMA_signal_14852, y0_1[70]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U611 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, mcs_out[199]}), .b ({w0_s2[71], w0_s1[71], w0_s0[71]}), .c ({new_AGEMA_signal_15837, new_AGEMA_signal_15836, y0_1[71]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U612 ( .a ({new_AGEMA_signal_16469, new_AGEMA_signal_16468, mcs_out[200]}), .b ({w0_s2[72], w0_s1[72], w0_s0[72]}), .c ({new_AGEMA_signal_16545, new_AGEMA_signal_16544, y0_1[72]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U613 ( .a ({new_AGEMA_signal_14221, new_AGEMA_signal_14220, mcs_out[201]}), .b ({w0_s2[73], w0_s1[73], w0_s0[73]}), .c ({new_AGEMA_signal_14381, new_AGEMA_signal_14380, y0_1[73]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U614 ( .a ({new_AGEMA_signal_15141, new_AGEMA_signal_15140, mcs_out[202]}), .b ({w0_s2[74], w0_s1[74], w0_s0[74]}), .c ({new_AGEMA_signal_15327, new_AGEMA_signal_15326, y0_1[74]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U615 ( .a ({new_AGEMA_signal_16101, new_AGEMA_signal_16100, mcs_out[203]}), .b ({w0_s2[75], w0_s1[75], w0_s0[75]}), .c ({new_AGEMA_signal_16227, new_AGEMA_signal_16226, y0_1[75]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U616 ( .a ({new_AGEMA_signal_16085, new_AGEMA_signal_16084, mcs_out[204]}), .b ({w0_s2[76], w0_s1[76], w0_s0[76]}), .c ({new_AGEMA_signal_16229, new_AGEMA_signal_16228, y0_1[76]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U617 ( .a ({new_AGEMA_signal_16083, new_AGEMA_signal_16082, mcs_out[205]}), .b ({w0_s2[77], w0_s1[77], w0_s0[77]}), .c ({new_AGEMA_signal_16231, new_AGEMA_signal_16230, y0_1[77]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U618 ( .a ({new_AGEMA_signal_16081, new_AGEMA_signal_16080, mcs_out[206]}), .b ({w0_s2[78], w0_s1[78], w0_s0[78]}), .c ({new_AGEMA_signal_16233, new_AGEMA_signal_16232, y0_1[78]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U619 ( .a ({new_AGEMA_signal_16079, new_AGEMA_signal_16078, mcs_out[207]}), .b ({w0_s2[79], w0_s1[79], w0_s0[79]}), .c ({new_AGEMA_signal_16235, new_AGEMA_signal_16234, y0_1[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U620 ( .a ({new_AGEMA_signal_15707, new_AGEMA_signal_15706, mcs_out[135]}), .b ({w0_s2[7], w0_s1[7], w0_s0[7]}), .c ({new_AGEMA_signal_15839, new_AGEMA_signal_15838, y0_1[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U621 ( .a ({new_AGEMA_signal_16063, new_AGEMA_signal_16062, mcs_out[208]}), .b ({w0_s2[80], w0_s1[80], w0_s0[80]}), .c ({new_AGEMA_signal_16237, new_AGEMA_signal_16236, y0_1[80]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U622 ( .a ({new_AGEMA_signal_15607, new_AGEMA_signal_15606, mcs_out[209]}), .b ({w0_s2[81], w0_s1[81], w0_s0[81]}), .c ({new_AGEMA_signal_15841, new_AGEMA_signal_15840, y0_1[81]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U623 ( .a ({new_AGEMA_signal_15605, new_AGEMA_signal_15604, mcs_out[210]}), .b ({w0_s2[82], w0_s1[82], w0_s0[82]}), .c ({new_AGEMA_signal_15843, new_AGEMA_signal_15842, y0_1[82]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U624 ( .a ({new_AGEMA_signal_15603, new_AGEMA_signal_15602, mcs_out[211]}), .b ({w0_s2[83], w0_s1[83], w0_s0[83]}), .c ({new_AGEMA_signal_15845, new_AGEMA_signal_15844, y0_1[83]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U625 ( .a ({new_AGEMA_signal_15567, new_AGEMA_signal_15566, mcs_out[212]}), .b ({w0_s2[84], w0_s1[84], w0_s0[84]}), .c ({new_AGEMA_signal_15847, new_AGEMA_signal_15846, y0_1[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U626 ( .a ({new_AGEMA_signal_15001, new_AGEMA_signal_15000, mcs_out[213]}), .b ({w0_s2[85], w0_s1[85], w0_s0[85]}), .c ({new_AGEMA_signal_15329, new_AGEMA_signal_15328, y0_1[85]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U627 ( .a ({new_AGEMA_signal_14513, new_AGEMA_signal_14512, mcs_out[214]}), .b ({w0_s2[86], w0_s1[86], w0_s0[86]}), .c ({new_AGEMA_signal_14855, new_AGEMA_signal_14854, y0_1[86]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U628 ( .a ({new_AGEMA_signal_15565, new_AGEMA_signal_15564, mcs_out[215]}), .b ({w0_s2[87], w0_s1[87], w0_s0[87]}), .c ({new_AGEMA_signal_15849, new_AGEMA_signal_15848, y0_1[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U629 ( .a ({new_AGEMA_signal_16465, new_AGEMA_signal_16464, mcs_out[216]}), .b ({w0_s2[88], w0_s1[88], w0_s0[88]}), .c ({new_AGEMA_signal_16547, new_AGEMA_signal_16546, y0_1[88]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U630 ( .a ({new_AGEMA_signal_14035, new_AGEMA_signal_14034, mcs_out[217]}), .b ({w0_s2[89], w0_s1[89], w0_s0[89]}), .c ({new_AGEMA_signal_14383, new_AGEMA_signal_14382, y0_1[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U631 ( .a ({new_AGEMA_signal_16377, new_AGEMA_signal_16376, mcs_out[136]}), .b ({w0_s2[8], w0_s1[8], w0_s0[8]}), .c ({new_AGEMA_signal_16439, new_AGEMA_signal_16438, y0_1[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U632 ( .a ({new_AGEMA_signal_14951, new_AGEMA_signal_14950, mcs_out[218]}), .b ({w0_s2[90], w0_s1[90], w0_s0[90]}), .c ({new_AGEMA_signal_15331, new_AGEMA_signal_15330, y0_1[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U633 ( .a ({new_AGEMA_signal_16027, new_AGEMA_signal_16026, mcs_out[219]}), .b ({w0_s2[91], w0_s1[91], w0_s0[91]}), .c ({new_AGEMA_signal_16239, new_AGEMA_signal_16238, y0_1[91]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U634 ( .a ({new_AGEMA_signal_16011, new_AGEMA_signal_16010, mcs_out[220]}), .b ({w0_s2[92], w0_s1[92], w0_s0[92]}), .c ({new_AGEMA_signal_16241, new_AGEMA_signal_16240, y0_1[92]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U635 ( .a ({new_AGEMA_signal_16009, new_AGEMA_signal_16008, mcs_out[221]}), .b ({w0_s2[93], w0_s1[93], w0_s0[93]}), .c ({new_AGEMA_signal_16243, new_AGEMA_signal_16242, y0_1[93]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U636 ( .a ({new_AGEMA_signal_16007, new_AGEMA_signal_16006, mcs_out[222]}), .b ({w0_s2[94], w0_s1[94], w0_s0[94]}), .c ({new_AGEMA_signal_16245, new_AGEMA_signal_16244, y0_1[94]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U637 ( .a ({new_AGEMA_signal_16005, new_AGEMA_signal_16004, mcs_out[223]}), .b ({w0_s2[95], w0_s1[95], w0_s0[95]}), .c ({new_AGEMA_signal_16247, new_AGEMA_signal_16246, y0_1[95]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U638 ( .a ({new_AGEMA_signal_15739, new_AGEMA_signal_15738, mcs_out[224]}), .b ({w0_s2[96], w0_s1[96], w0_s0[96]}), .c ({new_AGEMA_signal_15851, new_AGEMA_signal_15850, y0_1[96]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U639 ( .a ({new_AGEMA_signal_16135, new_AGEMA_signal_16134, mcs_out[225]}), .b ({w0_s2[97], w0_s1[97], w0_s0[97]}), .c ({new_AGEMA_signal_16249, new_AGEMA_signal_16248, y0_1[97]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U640 ( .a ({new_AGEMA_signal_14757, new_AGEMA_signal_14756, mcs_out[226]}), .b ({w0_s2[98], w0_s1[98], w0_s0[98]}), .c ({new_AGEMA_signal_14857, new_AGEMA_signal_14856, y0_1[98]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U641 ( .a ({new_AGEMA_signal_16133, new_AGEMA_signal_16132, mcs_out[227]}), .b ({w0_s2[99], w0_s1[99], w0_s0[99]}), .c ({new_AGEMA_signal_16251, new_AGEMA_signal_16250, y0_1[99]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U642 ( .a ({new_AGEMA_signal_14671, new_AGEMA_signal_14670, mcs_out[137]}), .b ({w0_s2[9], w0_s1[9], w0_s0[9]}), .c ({new_AGEMA_signal_14859, new_AGEMA_signal_14858, y0_1[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U643 ( .a ({temp_s2[0], temp_s1[0], temp_s0[0]}), .b ({temp_next_s2[0], temp_next_s1[0], temp_next_s0[0]}), .c ({y1_s2[0], y1_s1[0], y1_s0[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U644 ( .a ({temp_s2[100], temp_s1[100], temp_s0[100]}), .b ({temp_next_s2[100], temp_next_s1[100], temp_next_s0[100]}), .c ({y1_s2[100], y1_s1[100], y1_s0[100]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U645 ( .a ({temp_s2[101], temp_s1[101], temp_s0[101]}), .b ({temp_next_s2[101], temp_next_s1[101], temp_next_s0[101]}), .c ({y1_s2[101], y1_s1[101], y1_s0[101]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U646 ( .a ({temp_s2[102], temp_s1[102], temp_s0[102]}), .b ({temp_next_s2[102], temp_next_s1[102], temp_next_s0[102]}), .c ({y1_s2[102], y1_s1[102], y1_s0[102]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U647 ( .a ({temp_s2[103], temp_s1[103], temp_s0[103]}), .b ({temp_next_s2[103], temp_next_s1[103], temp_next_s0[103]}), .c ({y1_s2[103], y1_s1[103], y1_s0[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U648 ( .a ({temp_s2[104], temp_s1[104], temp_s0[104]}), .b ({temp_next_s2[104], temp_next_s1[104], temp_next_s0[104]}), .c ({y1_s2[104], y1_s1[104], y1_s0[104]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U649 ( .a ({temp_s2[105], temp_s1[105], temp_s0[105]}), .b ({temp_next_s2[105], temp_next_s1[105], temp_next_s0[105]}), .c ({y1_s2[105], y1_s1[105], y1_s0[105]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U650 ( .a ({temp_s2[106], temp_s1[106], temp_s0[106]}), .b ({temp_next_s2[106], temp_next_s1[106], temp_next_s0[106]}), .c ({y1_s2[106], y1_s1[106], y1_s0[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U651 ( .a ({temp_s2[107], temp_s1[107], temp_s0[107]}), .b ({temp_next_s2[107], temp_next_s1[107], temp_next_s0[107]}), .c ({y1_s2[107], y1_s1[107], y1_s0[107]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U652 ( .a ({temp_s2[108], temp_s1[108], temp_s0[108]}), .b ({temp_next_s2[108], temp_next_s1[108], temp_next_s0[108]}), .c ({y1_s2[108], y1_s1[108], y1_s0[108]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U653 ( .a ({temp_s2[109], temp_s1[109], temp_s0[109]}), .b ({temp_next_s2[109], temp_next_s1[109], temp_next_s0[109]}), .c ({y1_s2[109], y1_s1[109], y1_s0[109]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U654 ( .a ({temp_s2[10], temp_s1[10], temp_s0[10]}), .b ({temp_next_s2[10], temp_next_s1[10], temp_next_s0[10]}), .c ({y1_s2[10], y1_s1[10], y1_s0[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U655 ( .a ({temp_s2[110], temp_s1[110], temp_s0[110]}), .b ({temp_next_s2[110], temp_next_s1[110], temp_next_s0[110]}), .c ({y1_s2[110], y1_s1[110], y1_s0[110]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U656 ( .a ({temp_s2[111], temp_s1[111], temp_s0[111]}), .b ({temp_next_s2[111], temp_next_s1[111], temp_next_s0[111]}), .c ({y1_s2[111], y1_s1[111], y1_s0[111]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U657 ( .a ({temp_s2[112], temp_s1[112], temp_s0[112]}), .b ({temp_next_s2[112], temp_next_s1[112], temp_next_s0[112]}), .c ({y1_s2[112], y1_s1[112], y1_s0[112]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U658 ( .a ({temp_s2[113], temp_s1[113], temp_s0[113]}), .b ({temp_next_s2[113], temp_next_s1[113], temp_next_s0[113]}), .c ({y1_s2[113], y1_s1[113], y1_s0[113]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U659 ( .a ({temp_s2[114], temp_s1[114], temp_s0[114]}), .b ({temp_next_s2[114], temp_next_s1[114], temp_next_s0[114]}), .c ({y1_s2[114], y1_s1[114], y1_s0[114]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U660 ( .a ({temp_s2[115], temp_s1[115], temp_s0[115]}), .b ({temp_next_s2[115], temp_next_s1[115], temp_next_s0[115]}), .c ({y1_s2[115], y1_s1[115], y1_s0[115]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U661 ( .a ({temp_s2[116], temp_s1[116], temp_s0[116]}), .b ({temp_next_s2[116], temp_next_s1[116], temp_next_s0[116]}), .c ({y1_s2[116], y1_s1[116], y1_s0[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U662 ( .a ({temp_s2[117], temp_s1[117], temp_s0[117]}), .b ({temp_next_s2[117], temp_next_s1[117], temp_next_s0[117]}), .c ({y1_s2[117], y1_s1[117], y1_s0[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U663 ( .a ({temp_s2[118], temp_s1[118], temp_s0[118]}), .b ({temp_next_s2[118], temp_next_s1[118], temp_next_s0[118]}), .c ({y1_s2[118], y1_s1[118], y1_s0[118]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U664 ( .a ({temp_s2[119], temp_s1[119], temp_s0[119]}), .b ({temp_next_s2[119], temp_next_s1[119], temp_next_s0[119]}), .c ({y1_s2[119], y1_s1[119], y1_s0[119]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U665 ( .a ({temp_s2[11], temp_s1[11], temp_s0[11]}), .b ({temp_next_s2[11], temp_next_s1[11], temp_next_s0[11]}), .c ({y1_s2[11], y1_s1[11], y1_s0[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U666 ( .a ({temp_s2[120], temp_s1[120], temp_s0[120]}), .b ({temp_next_s2[120], temp_next_s1[120], temp_next_s0[120]}), .c ({y1_s2[120], y1_s1[120], y1_s0[120]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U667 ( .a ({temp_s2[121], temp_s1[121], temp_s0[121]}), .b ({temp_next_s2[121], temp_next_s1[121], temp_next_s0[121]}), .c ({y1_s2[121], y1_s1[121], y1_s0[121]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U668 ( .a ({temp_s2[122], temp_s1[122], temp_s0[122]}), .b ({temp_next_s2[122], temp_next_s1[122], temp_next_s0[122]}), .c ({y1_s2[122], y1_s1[122], y1_s0[122]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U669 ( .a ({temp_s2[123], temp_s1[123], temp_s0[123]}), .b ({temp_next_s2[123], temp_next_s1[123], temp_next_s0[123]}), .c ({y1_s2[123], y1_s1[123], y1_s0[123]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U670 ( .a ({temp_s2[124], temp_s1[124], temp_s0[124]}), .b ({temp_next_s2[124], temp_next_s1[124], temp_next_s0[124]}), .c ({y1_s2[124], y1_s1[124], y1_s0[124]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U671 ( .a ({temp_s2[125], temp_s1[125], temp_s0[125]}), .b ({temp_next_s2[125], temp_next_s1[125], temp_next_s0[125]}), .c ({y1_s2[125], y1_s1[125], y1_s0[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U672 ( .a ({temp_s2[126], temp_s1[126], temp_s0[126]}), .b ({temp_next_s2[126], temp_next_s1[126], temp_next_s0[126]}), .c ({y1_s2[126], y1_s1[126], y1_s0[126]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U673 ( .a ({temp_s2[127], temp_s1[127], temp_s0[127]}), .b ({temp_next_s2[127], temp_next_s1[127], temp_next_s0[127]}), .c ({y1_s2[127], y1_s1[127], y1_s0[127]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U674 ( .a ({temp_s2[12], temp_s1[12], temp_s0[12]}), .b ({temp_next_s2[12], temp_next_s1[12], temp_next_s0[12]}), .c ({y1_s2[12], y1_s1[12], y1_s0[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U675 ( .a ({temp_s2[13], temp_s1[13], temp_s0[13]}), .b ({temp_next_s2[13], temp_next_s1[13], temp_next_s0[13]}), .c ({y1_s2[13], y1_s1[13], y1_s0[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U676 ( .a ({temp_s2[14], temp_s1[14], temp_s0[14]}), .b ({temp_next_s2[14], temp_next_s1[14], temp_next_s0[14]}), .c ({y1_s2[14], y1_s1[14], y1_s0[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U677 ( .a ({temp_s2[15], temp_s1[15], temp_s0[15]}), .b ({temp_next_s2[15], temp_next_s1[15], temp_next_s0[15]}), .c ({y1_s2[15], y1_s1[15], y1_s0[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U678 ( .a ({temp_s2[16], temp_s1[16], temp_s0[16]}), .b ({temp_next_s2[16], temp_next_s1[16], temp_next_s0[16]}), .c ({y1_s2[16], y1_s1[16], y1_s0[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U679 ( .a ({temp_s2[17], temp_s1[17], temp_s0[17]}), .b ({temp_next_s2[17], temp_next_s1[17], temp_next_s0[17]}), .c ({y1_s2[17], y1_s1[17], y1_s0[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U680 ( .a ({temp_s2[18], temp_s1[18], temp_s0[18]}), .b ({temp_next_s2[18], temp_next_s1[18], temp_next_s0[18]}), .c ({y1_s2[18], y1_s1[18], y1_s0[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U681 ( .a ({temp_s2[19], temp_s1[19], temp_s0[19]}), .b ({temp_next_s2[19], temp_next_s1[19], temp_next_s0[19]}), .c ({y1_s2[19], y1_s1[19], y1_s0[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U682 ( .a ({temp_s2[1], temp_s1[1], temp_s0[1]}), .b ({temp_next_s2[1], temp_next_s1[1], temp_next_s0[1]}), .c ({y1_s2[1], y1_s1[1], y1_s0[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U683 ( .a ({temp_s2[20], temp_s1[20], temp_s0[20]}), .b ({temp_next_s2[20], temp_next_s1[20], temp_next_s0[20]}), .c ({y1_s2[20], y1_s1[20], y1_s0[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U684 ( .a ({temp_s2[21], temp_s1[21], temp_s0[21]}), .b ({temp_next_s2[21], temp_next_s1[21], temp_next_s0[21]}), .c ({y1_s2[21], y1_s1[21], y1_s0[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U685 ( .a ({temp_s2[22], temp_s1[22], temp_s0[22]}), .b ({temp_next_s2[22], temp_next_s1[22], temp_next_s0[22]}), .c ({y1_s2[22], y1_s1[22], y1_s0[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U686 ( .a ({temp_s2[23], temp_s1[23], temp_s0[23]}), .b ({temp_next_s2[23], temp_next_s1[23], temp_next_s0[23]}), .c ({y1_s2[23], y1_s1[23], y1_s0[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U687 ( .a ({temp_s2[24], temp_s1[24], temp_s0[24]}), .b ({temp_next_s2[24], temp_next_s1[24], temp_next_s0[24]}), .c ({y1_s2[24], y1_s1[24], y1_s0[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U688 ( .a ({temp_s2[25], temp_s1[25], temp_s0[25]}), .b ({temp_next_s2[25], temp_next_s1[25], temp_next_s0[25]}), .c ({y1_s2[25], y1_s1[25], y1_s0[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U689 ( .a ({temp_s2[26], temp_s1[26], temp_s0[26]}), .b ({temp_next_s2[26], temp_next_s1[26], temp_next_s0[26]}), .c ({y1_s2[26], y1_s1[26], y1_s0[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U690 ( .a ({temp_s2[27], temp_s1[27], temp_s0[27]}), .b ({temp_next_s2[27], temp_next_s1[27], temp_next_s0[27]}), .c ({y1_s2[27], y1_s1[27], y1_s0[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U691 ( .a ({temp_s2[28], temp_s1[28], temp_s0[28]}), .b ({temp_next_s2[28], temp_next_s1[28], temp_next_s0[28]}), .c ({y1_s2[28], y1_s1[28], y1_s0[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U692 ( .a ({temp_s2[29], temp_s1[29], temp_s0[29]}), .b ({temp_next_s2[29], temp_next_s1[29], temp_next_s0[29]}), .c ({y1_s2[29], y1_s1[29], y1_s0[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U693 ( .a ({temp_s2[2], temp_s1[2], temp_s0[2]}), .b ({temp_next_s2[2], temp_next_s1[2], temp_next_s0[2]}), .c ({y1_s2[2], y1_s1[2], y1_s0[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U694 ( .a ({temp_s2[30], temp_s1[30], temp_s0[30]}), .b ({temp_next_s2[30], temp_next_s1[30], temp_next_s0[30]}), .c ({y1_s2[30], y1_s1[30], y1_s0[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U695 ( .a ({temp_s2[31], temp_s1[31], temp_s0[31]}), .b ({temp_next_s2[31], temp_next_s1[31], temp_next_s0[31]}), .c ({y1_s2[31], y1_s1[31], y1_s0[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U696 ( .a ({temp_s2[32], temp_s1[32], temp_s0[32]}), .b ({temp_next_s2[32], temp_next_s1[32], temp_next_s0[32]}), .c ({y1_s2[32], y1_s1[32], y1_s0[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U697 ( .a ({temp_s2[33], temp_s1[33], temp_s0[33]}), .b ({temp_next_s2[33], temp_next_s1[33], temp_next_s0[33]}), .c ({y1_s2[33], y1_s1[33], y1_s0[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U698 ( .a ({temp_s2[34], temp_s1[34], temp_s0[34]}), .b ({temp_next_s2[34], temp_next_s1[34], temp_next_s0[34]}), .c ({y1_s2[34], y1_s1[34], y1_s0[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U699 ( .a ({temp_s2[35], temp_s1[35], temp_s0[35]}), .b ({temp_next_s2[35], temp_next_s1[35], temp_next_s0[35]}), .c ({y1_s2[35], y1_s1[35], y1_s0[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U700 ( .a ({temp_s2[36], temp_s1[36], temp_s0[36]}), .b ({temp_next_s2[36], temp_next_s1[36], temp_next_s0[36]}), .c ({y1_s2[36], y1_s1[36], y1_s0[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U701 ( .a ({temp_s2[37], temp_s1[37], temp_s0[37]}), .b ({temp_next_s2[37], temp_next_s1[37], temp_next_s0[37]}), .c ({y1_s2[37], y1_s1[37], y1_s0[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U702 ( .a ({temp_s2[38], temp_s1[38], temp_s0[38]}), .b ({temp_next_s2[38], temp_next_s1[38], temp_next_s0[38]}), .c ({y1_s2[38], y1_s1[38], y1_s0[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U703 ( .a ({temp_s2[39], temp_s1[39], temp_s0[39]}), .b ({temp_next_s2[39], temp_next_s1[39], temp_next_s0[39]}), .c ({y1_s2[39], y1_s1[39], y1_s0[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U704 ( .a ({temp_s2[3], temp_s1[3], temp_s0[3]}), .b ({temp_next_s2[3], temp_next_s1[3], temp_next_s0[3]}), .c ({y1_s2[3], y1_s1[3], y1_s0[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U705 ( .a ({temp_s2[40], temp_s1[40], temp_s0[40]}), .b ({temp_next_s2[40], temp_next_s1[40], temp_next_s0[40]}), .c ({y1_s2[40], y1_s1[40], y1_s0[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U706 ( .a ({temp_s2[41], temp_s1[41], temp_s0[41]}), .b ({temp_next_s2[41], temp_next_s1[41], temp_next_s0[41]}), .c ({y1_s2[41], y1_s1[41], y1_s0[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U707 ( .a ({temp_s2[42], temp_s1[42], temp_s0[42]}), .b ({temp_next_s2[42], temp_next_s1[42], temp_next_s0[42]}), .c ({y1_s2[42], y1_s1[42], y1_s0[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U708 ( .a ({temp_s2[43], temp_s1[43], temp_s0[43]}), .b ({temp_next_s2[43], temp_next_s1[43], temp_next_s0[43]}), .c ({y1_s2[43], y1_s1[43], y1_s0[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U709 ( .a ({temp_s2[44], temp_s1[44], temp_s0[44]}), .b ({temp_next_s2[44], temp_next_s1[44], temp_next_s0[44]}), .c ({y1_s2[44], y1_s1[44], y1_s0[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U710 ( .a ({temp_s2[45], temp_s1[45], temp_s0[45]}), .b ({temp_next_s2[45], temp_next_s1[45], temp_next_s0[45]}), .c ({y1_s2[45], y1_s1[45], y1_s0[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U711 ( .a ({temp_s2[46], temp_s1[46], temp_s0[46]}), .b ({temp_next_s2[46], temp_next_s1[46], temp_next_s0[46]}), .c ({y1_s2[46], y1_s1[46], y1_s0[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U712 ( .a ({temp_s2[47], temp_s1[47], temp_s0[47]}), .b ({temp_next_s2[47], temp_next_s1[47], temp_next_s0[47]}), .c ({y1_s2[47], y1_s1[47], y1_s0[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U713 ( .a ({temp_s2[48], temp_s1[48], temp_s0[48]}), .b ({temp_next_s2[48], temp_next_s1[48], temp_next_s0[48]}), .c ({y1_s2[48], y1_s1[48], y1_s0[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U714 ( .a ({temp_s2[49], temp_s1[49], temp_s0[49]}), .b ({temp_next_s2[49], temp_next_s1[49], temp_next_s0[49]}), .c ({y1_s2[49], y1_s1[49], y1_s0[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U715 ( .a ({temp_s2[4], temp_s1[4], temp_s0[4]}), .b ({temp_next_s2[4], temp_next_s1[4], temp_next_s0[4]}), .c ({y1_s2[4], y1_s1[4], y1_s0[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U716 ( .a ({temp_s2[50], temp_s1[50], temp_s0[50]}), .b ({temp_next_s2[50], temp_next_s1[50], temp_next_s0[50]}), .c ({y1_s2[50], y1_s1[50], y1_s0[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U717 ( .a ({temp_s2[51], temp_s1[51], temp_s0[51]}), .b ({temp_next_s2[51], temp_next_s1[51], temp_next_s0[51]}), .c ({y1_s2[51], y1_s1[51], y1_s0[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U718 ( .a ({temp_s2[52], temp_s1[52], temp_s0[52]}), .b ({temp_next_s2[52], temp_next_s1[52], temp_next_s0[52]}), .c ({y1_s2[52], y1_s1[52], y1_s0[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U719 ( .a ({temp_s2[53], temp_s1[53], temp_s0[53]}), .b ({temp_next_s2[53], temp_next_s1[53], temp_next_s0[53]}), .c ({y1_s2[53], y1_s1[53], y1_s0[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U720 ( .a ({temp_s2[54], temp_s1[54], temp_s0[54]}), .b ({temp_next_s2[54], temp_next_s1[54], temp_next_s0[54]}), .c ({y1_s2[54], y1_s1[54], y1_s0[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U721 ( .a ({temp_s2[55], temp_s1[55], temp_s0[55]}), .b ({temp_next_s2[55], temp_next_s1[55], temp_next_s0[55]}), .c ({y1_s2[55], y1_s1[55], y1_s0[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U722 ( .a ({temp_s2[56], temp_s1[56], temp_s0[56]}), .b ({temp_next_s2[56], temp_next_s1[56], temp_next_s0[56]}), .c ({y1_s2[56], y1_s1[56], y1_s0[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U723 ( .a ({temp_s2[57], temp_s1[57], temp_s0[57]}), .b ({temp_next_s2[57], temp_next_s1[57], temp_next_s0[57]}), .c ({y1_s2[57], y1_s1[57], y1_s0[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U724 ( .a ({temp_s2[58], temp_s1[58], temp_s0[58]}), .b ({temp_next_s2[58], temp_next_s1[58], temp_next_s0[58]}), .c ({y1_s2[58], y1_s1[58], y1_s0[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U725 ( .a ({temp_s2[59], temp_s1[59], temp_s0[59]}), .b ({temp_next_s2[59], temp_next_s1[59], temp_next_s0[59]}), .c ({y1_s2[59], y1_s1[59], y1_s0[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U726 ( .a ({temp_s2[5], temp_s1[5], temp_s0[5]}), .b ({temp_next_s2[5], temp_next_s1[5], temp_next_s0[5]}), .c ({y1_s2[5], y1_s1[5], y1_s0[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U727 ( .a ({temp_s2[60], temp_s1[60], temp_s0[60]}), .b ({temp_next_s2[60], temp_next_s1[60], temp_next_s0[60]}), .c ({y1_s2[60], y1_s1[60], y1_s0[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U728 ( .a ({temp_s2[61], temp_s1[61], temp_s0[61]}), .b ({temp_next_s2[61], temp_next_s1[61], temp_next_s0[61]}), .c ({y1_s2[61], y1_s1[61], y1_s0[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U729 ( .a ({temp_s2[62], temp_s1[62], temp_s0[62]}), .b ({temp_next_s2[62], temp_next_s1[62], temp_next_s0[62]}), .c ({y1_s2[62], y1_s1[62], y1_s0[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U730 ( .a ({temp_s2[63], temp_s1[63], temp_s0[63]}), .b ({temp_next_s2[63], temp_next_s1[63], temp_next_s0[63]}), .c ({y1_s2[63], y1_s1[63], y1_s0[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U731 ( .a ({temp_s2[64], temp_s1[64], temp_s0[64]}), .b ({temp_next_s2[64], temp_next_s1[64], temp_next_s0[64]}), .c ({y1_s2[64], y1_s1[64], y1_s0[64]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U732 ( .a ({temp_s2[65], temp_s1[65], temp_s0[65]}), .b ({temp_next_s2[65], temp_next_s1[65], temp_next_s0[65]}), .c ({y1_s2[65], y1_s1[65], y1_s0[65]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U733 ( .a ({temp_s2[66], temp_s1[66], temp_s0[66]}), .b ({temp_next_s2[66], temp_next_s1[66], temp_next_s0[66]}), .c ({y1_s2[66], y1_s1[66], y1_s0[66]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U734 ( .a ({temp_s2[67], temp_s1[67], temp_s0[67]}), .b ({temp_next_s2[67], temp_next_s1[67], temp_next_s0[67]}), .c ({y1_s2[67], y1_s1[67], y1_s0[67]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U735 ( .a ({temp_s2[68], temp_s1[68], temp_s0[68]}), .b ({temp_next_s2[68], temp_next_s1[68], temp_next_s0[68]}), .c ({y1_s2[68], y1_s1[68], y1_s0[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U736 ( .a ({temp_s2[69], temp_s1[69], temp_s0[69]}), .b ({temp_next_s2[69], temp_next_s1[69], temp_next_s0[69]}), .c ({y1_s2[69], y1_s1[69], y1_s0[69]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U737 ( .a ({temp_s2[6], temp_s1[6], temp_s0[6]}), .b ({temp_next_s2[6], temp_next_s1[6], temp_next_s0[6]}), .c ({y1_s2[6], y1_s1[6], y1_s0[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U738 ( .a ({temp_s2[70], temp_s1[70], temp_s0[70]}), .b ({temp_next_s2[70], temp_next_s1[70], temp_next_s0[70]}), .c ({y1_s2[70], y1_s1[70], y1_s0[70]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U739 ( .a ({temp_s2[71], temp_s1[71], temp_s0[71]}), .b ({temp_next_s2[71], temp_next_s1[71], temp_next_s0[71]}), .c ({y1_s2[71], y1_s1[71], y1_s0[71]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U740 ( .a ({temp_s2[72], temp_s1[72], temp_s0[72]}), .b ({temp_next_s2[72], temp_next_s1[72], temp_next_s0[72]}), .c ({y1_s2[72], y1_s1[72], y1_s0[72]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U741 ( .a ({temp_s2[73], temp_s1[73], temp_s0[73]}), .b ({temp_next_s2[73], temp_next_s1[73], temp_next_s0[73]}), .c ({y1_s2[73], y1_s1[73], y1_s0[73]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U742 ( .a ({temp_s2[74], temp_s1[74], temp_s0[74]}), .b ({temp_next_s2[74], temp_next_s1[74], temp_next_s0[74]}), .c ({y1_s2[74], y1_s1[74], y1_s0[74]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U743 ( .a ({temp_s2[75], temp_s1[75], temp_s0[75]}), .b ({temp_next_s2[75], temp_next_s1[75], temp_next_s0[75]}), .c ({y1_s2[75], y1_s1[75], y1_s0[75]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U744 ( .a ({temp_s2[76], temp_s1[76], temp_s0[76]}), .b ({temp_next_s2[76], temp_next_s1[76], temp_next_s0[76]}), .c ({y1_s2[76], y1_s1[76], y1_s0[76]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U745 ( .a ({temp_s2[77], temp_s1[77], temp_s0[77]}), .b ({temp_next_s2[77], temp_next_s1[77], temp_next_s0[77]}), .c ({y1_s2[77], y1_s1[77], y1_s0[77]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U746 ( .a ({temp_s2[78], temp_s1[78], temp_s0[78]}), .b ({temp_next_s2[78], temp_next_s1[78], temp_next_s0[78]}), .c ({y1_s2[78], y1_s1[78], y1_s0[78]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U747 ( .a ({temp_s2[79], temp_s1[79], temp_s0[79]}), .b ({temp_next_s2[79], temp_next_s1[79], temp_next_s0[79]}), .c ({y1_s2[79], y1_s1[79], y1_s0[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U748 ( .a ({temp_s2[7], temp_s1[7], temp_s0[7]}), .b ({temp_next_s2[7], temp_next_s1[7], temp_next_s0[7]}), .c ({y1_s2[7], y1_s1[7], y1_s0[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U749 ( .a ({temp_s2[80], temp_s1[80], temp_s0[80]}), .b ({temp_next_s2[80], temp_next_s1[80], temp_next_s0[80]}), .c ({y1_s2[80], y1_s1[80], y1_s0[80]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U750 ( .a ({temp_s2[81], temp_s1[81], temp_s0[81]}), .b ({temp_next_s2[81], temp_next_s1[81], temp_next_s0[81]}), .c ({y1_s2[81], y1_s1[81], y1_s0[81]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U751 ( .a ({temp_s2[82], temp_s1[82], temp_s0[82]}), .b ({temp_next_s2[82], temp_next_s1[82], temp_next_s0[82]}), .c ({y1_s2[82], y1_s1[82], y1_s0[82]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U752 ( .a ({temp_s2[83], temp_s1[83], temp_s0[83]}), .b ({temp_next_s2[83], temp_next_s1[83], temp_next_s0[83]}), .c ({y1_s2[83], y1_s1[83], y1_s0[83]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U753 ( .a ({temp_s2[84], temp_s1[84], temp_s0[84]}), .b ({temp_next_s2[84], temp_next_s1[84], temp_next_s0[84]}), .c ({y1_s2[84], y1_s1[84], y1_s0[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U754 ( .a ({temp_s2[85], temp_s1[85], temp_s0[85]}), .b ({temp_next_s2[85], temp_next_s1[85], temp_next_s0[85]}), .c ({y1_s2[85], y1_s1[85], y1_s0[85]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U755 ( .a ({temp_s2[86], temp_s1[86], temp_s0[86]}), .b ({temp_next_s2[86], temp_next_s1[86], temp_next_s0[86]}), .c ({y1_s2[86], y1_s1[86], y1_s0[86]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U756 ( .a ({temp_s2[87], temp_s1[87], temp_s0[87]}), .b ({temp_next_s2[87], temp_next_s1[87], temp_next_s0[87]}), .c ({y1_s2[87], y1_s1[87], y1_s0[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U757 ( .a ({temp_s2[88], temp_s1[88], temp_s0[88]}), .b ({temp_next_s2[88], temp_next_s1[88], temp_next_s0[88]}), .c ({y1_s2[88], y1_s1[88], y1_s0[88]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U758 ( .a ({temp_s2[89], temp_s1[89], temp_s0[89]}), .b ({temp_next_s2[89], temp_next_s1[89], temp_next_s0[89]}), .c ({y1_s2[89], y1_s1[89], y1_s0[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U759 ( .a ({temp_s2[8], temp_s1[8], temp_s0[8]}), .b ({temp_next_s2[8], temp_next_s1[8], temp_next_s0[8]}), .c ({y1_s2[8], y1_s1[8], y1_s0[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U760 ( .a ({temp_s2[90], temp_s1[90], temp_s0[90]}), .b ({temp_next_s2[90], temp_next_s1[90], temp_next_s0[90]}), .c ({y1_s2[90], y1_s1[90], y1_s0[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U761 ( .a ({temp_s2[91], temp_s1[91], temp_s0[91]}), .b ({temp_next_s2[91], temp_next_s1[91], temp_next_s0[91]}), .c ({y1_s2[91], y1_s1[91], y1_s0[91]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U762 ( .a ({temp_s2[92], temp_s1[92], temp_s0[92]}), .b ({temp_next_s2[92], temp_next_s1[92], temp_next_s0[92]}), .c ({y1_s2[92], y1_s1[92], y1_s0[92]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U763 ( .a ({temp_s2[93], temp_s1[93], temp_s0[93]}), .b ({temp_next_s2[93], temp_next_s1[93], temp_next_s0[93]}), .c ({y1_s2[93], y1_s1[93], y1_s0[93]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U764 ( .a ({temp_s2[94], temp_s1[94], temp_s0[94]}), .b ({temp_next_s2[94], temp_next_s1[94], temp_next_s0[94]}), .c ({y1_s2[94], y1_s1[94], y1_s0[94]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U765 ( .a ({temp_s2[95], temp_s1[95], temp_s0[95]}), .b ({temp_next_s2[95], temp_next_s1[95], temp_next_s0[95]}), .c ({y1_s2[95], y1_s1[95], y1_s0[95]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U766 ( .a ({temp_s2[96], temp_s1[96], temp_s0[96]}), .b ({temp_next_s2[96], temp_next_s1[96], temp_next_s0[96]}), .c ({y1_s2[96], y1_s1[96], y1_s0[96]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U767 ( .a ({temp_s2[97], temp_s1[97], temp_s0[97]}), .b ({temp_next_s2[97], temp_next_s1[97], temp_next_s0[97]}), .c ({y1_s2[97], y1_s1[97], y1_s0[97]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U768 ( .a ({temp_s2[98], temp_s1[98], temp_s0[98]}), .b ({temp_next_s2[98], temp_next_s1[98], temp_next_s0[98]}), .c ({y1_s2[98], y1_s1[98], y1_s0[98]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U769 ( .a ({temp_s2[99], temp_s1[99], temp_s0[99]}), .b ({temp_next_s2[99], temp_next_s1[99], temp_next_s0[99]}), .c ({y1_s2[99], y1_s1[99], y1_s0[99]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U770 ( .a ({temp_s2[9], temp_s1[9], temp_s0[9]}), .b ({temp_next_s2[9], temp_next_s1[9], temp_next_s0[9]}), .c ({y1_s2[9], y1_s1[9], y1_s0[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U96 ( .a ({new_AGEMA_signal_12997, new_AGEMA_signal_12996, mcs1_mcs_mat1_0_n128}), .b ({new_AGEMA_signal_13989, new_AGEMA_signal_13988, mcs1_mcs_mat1_0_n127}), .c ({temp_next_s2[93], temp_next_s1[93], temp_next_s0[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U95 ( .a ({new_AGEMA_signal_11515, new_AGEMA_signal_11514, mcs1_mcs_mat1_0_mcs_out[41]}), .b ({new_AGEMA_signal_13541, new_AGEMA_signal_13540, mcs1_mcs_mat1_0_mcs_out[45]}), .c ({new_AGEMA_signal_13989, new_AGEMA_signal_13988, mcs1_mcs_mat1_0_n127}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U94 ( .a ({new_AGEMA_signal_8765, new_AGEMA_signal_8764, mcs1_mcs_mat1_0_mcs_out[33]}), .b ({new_AGEMA_signal_12437, new_AGEMA_signal_12436, mcs1_mcs_mat1_0_mcs_out[37]}), .c ({new_AGEMA_signal_12997, new_AGEMA_signal_12996, mcs1_mcs_mat1_0_n128}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U93 ( .a ({new_AGEMA_signal_13505, new_AGEMA_signal_13504, mcs1_mcs_mat1_0_n126}), .b ({new_AGEMA_signal_15997, new_AGEMA_signal_15996, mcs1_mcs_mat1_0_n125}), .c ({temp_next_s2[92], temp_next_s1[92], temp_next_s0[92]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U92 ( .a ({new_AGEMA_signal_10547, new_AGEMA_signal_10546, mcs1_mcs_mat1_0_mcs_out[40]}), .b ({new_AGEMA_signal_15519, new_AGEMA_signal_15518, mcs1_mcs_mat1_0_mcs_out[44]}), .c ({new_AGEMA_signal_15997, new_AGEMA_signal_15996, mcs1_mcs_mat1_0_n125}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U91 ( .a ({new_AGEMA_signal_13051, new_AGEMA_signal_13050, mcs1_mcs_mat1_0_mcs_out[32]}), .b ({new_AGEMA_signal_10551, new_AGEMA_signal_10550, mcs1_mcs_mat1_0_mcs_out[36]}), .c ({new_AGEMA_signal_13505, new_AGEMA_signal_13504, mcs1_mcs_mat1_0_n126}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U90 ( .a ({new_AGEMA_signal_11429, new_AGEMA_signal_11428, mcs1_mcs_mat1_0_n124}), .b ({new_AGEMA_signal_15485, new_AGEMA_signal_15484, mcs1_mcs_mat1_0_n123}), .c ({temp_next_s2[63], temp_next_s1[63], temp_next_s0[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U89 ( .a ({new_AGEMA_signal_10559, new_AGEMA_signal_10558, mcs1_mcs_mat1_0_mcs_out[27]}), .b ({new_AGEMA_signal_14929, new_AGEMA_signal_14928, mcs1_mcs_mat1_0_mcs_out[31]}), .c ({new_AGEMA_signal_15485, new_AGEMA_signal_15484, mcs1_mcs_mat1_0_n123}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U88 ( .a ({new_AGEMA_signal_10571, new_AGEMA_signal_10570, mcs1_mcs_mat1_0_mcs_out[19]}), .b ({new_AGEMA_signal_10565, new_AGEMA_signal_10564, mcs1_mcs_mat1_0_mcs_out[23]}), .c ({new_AGEMA_signal_11429, new_AGEMA_signal_11428, mcs1_mcs_mat1_0_n124}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U87 ( .a ({new_AGEMA_signal_12389, new_AGEMA_signal_12388, mcs1_mcs_mat1_0_n122}), .b ({new_AGEMA_signal_14893, new_AGEMA_signal_14892, mcs1_mcs_mat1_0_n121}), .c ({temp_next_s2[62], temp_next_s1[62], temp_next_s0[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U86 ( .a ({new_AGEMA_signal_11525, new_AGEMA_signal_11524, mcs1_mcs_mat1_0_mcs_out[26]}), .b ({new_AGEMA_signal_14443, new_AGEMA_signal_14442, mcs1_mcs_mat1_0_mcs_out[30]}), .c ({new_AGEMA_signal_14893, new_AGEMA_signal_14892, mcs1_mcs_mat1_0_n121}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U85 ( .a ({new_AGEMA_signal_11533, new_AGEMA_signal_11532, mcs1_mcs_mat1_0_mcs_out[18]}), .b ({new_AGEMA_signal_11529, new_AGEMA_signal_11528, mcs1_mcs_mat1_0_mcs_out[22]}), .c ({new_AGEMA_signal_12389, new_AGEMA_signal_12388, mcs1_mcs_mat1_0_n122}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U84 ( .a ({new_AGEMA_signal_12999, new_AGEMA_signal_12998, mcs1_mcs_mat1_0_n120}), .b ({new_AGEMA_signal_14411, new_AGEMA_signal_14410, mcs1_mcs_mat1_0_n119}), .c ({temp_next_s2[61], temp_next_s1[61], temp_next_s0[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U83 ( .a ({new_AGEMA_signal_12441, new_AGEMA_signal_12440, mcs1_mcs_mat1_0_mcs_out[25]}), .b ({new_AGEMA_signal_14023, new_AGEMA_signal_14022, mcs1_mcs_mat1_0_mcs_out[29]}), .c ({new_AGEMA_signal_14411, new_AGEMA_signal_14410, mcs1_mcs_mat1_0_n119}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U82 ( .a ({new_AGEMA_signal_12445, new_AGEMA_signal_12444, mcs1_mcs_mat1_0_mcs_out[17]}), .b ({new_AGEMA_signal_12443, new_AGEMA_signal_12442, mcs1_mcs_mat1_0_mcs_out[21]}), .c ({new_AGEMA_signal_12999, new_AGEMA_signal_12998, mcs1_mcs_mat1_0_n120}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U81 ( .a ({new_AGEMA_signal_11431, new_AGEMA_signal_11430, mcs1_mcs_mat1_0_n118}), .b ({new_AGEMA_signal_15489, new_AGEMA_signal_15488, mcs1_mcs_mat1_0_n117}), .c ({temp_next_s2[60], temp_next_s1[60], temp_next_s0[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U80 ( .a ({new_AGEMA_signal_10563, new_AGEMA_signal_10562, mcs1_mcs_mat1_0_mcs_out[24]}), .b ({new_AGEMA_signal_14931, new_AGEMA_signal_14930, mcs1_mcs_mat1_0_mcs_out[28]}), .c ({new_AGEMA_signal_15489, new_AGEMA_signal_15488, mcs1_mcs_mat1_0_n117}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U79 ( .a ({new_AGEMA_signal_10575, new_AGEMA_signal_10574, mcs1_mcs_mat1_0_mcs_out[16]}), .b ({new_AGEMA_signal_10569, new_AGEMA_signal_10568, mcs1_mcs_mat1_0_mcs_out[20]}), .c ({new_AGEMA_signal_11431, new_AGEMA_signal_11430, mcs1_mcs_mat1_0_n118}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U78 ( .a ({new_AGEMA_signal_15491, new_AGEMA_signal_15490, mcs1_mcs_mat1_0_n116}), .b ({new_AGEMA_signal_13001, new_AGEMA_signal_13000, mcs1_mcs_mat1_0_n115}), .c ({temp_next_s2[31], temp_next_s1[31], temp_next_s0[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U77 ( .a ({new_AGEMA_signal_10585, new_AGEMA_signal_10584, mcs1_mcs_mat1_0_mcs_out[3]}), .b ({new_AGEMA_signal_12451, new_AGEMA_signal_12450, mcs1_mcs_mat1_0_mcs_out[7]}), .c ({new_AGEMA_signal_13001, new_AGEMA_signal_13000, mcs1_mcs_mat1_0_n115}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U76 ( .a ({new_AGEMA_signal_8957, new_AGEMA_signal_8956, mcs1_mcs_mat1_0_mcs_out[11]}), .b ({new_AGEMA_signal_14933, new_AGEMA_signal_14932, mcs1_mcs_mat1_0_mcs_out[15]}), .c ({new_AGEMA_signal_15491, new_AGEMA_signal_15490, mcs1_mcs_mat1_0_n116}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U75 ( .a ({new_AGEMA_signal_13005, new_AGEMA_signal_13004, mcs1_mcs_mat1_0_n114}), .b ({new_AGEMA_signal_13003, new_AGEMA_signal_13002, mcs1_mcs_mat1_0_n113}), .c ({new_AGEMA_signal_13507, new_AGEMA_signal_13506, mcs_out[255]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U74 ( .a ({new_AGEMA_signal_12405, new_AGEMA_signal_12404, mcs1_mcs_mat1_0_mcs_out[123]}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_13003, new_AGEMA_signal_13002, mcs1_mcs_mat1_0_n113}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U73 ( .a ({new_AGEMA_signal_11457, new_AGEMA_signal_11456, mcs1_mcs_mat1_0_mcs_out[115]}), .b ({new_AGEMA_signal_12409, new_AGEMA_signal_12408, mcs1_mcs_mat1_0_mcs_out[119]}), .c ({new_AGEMA_signal_13005, new_AGEMA_signal_13004, mcs1_mcs_mat1_0_n114}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U72 ( .a ({new_AGEMA_signal_13007, new_AGEMA_signal_13006, mcs1_mcs_mat1_0_n112}), .b ({new_AGEMA_signal_13509, new_AGEMA_signal_13508, mcs1_mcs_mat1_0_n111}), .c ({new_AGEMA_signal_13991, new_AGEMA_signal_13990, mcs_out[254]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U71 ( .a ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, mcs1_mcs_mat1_0_mcs_out[122]}), .b ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_13509, new_AGEMA_signal_13508, mcs1_mcs_mat1_0_n111}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U70 ( .a ({new_AGEMA_signal_10481, new_AGEMA_signal_10480, mcs1_mcs_mat1_0_mcs_out[114]}), .b ({new_AGEMA_signal_12411, new_AGEMA_signal_12410, mcs1_mcs_mat1_0_mcs_out[118]}), .c ({new_AGEMA_signal_13007, new_AGEMA_signal_13006, mcs1_mcs_mat1_0_n112}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U69 ( .a ({new_AGEMA_signal_14897, new_AGEMA_signal_14896, mcs1_mcs_mat1_0_n110}), .b ({new_AGEMA_signal_11433, new_AGEMA_signal_11432, mcs1_mcs_mat1_0_n109}), .c ({temp_next_s2[30], temp_next_s1[30], temp_next_s0[30]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U68 ( .a ({new_AGEMA_signal_10587, new_AGEMA_signal_10586, mcs1_mcs_mat1_0_mcs_out[2]}), .b ({new_AGEMA_signal_10583, new_AGEMA_signal_10582, mcs1_mcs_mat1_0_mcs_out[6]}), .c ({new_AGEMA_signal_11433, new_AGEMA_signal_11432, mcs1_mcs_mat1_0_n109}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U67 ( .a ({new_AGEMA_signal_11539, new_AGEMA_signal_11538, mcs1_mcs_mat1_0_mcs_out[10]}), .b ({new_AGEMA_signal_14447, new_AGEMA_signal_14446, mcs1_mcs_mat1_0_mcs_out[14]}), .c ({new_AGEMA_signal_14897, new_AGEMA_signal_14896, mcs1_mcs_mat1_0_n110}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U66 ( .a ({new_AGEMA_signal_12391, new_AGEMA_signal_12390, mcs1_mcs_mat1_0_n108}), .b ({new_AGEMA_signal_13511, new_AGEMA_signal_13510, mcs1_mcs_mat1_0_n107}), .c ({new_AGEMA_signal_13993, new_AGEMA_signal_13992, mcs_out[253]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U65 ( .a ({new_AGEMA_signal_12407, new_AGEMA_signal_12406, mcs1_mcs_mat1_0_mcs_out[121]}), .b ({new_AGEMA_signal_13029, new_AGEMA_signal_13028, mcs1_mcs_mat1_0_mcs_out[125]}), .c ({new_AGEMA_signal_13511, new_AGEMA_signal_13510, mcs1_mcs_mat1_0_n107}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U64 ( .a ({new_AGEMA_signal_9523, new_AGEMA_signal_9522, mcs1_mcs_mat1_0_mcs_out[113]}), .b ({new_AGEMA_signal_11455, new_AGEMA_signal_11454, mcs1_mcs_mat1_0_mcs_out[117]}), .c ({new_AGEMA_signal_12391, new_AGEMA_signal_12390, mcs1_mcs_mat1_0_n108}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U63 ( .a ({new_AGEMA_signal_13011, new_AGEMA_signal_13010, mcs1_mcs_mat1_0_n106}), .b ({new_AGEMA_signal_13009, new_AGEMA_signal_13008, mcs1_mcs_mat1_0_n105}), .c ({new_AGEMA_signal_13513, new_AGEMA_signal_13512, mcs_out[252]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U62 ( .a ({new_AGEMA_signal_11449, new_AGEMA_signal_11448, mcs1_mcs_mat1_0_mcs_out[120]}), .b ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_13009, new_AGEMA_signal_13008, mcs1_mcs_mat1_0_n105}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U61 ( .a ({new_AGEMA_signal_12413, new_AGEMA_signal_12412, mcs1_mcs_mat1_0_mcs_out[112]}), .b ({new_AGEMA_signal_10479, new_AGEMA_signal_10478, mcs1_mcs_mat1_0_mcs_out[116]}), .c ({new_AGEMA_signal_13011, new_AGEMA_signal_13010, mcs1_mcs_mat1_0_n106}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U60 ( .a ({new_AGEMA_signal_12393, new_AGEMA_signal_12392, mcs1_mcs_mat1_0_n104}), .b ({new_AGEMA_signal_15495, new_AGEMA_signal_15494, mcs1_mcs_mat1_0_n103}), .c ({new_AGEMA_signal_16005, new_AGEMA_signal_16004, mcs_out[223]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U59 ( .a ({new_AGEMA_signal_14913, new_AGEMA_signal_14912, mcs1_mcs_mat1_0_mcs_out[111]}), .b ({new_AGEMA_signal_12417, new_AGEMA_signal_12416, mcs1_mcs_mat1_0_mcs_out[99]}), .c ({new_AGEMA_signal_15495, new_AGEMA_signal_15494, mcs1_mcs_mat1_0_n103}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U58 ( .a ({new_AGEMA_signal_11471, new_AGEMA_signal_11470, mcs1_mcs_mat1_0_mcs_out[103]}), .b ({new_AGEMA_signal_11463, new_AGEMA_signal_11462, mcs1_mcs_mat1_0_mcs_out[107]}), .c ({new_AGEMA_signal_12393, new_AGEMA_signal_12392, mcs1_mcs_mat1_0_n104}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U57 ( .a ({new_AGEMA_signal_12395, new_AGEMA_signal_12394, mcs1_mcs_mat1_0_n102}), .b ({new_AGEMA_signal_15497, new_AGEMA_signal_15496, mcs1_mcs_mat1_0_n101}), .c ({new_AGEMA_signal_16007, new_AGEMA_signal_16006, mcs_out[222]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U56 ( .a ({new_AGEMA_signal_14915, new_AGEMA_signal_14914, mcs1_mcs_mat1_0_mcs_out[110]}), .b ({new_AGEMA_signal_10499, new_AGEMA_signal_10498, mcs1_mcs_mat1_0_mcs_out[98]}), .c ({new_AGEMA_signal_15497, new_AGEMA_signal_15496, mcs1_mcs_mat1_0_n101}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U55 ( .a ({new_AGEMA_signal_9533, new_AGEMA_signal_9532, mcs1_mcs_mat1_0_mcs_out[102]}), .b ({new_AGEMA_signal_11465, new_AGEMA_signal_11464, mcs1_mcs_mat1_0_mcs_out[106]}), .c ({new_AGEMA_signal_12395, new_AGEMA_signal_12394, mcs1_mcs_mat1_0_n102}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U54 ( .a ({new_AGEMA_signal_12397, new_AGEMA_signal_12396, mcs1_mcs_mat1_0_n100}), .b ({new_AGEMA_signal_15499, new_AGEMA_signal_15498, mcs1_mcs_mat1_0_n99}), .c ({new_AGEMA_signal_16009, new_AGEMA_signal_16008, mcs_out[221]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U53 ( .a ({new_AGEMA_signal_14917, new_AGEMA_signal_14916, mcs1_mcs_mat1_0_mcs_out[109]}), .b ({new_AGEMA_signal_8915, new_AGEMA_signal_8914, mcs1_mcs_mat1_0_mcs_out[97]}), .c ({new_AGEMA_signal_15499, new_AGEMA_signal_15498, mcs1_mcs_mat1_0_n99}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U52 ( .a ({new_AGEMA_signal_10495, new_AGEMA_signal_10494, mcs1_mcs_mat1_0_mcs_out[101]}), .b ({new_AGEMA_signal_11467, new_AGEMA_signal_11466, mcs1_mcs_mat1_0_mcs_out[105]}), .c ({new_AGEMA_signal_12397, new_AGEMA_signal_12396, mcs1_mcs_mat1_0_n100}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U51 ( .a ({new_AGEMA_signal_13013, new_AGEMA_signal_13012, mcs1_mcs_mat1_0_n98}), .b ({new_AGEMA_signal_15501, new_AGEMA_signal_15500, mcs1_mcs_mat1_0_n97}), .c ({new_AGEMA_signal_16011, new_AGEMA_signal_16010, mcs_out[220]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U50 ( .a ({new_AGEMA_signal_14919, new_AGEMA_signal_14918, mcs1_mcs_mat1_0_mcs_out[108]}), .b ({new_AGEMA_signal_13525, new_AGEMA_signal_13524, mcs1_mcs_mat1_0_mcs_out[96]}), .c ({new_AGEMA_signal_15501, new_AGEMA_signal_15500, mcs1_mcs_mat1_0_n97}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U49 ( .a ({new_AGEMA_signal_11473, new_AGEMA_signal_11472, mcs1_mcs_mat1_0_mcs_out[100]}), .b ({new_AGEMA_signal_12415, new_AGEMA_signal_12414, mcs1_mcs_mat1_0_mcs_out[104]}), .c ({new_AGEMA_signal_13013, new_AGEMA_signal_13012, mcs1_mcs_mat1_0_n98}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U48 ( .a ({new_AGEMA_signal_11435, new_AGEMA_signal_11434, mcs1_mcs_mat1_0_n96}), .b ({new_AGEMA_signal_14899, new_AGEMA_signal_14898, mcs1_mcs_mat1_0_n95}), .c ({new_AGEMA_signal_15503, new_AGEMA_signal_15502, mcs_out[191]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U47 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_14427, new_AGEMA_signal_14426, mcs1_mcs_mat1_0_mcs_out[95]}), .c ({new_AGEMA_signal_14899, new_AGEMA_signal_14898, mcs1_mcs_mat1_0_n95}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U46 ( .a ({new_AGEMA_signal_10505, new_AGEMA_signal_10504, mcs1_mcs_mat1_0_mcs_out[83]}), .b ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, mcs1_mcs_mat1_0_mcs_out[87]}), .c ({new_AGEMA_signal_11435, new_AGEMA_signal_11434, mcs1_mcs_mat1_0_n96}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U45 ( .a ({new_AGEMA_signal_11437, new_AGEMA_signal_11436, mcs1_mcs_mat1_0_n94}), .b ({new_AGEMA_signal_13995, new_AGEMA_signal_13994, mcs1_mcs_mat1_0_n93}), .c ({new_AGEMA_signal_14413, new_AGEMA_signal_14412, mcs_out[190]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U43 ( .a ({new_AGEMA_signal_10507, new_AGEMA_signal_10506, mcs1_mcs_mat1_0_mcs_out[82]}), .b ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_11437, new_AGEMA_signal_11436, mcs1_mcs_mat1_0_n94}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U42 ( .a ({new_AGEMA_signal_11439, new_AGEMA_signal_11438, mcs1_mcs_mat1_0_n92}), .b ({new_AGEMA_signal_13997, new_AGEMA_signal_13996, mcs1_mcs_mat1_0_n91}), .c ({new_AGEMA_signal_14415, new_AGEMA_signal_14414, mcs_out[189]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U41 ( .a ({new_AGEMA_signal_8921, new_AGEMA_signal_8920, mcs1_mcs_mat1_0_mcs_out[89]}), .b ({new_AGEMA_signal_13529, new_AGEMA_signal_13528, mcs1_mcs_mat1_0_mcs_out[93]}), .c ({new_AGEMA_signal_13997, new_AGEMA_signal_13996, mcs1_mcs_mat1_0_n91}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U40 ( .a ({new_AGEMA_signal_10509, new_AGEMA_signal_10508, mcs1_mcs_mat1_0_mcs_out[81]}), .b ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_11439, new_AGEMA_signal_11438, mcs1_mcs_mat1_0_n92}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U39 ( .a ({new_AGEMA_signal_12399, new_AGEMA_signal_12398, mcs1_mcs_mat1_0_n90}), .b ({new_AGEMA_signal_15505, new_AGEMA_signal_15504, mcs1_mcs_mat1_0_n89}), .c ({new_AGEMA_signal_16013, new_AGEMA_signal_16012, mcs_out[188]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U38 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_14921, new_AGEMA_signal_14920, mcs1_mcs_mat1_0_mcs_out[92]}), .c ({new_AGEMA_signal_15505, new_AGEMA_signal_15504, mcs1_mcs_mat1_0_n89}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U37 ( .a ({new_AGEMA_signal_11479, new_AGEMA_signal_11478, mcs1_mcs_mat1_0_mcs_out[80]}), .b ({new_AGEMA_signal_10503, new_AGEMA_signal_10502, mcs1_mcs_mat1_0_mcs_out[84]}), .c ({new_AGEMA_signal_12399, new_AGEMA_signal_12398, mcs1_mcs_mat1_0_n90}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U36 ( .a ({new_AGEMA_signal_14901, new_AGEMA_signal_14900, mcs1_mcs_mat1_0_n88}), .b ({new_AGEMA_signal_11441, new_AGEMA_signal_11440, mcs1_mcs_mat1_0_n87}), .c ({temp_next_s2[29], temp_next_s1[29], temp_next_s0[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U35 ( .a ({new_AGEMA_signal_8961, new_AGEMA_signal_8960, mcs1_mcs_mat1_0_mcs_out[5]}), .b ({new_AGEMA_signal_10579, new_AGEMA_signal_10578, mcs1_mcs_mat1_0_mcs_out[9]}), .c ({new_AGEMA_signal_11441, new_AGEMA_signal_11440, mcs1_mcs_mat1_0_n87}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U34 ( .a ({new_AGEMA_signal_14449, new_AGEMA_signal_14448, mcs1_mcs_mat1_0_mcs_out[13]}), .b ({new_AGEMA_signal_11545, new_AGEMA_signal_11544, mcs1_mcs_mat1_0_mcs_out[1]}), .c ({new_AGEMA_signal_14901, new_AGEMA_signal_14900, mcs1_mcs_mat1_0_n88}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U33 ( .a ({new_AGEMA_signal_13015, new_AGEMA_signal_13014, mcs1_mcs_mat1_0_n86}), .b ({new_AGEMA_signal_14903, new_AGEMA_signal_14902, mcs1_mcs_mat1_0_n85}), .c ({new_AGEMA_signal_15509, new_AGEMA_signal_15508, mcs_out[159]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U32 ( .a ({new_AGEMA_signal_9553, new_AGEMA_signal_9552, mcs1_mcs_mat1_0_mcs_out[75]}), .b ({new_AGEMA_signal_14431, new_AGEMA_signal_14430, mcs1_mcs_mat1_0_mcs_out[79]}), .c ({new_AGEMA_signal_14903, new_AGEMA_signal_14902, mcs1_mcs_mat1_0_n85}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U31 ( .a ({new_AGEMA_signal_12427, new_AGEMA_signal_12426, mcs1_mcs_mat1_0_mcs_out[67]}), .b ({new_AGEMA_signal_11489, new_AGEMA_signal_11488, mcs1_mcs_mat1_0_mcs_out[71]}), .c ({new_AGEMA_signal_13015, new_AGEMA_signal_13014, mcs1_mcs_mat1_0_n86}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U30 ( .a ({new_AGEMA_signal_13019, new_AGEMA_signal_13018, mcs1_mcs_mat1_0_n84}), .b ({new_AGEMA_signal_13017, new_AGEMA_signal_13016, mcs1_mcs_mat1_0_n83}), .c ({new_AGEMA_signal_13515, new_AGEMA_signal_13514, mcs_out[158]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U29 ( .a ({new_AGEMA_signal_12419, new_AGEMA_signal_12418, mcs1_mcs_mat1_0_mcs_out[74]}), .b ({new_AGEMA_signal_11481, new_AGEMA_signal_11480, mcs1_mcs_mat1_0_mcs_out[78]}), .c ({new_AGEMA_signal_13017, new_AGEMA_signal_13016, mcs1_mcs_mat1_0_n83}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U28 ( .a ({new_AGEMA_signal_11495, new_AGEMA_signal_11494, mcs1_mcs_mat1_0_mcs_out[66]}), .b ({new_AGEMA_signal_12423, new_AGEMA_signal_12422, mcs1_mcs_mat1_0_mcs_out[70]}), .c ({new_AGEMA_signal_13019, new_AGEMA_signal_13018, mcs1_mcs_mat1_0_n84}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U27 ( .a ({new_AGEMA_signal_13021, new_AGEMA_signal_13020, mcs1_mcs_mat1_0_n82}), .b ({new_AGEMA_signal_13999, new_AGEMA_signal_13998, mcs1_mcs_mat1_0_n81}), .c ({new_AGEMA_signal_14417, new_AGEMA_signal_14416, mcs_out[157]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U26 ( .a ({new_AGEMA_signal_10515, new_AGEMA_signal_10514, mcs1_mcs_mat1_0_mcs_out[73]}), .b ({new_AGEMA_signal_13533, new_AGEMA_signal_13532, mcs1_mcs_mat1_0_mcs_out[77]}), .c ({new_AGEMA_signal_13999, new_AGEMA_signal_13998, mcs1_mcs_mat1_0_n81}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U25 ( .a ({new_AGEMA_signal_9565, new_AGEMA_signal_9564, mcs1_mcs_mat1_0_mcs_out[65]}), .b ({new_AGEMA_signal_12425, new_AGEMA_signal_12424, mcs1_mcs_mat1_0_mcs_out[69]}), .c ({new_AGEMA_signal_13021, new_AGEMA_signal_13020, mcs1_mcs_mat1_0_n82}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U24 ( .a ({new_AGEMA_signal_13517, new_AGEMA_signal_13516, mcs1_mcs_mat1_0_n80}), .b ({new_AGEMA_signal_15511, new_AGEMA_signal_15510, mcs1_mcs_mat1_0_n79}), .c ({new_AGEMA_signal_16015, new_AGEMA_signal_16014, mcs_out[156]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U23 ( .a ({new_AGEMA_signal_12421, new_AGEMA_signal_12420, mcs1_mcs_mat1_0_mcs_out[72]}), .b ({new_AGEMA_signal_14923, new_AGEMA_signal_14922, mcs1_mcs_mat1_0_mcs_out[76]}), .c ({new_AGEMA_signal_15511, new_AGEMA_signal_15510, mcs1_mcs_mat1_0_n79}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U22 ( .a ({new_AGEMA_signal_13043, new_AGEMA_signal_13042, mcs1_mcs_mat1_0_mcs_out[64]}), .b ({new_AGEMA_signal_11493, new_AGEMA_signal_11492, mcs1_mcs_mat1_0_mcs_out[68]}), .c ({new_AGEMA_signal_13517, new_AGEMA_signal_13516, mcs1_mcs_mat1_0_n80}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U21 ( .a ({new_AGEMA_signal_12401, new_AGEMA_signal_12400, mcs1_mcs_mat1_0_n78}), .b ({new_AGEMA_signal_14905, new_AGEMA_signal_14904, mcs1_mcs_mat1_0_n77}), .c ({temp_next_s2[127], temp_next_s1[127], temp_next_s0[127]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U20 ( .a ({new_AGEMA_signal_10527, new_AGEMA_signal_10526, mcs1_mcs_mat1_0_mcs_out[59]}), .b ({new_AGEMA_signal_14435, new_AGEMA_signal_14434, mcs1_mcs_mat1_0_mcs_out[63]}), .c ({new_AGEMA_signal_14905, new_AGEMA_signal_14904, mcs1_mcs_mat1_0_n77}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U19 ( .a ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, mcs1_mcs_mat1_0_mcs_out[51]}), .b ({new_AGEMA_signal_11503, new_AGEMA_signal_11502, mcs1_mcs_mat1_0_mcs_out[55]}), .c ({new_AGEMA_signal_12401, new_AGEMA_signal_12400, mcs1_mcs_mat1_0_n78}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U18 ( .a ({new_AGEMA_signal_13023, new_AGEMA_signal_13022, mcs1_mcs_mat1_0_n76}), .b ({new_AGEMA_signal_14419, new_AGEMA_signal_14418, mcs1_mcs_mat1_0_n75}), .c ({temp_next_s2[126], temp_next_s1[126], temp_next_s0[126]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U17 ( .a ({new_AGEMA_signal_9569, new_AGEMA_signal_9568, mcs1_mcs_mat1_0_mcs_out[58]}), .b ({new_AGEMA_signal_14013, new_AGEMA_signal_14012, mcs1_mcs_mat1_0_mcs_out[62]}), .c ({new_AGEMA_signal_14419, new_AGEMA_signal_14418, mcs1_mcs_mat1_0_n75}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U16 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_12431, new_AGEMA_signal_12430, mcs1_mcs_mat1_0_mcs_out[54]}), .c ({new_AGEMA_signal_13023, new_AGEMA_signal_13022, mcs1_mcs_mat1_0_n76}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U15 ( .a ({new_AGEMA_signal_13025, new_AGEMA_signal_13024, mcs1_mcs_mat1_0_n74}), .b ({new_AGEMA_signal_14421, new_AGEMA_signal_14420, mcs1_mcs_mat1_0_n73}), .c ({temp_next_s2[125], temp_next_s1[125], temp_next_s0[125]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U14 ( .a ({new_AGEMA_signal_10529, new_AGEMA_signal_10528, mcs1_mcs_mat1_0_mcs_out[57]}), .b ({new_AGEMA_signal_14015, new_AGEMA_signal_14014, mcs1_mcs_mat1_0_mcs_out[61]}), .c ({new_AGEMA_signal_14421, new_AGEMA_signal_14420, mcs1_mcs_mat1_0_n73}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U13 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_12433, new_AGEMA_signal_12432, mcs1_mcs_mat1_0_mcs_out[53]}), .c ({new_AGEMA_signal_13025, new_AGEMA_signal_13024, mcs1_mcs_mat1_0_n74}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U12 ( .a ({new_AGEMA_signal_12403, new_AGEMA_signal_12402, mcs1_mcs_mat1_0_n72}), .b ({new_AGEMA_signal_15515, new_AGEMA_signal_15514, mcs1_mcs_mat1_0_n71}), .c ({temp_next_s2[124], temp_next_s1[124], temp_next_s0[124]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U11 ( .a ({new_AGEMA_signal_11501, new_AGEMA_signal_11500, mcs1_mcs_mat1_0_mcs_out[56]}), .b ({new_AGEMA_signal_14925, new_AGEMA_signal_14924, mcs1_mcs_mat1_0_mcs_out[60]}), .c ({new_AGEMA_signal_15515, new_AGEMA_signal_15514, mcs1_mcs_mat1_0_n71}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U10 ( .a ({new_AGEMA_signal_10537, new_AGEMA_signal_10536, mcs1_mcs_mat1_0_mcs_out[48]}), .b ({new_AGEMA_signal_11507, new_AGEMA_signal_11506, mcs1_mcs_mat1_0_mcs_out[52]}), .c ({new_AGEMA_signal_12403, new_AGEMA_signal_12402, mcs1_mcs_mat1_0_n72}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U9 ( .a ({new_AGEMA_signal_13027, new_AGEMA_signal_13026, mcs1_mcs_mat1_0_n70}), .b ({new_AGEMA_signal_14911, new_AGEMA_signal_14910, mcs1_mcs_mat1_0_n69}), .c ({temp_next_s2[95], temp_next_s1[95], temp_next_s0[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U8 ( .a ({new_AGEMA_signal_11511, new_AGEMA_signal_11510, mcs1_mcs_mat1_0_mcs_out[43]}), .b ({new_AGEMA_signal_14439, new_AGEMA_signal_14438, mcs1_mcs_mat1_0_mcs_out[47]}), .c ({new_AGEMA_signal_14911, new_AGEMA_signal_14910, mcs1_mcs_mat1_0_n69}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U7 ( .a ({new_AGEMA_signal_11519, new_AGEMA_signal_11518, mcs1_mcs_mat1_0_mcs_out[35]}), .b ({new_AGEMA_signal_12435, new_AGEMA_signal_12434, mcs1_mcs_mat1_0_mcs_out[39]}), .c ({new_AGEMA_signal_13027, new_AGEMA_signal_13026, mcs1_mcs_mat1_0_n70}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U6 ( .a ({new_AGEMA_signal_11443, new_AGEMA_signal_11442, mcs1_mcs_mat1_0_n68}), .b ({new_AGEMA_signal_13519, new_AGEMA_signal_13518, mcs1_mcs_mat1_0_n67}), .c ({temp_next_s2[94], temp_next_s1[94], temp_next_s0[94]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U5 ( .a ({new_AGEMA_signal_11513, new_AGEMA_signal_11512, mcs1_mcs_mat1_0_mcs_out[42]}), .b ({new_AGEMA_signal_13047, new_AGEMA_signal_13046, mcs1_mcs_mat1_0_mcs_out[46]}), .c ({new_AGEMA_signal_13519, new_AGEMA_signal_13518, mcs1_mcs_mat1_0_n67}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U4 ( .a ({new_AGEMA_signal_10553, new_AGEMA_signal_10552, mcs1_mcs_mat1_0_mcs_out[34]}), .b ({new_AGEMA_signal_9593, new_AGEMA_signal_9592, mcs1_mcs_mat1_0_mcs_out[38]}), .c ({new_AGEMA_signal_11443, new_AGEMA_signal_11442, mcs1_mcs_mat1_0_n68}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U3 ( .a ({new_AGEMA_signal_16019, new_AGEMA_signal_16018, mcs1_mcs_mat1_0_n66}), .b ({new_AGEMA_signal_14003, new_AGEMA_signal_14002, mcs1_mcs_mat1_0_n65}), .c ({temp_next_s2[28], temp_next_s1[28], temp_next_s0[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U2 ( .a ({new_AGEMA_signal_13555, new_AGEMA_signal_13554, mcs1_mcs_mat1_0_mcs_out[4]}), .b ({new_AGEMA_signal_12449, new_AGEMA_signal_12448, mcs1_mcs_mat1_0_mcs_out[8]}), .c ({new_AGEMA_signal_14003, new_AGEMA_signal_14002, mcs1_mcs_mat1_0_n65}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_U1 ( .a ({new_AGEMA_signal_11547, new_AGEMA_signal_11546, mcs1_mcs_mat1_0_mcs_out[0]}), .b ({new_AGEMA_signal_15521, new_AGEMA_signal_15520, mcs1_mcs_mat1_0_mcs_out[12]}), .c ({new_AGEMA_signal_16019, new_AGEMA_signal_16018, mcs1_mcs_mat1_0_n66}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_11445, new_AGEMA_signal_11444, mcs1_mcs_mat1_0_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_12405, new_AGEMA_signal_12404, mcs1_mcs_mat1_0_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_10473, new_AGEMA_signal_10472, mcs1_mcs_mat1_0_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_7669, new_AGEMA_signal_7668, mcs1_mcs_mat1_0_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_11445, new_AGEMA_signal_11444, mcs1_mcs_mat1_0_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_8173, new_AGEMA_signal_8172, mcs1_mcs_mat1_0_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_8893, new_AGEMA_signal_8892, mcs1_mcs_mat1_0_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, mcs1_mcs_mat1_0_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_8175, new_AGEMA_signal_8174, mcs1_mcs_mat1_0_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .c ({new_AGEMA_signal_8893, new_AGEMA_signal_8892, mcs1_mcs_mat1_0_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_11447, new_AGEMA_signal_11446, mcs1_mcs_mat1_0_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .c ({new_AGEMA_signal_12407, new_AGEMA_signal_12406, mcs1_mcs_mat1_0_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_10473, new_AGEMA_signal_10472, mcs1_mcs_mat1_0_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_11447, new_AGEMA_signal_11446, mcs1_mcs_mat1_0_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_9515, new_AGEMA_signal_9514, mcs1_mcs_mat1_0_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_8895, new_AGEMA_signal_8894, mcs1_mcs_mat1_0_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_10473, new_AGEMA_signal_10472, mcs1_mcs_mat1_0_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_10475, new_AGEMA_signal_10474, mcs1_mcs_mat1_0_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_11449, new_AGEMA_signal_11448, mcs1_mcs_mat1_0_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_9515, new_AGEMA_signal_9514, mcs1_mcs_mat1_0_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_8175, new_AGEMA_signal_8174, mcs1_mcs_mat1_0_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_10475, new_AGEMA_signal_10474, mcs1_mcs_mat1_0_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_9515, new_AGEMA_signal_9514, mcs1_mcs_mat1_0_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347]}), .c ({new_AGEMA_signal_8175, new_AGEMA_signal_8174, mcs1_mcs_mat1_0_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_8895, new_AGEMA_signal_8894, mcs1_mcs_mat1_0_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_11451, new_AGEMA_signal_11450, mcs1_mcs_mat1_0_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .c ({new_AGEMA_signal_12409, new_AGEMA_signal_12408, mcs1_mcs_mat1_0_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_10477, new_AGEMA_signal_10476, mcs1_mcs_mat1_0_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_8901, new_AGEMA_signal_8900, mcs1_mcs_mat1_0_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_11451, new_AGEMA_signal_11450, mcs1_mcs_mat1_0_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_11453, new_AGEMA_signal_11452, mcs1_mcs_mat1_0_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, mcs1_mcs_mat1_0_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_12411, new_AGEMA_signal_12410, mcs1_mcs_mat1_0_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_10477, new_AGEMA_signal_10476, mcs1_mcs_mat1_0_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .c ({new_AGEMA_signal_11453, new_AGEMA_signal_11452, mcs1_mcs_mat1_0_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_10477, new_AGEMA_signal_10476, mcs1_mcs_mat1_0_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9517, new_AGEMA_signal_9516, mcs1_mcs_mat1_0_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_11455, new_AGEMA_signal_11454, mcs1_mcs_mat1_0_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_9521, new_AGEMA_signal_9520, mcs1_mcs_mat1_0_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_8177, new_AGEMA_signal_8176, mcs1_mcs_mat1_0_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_10477, new_AGEMA_signal_10476, mcs1_mcs_mat1_0_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_8899, new_AGEMA_signal_8898, mcs1_mcs_mat1_0_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, mcs1_mcs_mat1_0_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_10479, new_AGEMA_signal_10478, mcs1_mcs_mat1_0_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_7671, new_AGEMA_signal_7670, mcs1_mcs_mat1_0_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_8901, new_AGEMA_signal_8900, mcs1_mcs_mat1_0_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, mcs1_mcs_mat1_0_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_8177, new_AGEMA_signal_8176, mcs1_mcs_mat1_0_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_8899, new_AGEMA_signal_8898, mcs1_mcs_mat1_0_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353]}), .c ({new_AGEMA_signal_9521, new_AGEMA_signal_9520, mcs1_mcs_mat1_0_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_8177, new_AGEMA_signal_8176, mcs1_mcs_mat1_0_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359]}), .c ({new_AGEMA_signal_8901, new_AGEMA_signal_8900, mcs1_mcs_mat1_0_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_10483, new_AGEMA_signal_10482, mcs1_mcs_mat1_0_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_8179, new_AGEMA_signal_8178, mcs1_mcs_mat1_0_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_11457, new_AGEMA_signal_11456, mcs1_mcs_mat1_0_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_8903, new_AGEMA_signal_8902, mcs1_mcs_mat1_0_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_8905, new_AGEMA_signal_8904, mcs1_mcs_mat1_0_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_9523, new_AGEMA_signal_9522, mcs1_mcs_mat1_0_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_10485, new_AGEMA_signal_10484, mcs1_mcs_mat1_0_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_11459, new_AGEMA_signal_11458, mcs1_mcs_mat1_0_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_12413, new_AGEMA_signal_12412, mcs1_mcs_mat1_0_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_10483, new_AGEMA_signal_10482, mcs1_mcs_mat1_0_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_11459, new_AGEMA_signal_11458, mcs1_mcs_mat1_0_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_7673, new_AGEMA_signal_7672, mcs1_mcs_mat1_0_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9527, new_AGEMA_signal_9526, mcs1_mcs_mat1_0_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_10483, new_AGEMA_signal_10482, mcs1_mcs_mat1_0_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_8181, new_AGEMA_signal_8180, mcs1_mcs_mat1_0_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, mcs1_mcs_mat1_0_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_10485, new_AGEMA_signal_10484, mcs1_mcs_mat1_0_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_9527, new_AGEMA_signal_9526, mcs1_mcs_mat1_0_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365]}), .c ({new_AGEMA_signal_8181, new_AGEMA_signal_8180, mcs1_mcs_mat1_0_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_8905, new_AGEMA_signal_8904, mcs1_mcs_mat1_0_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({new_AGEMA_signal_14423, new_AGEMA_signal_14422, mcs1_mcs_mat1_0_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_14913, new_AGEMA_signal_14912, mcs1_mcs_mat1_0_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({new_AGEMA_signal_14425, new_AGEMA_signal_14424, mcs1_mcs_mat1_0_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_14915, new_AGEMA_signal_14914, mcs1_mcs_mat1_0_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_13031, new_AGEMA_signal_13030, mcs1_mcs_mat1_0_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_14423, new_AGEMA_signal_14422, mcs1_mcs_mat1_0_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_14917, new_AGEMA_signal_14916, mcs1_mcs_mat1_0_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_11461, new_AGEMA_signal_11460, mcs1_mcs_mat1_0_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_14005, new_AGEMA_signal_14004, mcs1_mcs_mat1_0_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_14423, new_AGEMA_signal_14422, mcs1_mcs_mat1_0_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_13521, new_AGEMA_signal_13520, mcs1_mcs_mat1_0_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_14425, new_AGEMA_signal_14424, mcs1_mcs_mat1_0_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_14919, new_AGEMA_signal_14918, mcs1_mcs_mat1_0_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_14007, new_AGEMA_signal_14006, mcs1_mcs_mat1_0_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_14425, new_AGEMA_signal_14424, mcs1_mcs_mat1_0_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_13031, new_AGEMA_signal_13030, mcs1_mcs_mat1_0_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_13523, new_AGEMA_signal_13522, mcs1_mcs_mat1_0_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_14007, new_AGEMA_signal_14006, mcs1_mcs_mat1_0_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371]}), .c ({new_AGEMA_signal_13523, new_AGEMA_signal_13522, mcs1_mcs_mat1_0_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_11461, new_AGEMA_signal_11460, mcs1_mcs_mat1_0_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377]}), .c ({new_AGEMA_signal_13031, new_AGEMA_signal_13030, mcs1_mcs_mat1_0_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_10491, new_AGEMA_signal_10490, mcs1_mcs_mat1_0_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_10489, new_AGEMA_signal_10488, mcs1_mcs_mat1_0_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_11463, new_AGEMA_signal_11462, mcs1_mcs_mat1_0_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_10489, new_AGEMA_signal_10488, mcs1_mcs_mat1_0_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_8907, new_AGEMA_signal_8906, mcs1_mcs_mat1_0_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_11465, new_AGEMA_signal_11464, mcs1_mcs_mat1_0_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_8183, new_AGEMA_signal_8182, mcs1_mcs_mat1_0_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .c ({new_AGEMA_signal_8907, new_AGEMA_signal_8906, mcs1_mcs_mat1_0_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_10489, new_AGEMA_signal_10488, mcs1_mcs_mat1_0_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_11467, new_AGEMA_signal_11466, mcs1_mcs_mat1_0_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, mcs1_mcs_mat1_0_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_7675, new_AGEMA_signal_7674, mcs1_mcs_mat1_0_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_10489, new_AGEMA_signal_10488, mcs1_mcs_mat1_0_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_11469, new_AGEMA_signal_11468, mcs1_mcs_mat1_0_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_12415, new_AGEMA_signal_12414, mcs1_mcs_mat1_0_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_10491, new_AGEMA_signal_10490, mcs1_mcs_mat1_0_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, mcs1_mcs_mat1_0_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_11469, new_AGEMA_signal_11468, mcs1_mcs_mat1_0_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_9529, new_AGEMA_signal_9528, mcs1_mcs_mat1_0_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .c ({new_AGEMA_signal_10491, new_AGEMA_signal_10490, mcs1_mcs_mat1_0_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_8183, new_AGEMA_signal_8182, mcs1_mcs_mat1_0_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_8909, new_AGEMA_signal_8908, mcs1_mcs_mat1_0_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_9529, new_AGEMA_signal_9528, mcs1_mcs_mat1_0_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, mcs1_mcs_mat1_0_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383]}), .c ({new_AGEMA_signal_8183, new_AGEMA_signal_8182, mcs1_mcs_mat1_0_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_8909, new_AGEMA_signal_8908, mcs1_mcs_mat1_0_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_8911, new_AGEMA_signal_8910, mcs1_mcs_mat1_0_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_10493, new_AGEMA_signal_10492, mcs1_mcs_mat1_0_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_11471, new_AGEMA_signal_11470, mcs1_mcs_mat1_0_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_9539, new_AGEMA_signal_9538, mcs1_mcs_mat1_0_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_10493, new_AGEMA_signal_10492, mcs1_mcs_mat1_0_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_9535, new_AGEMA_signal_9534, mcs1_mcs_mat1_0_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_8913, new_AGEMA_signal_8912, mcs1_mcs_mat1_0_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_10495, new_AGEMA_signal_10494, mcs1_mcs_mat1_0_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, mcs1_mcs_mat1_0_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_10497, new_AGEMA_signal_10496, mcs1_mcs_mat1_0_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_11473, new_AGEMA_signal_11472, mcs1_mcs_mat1_0_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_7677, new_AGEMA_signal_7676, mcs1_mcs_mat1_0_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_9539, new_AGEMA_signal_9538, mcs1_mcs_mat1_0_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_10497, new_AGEMA_signal_10496, mcs1_mcs_mat1_0_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_8185, new_AGEMA_signal_8184, mcs1_mcs_mat1_0_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .c ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, mcs1_mcs_mat1_0_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389]}), .c ({new_AGEMA_signal_9539, new_AGEMA_signal_9538, mcs1_mcs_mat1_0_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_8185, new_AGEMA_signal_8184, mcs1_mcs_mat1_0_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395]}), .c ({new_AGEMA_signal_8913, new_AGEMA_signal_8912, mcs1_mcs_mat1_0_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_13033, new_AGEMA_signal_13032, mcs1_mcs_mat1_0_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_8917, new_AGEMA_signal_8916, mcs1_mcs_mat1_0_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_13525, new_AGEMA_signal_13524, mcs1_mcs_mat1_0_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_12417, new_AGEMA_signal_12416, mcs1_mcs_mat1_0_mcs_out[99]}), .b ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .c ({new_AGEMA_signal_13033, new_AGEMA_signal_13032, mcs1_mcs_mat1_0_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_11475, new_AGEMA_signal_11474, mcs1_mcs_mat1_0_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .c ({new_AGEMA_signal_12417, new_AGEMA_signal_12416, mcs1_mcs_mat1_0_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_10499, new_AGEMA_signal_10498, mcs1_mcs_mat1_0_mcs_out[98]}), .b ({new_AGEMA_signal_8189, new_AGEMA_signal_8188, mcs1_mcs_mat1_0_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_11475, new_AGEMA_signal_11474, mcs1_mcs_mat1_0_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_8187, new_AGEMA_signal_8186, mcs1_mcs_mat1_0_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_9541, new_AGEMA_signal_9540, mcs1_mcs_mat1_0_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_10499, new_AGEMA_signal_10498, mcs1_mcs_mat1_0_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_9541, new_AGEMA_signal_9540, mcs1_mcs_mat1_0_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401]}), .c ({new_AGEMA_signal_8189, new_AGEMA_signal_8188, mcs1_mcs_mat1_0_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_8917, new_AGEMA_signal_8916, mcs1_mcs_mat1_0_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_14009, new_AGEMA_signal_14008, mcs1_mcs_mat1_0_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_14427, new_AGEMA_signal_14426, mcs1_mcs_mat1_0_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_13037, new_AGEMA_signal_13036, mcs1_mcs_mat1_0_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_13039, new_AGEMA_signal_13038, mcs1_mcs_mat1_0_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_13529, new_AGEMA_signal_13528, mcs1_mcs_mat1_0_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_14429, new_AGEMA_signal_14428, mcs1_mcs_mat1_0_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_11477, new_AGEMA_signal_11476, mcs1_mcs_mat1_0_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_14921, new_AGEMA_signal_14920, mcs1_mcs_mat1_0_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_14009, new_AGEMA_signal_14008, mcs1_mcs_mat1_0_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_14429, new_AGEMA_signal_14428, mcs1_mcs_mat1_0_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_10501, new_AGEMA_signal_10500, mcs1_mcs_mat1_0_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_13531, new_AGEMA_signal_13530, mcs1_mcs_mat1_0_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_14009, new_AGEMA_signal_14008, mcs1_mcs_mat1_0_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407]}), .c ({new_AGEMA_signal_13531, new_AGEMA_signal_13530, mcs1_mcs_mat1_0_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_11477, new_AGEMA_signal_11476, mcs1_mcs_mat1_0_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413]}), .c ({new_AGEMA_signal_13039, new_AGEMA_signal_13038, mcs1_mcs_mat1_0_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, mcs1_mcs_mat1_0_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_9551, new_AGEMA_signal_9550, mcs1_mcs_mat1_0_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_10505, new_AGEMA_signal_10504, mcs1_mcs_mat1_0_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_9545, new_AGEMA_signal_9544, mcs1_mcs_mat1_0_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_7681, new_AGEMA_signal_7680, mcs1_mcs_mat1_0_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_10507, new_AGEMA_signal_10506, mcs1_mcs_mat1_0_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_8923, new_AGEMA_signal_8922, mcs1_mcs_mat1_0_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_9545, new_AGEMA_signal_9544, mcs1_mcs_mat1_0_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_9547, new_AGEMA_signal_9546, mcs1_mcs_mat1_0_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_10509, new_AGEMA_signal_10508, mcs1_mcs_mat1_0_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_8191, new_AGEMA_signal_8190, mcs1_mcs_mat1_0_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_8923, new_AGEMA_signal_8922, mcs1_mcs_mat1_0_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_9547, new_AGEMA_signal_9546, mcs1_mcs_mat1_0_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_10511, new_AGEMA_signal_10510, mcs1_mcs_mat1_0_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .c ({new_AGEMA_signal_11479, new_AGEMA_signal_11478, mcs1_mcs_mat1_0_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, mcs1_mcs_mat1_0_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_8191, new_AGEMA_signal_8190, mcs1_mcs_mat1_0_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_10511, new_AGEMA_signal_10510, mcs1_mcs_mat1_0_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_9551, new_AGEMA_signal_9550, mcs1_mcs_mat1_0_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419]}), .c ({new_AGEMA_signal_8191, new_AGEMA_signal_8190, mcs1_mcs_mat1_0_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_8923, new_AGEMA_signal_8922, mcs1_mcs_mat1_0_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_14011, new_AGEMA_signal_14010, mcs1_mcs_mat1_0_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_14431, new_AGEMA_signal_14430, mcs1_mcs_mat1_0_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_13041, new_AGEMA_signal_13040, mcs1_mcs_mat1_0_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_13533, new_AGEMA_signal_13532, mcs1_mcs_mat1_0_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_14433, new_AGEMA_signal_14432, mcs1_mcs_mat1_0_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_11483, new_AGEMA_signal_11482, mcs1_mcs_mat1_0_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_14923, new_AGEMA_signal_14922, mcs1_mcs_mat1_0_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_14011, new_AGEMA_signal_14010, mcs1_mcs_mat1_0_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .c ({new_AGEMA_signal_14433, new_AGEMA_signal_14432, mcs1_mcs_mat1_0_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_10513, new_AGEMA_signal_10512, mcs1_mcs_mat1_0_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_13535, new_AGEMA_signal_13534, mcs1_mcs_mat1_0_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_14011, new_AGEMA_signal_14010, mcs1_mcs_mat1_0_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425]}), .c ({new_AGEMA_signal_13535, new_AGEMA_signal_13534, mcs1_mcs_mat1_0_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_11483, new_AGEMA_signal_11482, mcs1_mcs_mat1_0_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431]}), .c ({new_AGEMA_signal_13041, new_AGEMA_signal_13040, mcs1_mcs_mat1_0_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_11485, new_AGEMA_signal_11484, mcs1_mcs_mat1_0_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_12419, new_AGEMA_signal_12418, mcs1_mcs_mat1_0_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_10517, new_AGEMA_signal_10516, mcs1_mcs_mat1_0_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, mcs1_mcs_mat1_0_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_11485, new_AGEMA_signal_11484, mcs1_mcs_mat1_0_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_8761, new_AGEMA_signal_8760, mcs1_mcs_mat1_0_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_9553, new_AGEMA_signal_9552, mcs1_mcs_mat1_0_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, mcs1_mcs_mat1_0_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_8761, new_AGEMA_signal_8760, mcs1_mcs_mat1_0_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_10515, new_AGEMA_signal_10514, mcs1_mcs_mat1_0_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_8193, new_AGEMA_signal_8192, mcs1_mcs_mat1_0_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_8195, new_AGEMA_signal_8194, mcs1_mcs_mat1_0_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_8761, new_AGEMA_signal_8760, mcs1_mcs_mat1_0_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_8925, new_AGEMA_signal_8924, mcs1_mcs_mat1_0_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .c ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, mcs1_mcs_mat1_0_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_11487, new_AGEMA_signal_11486, mcs1_mcs_mat1_0_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_8193, new_AGEMA_signal_8192, mcs1_mcs_mat1_0_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_12421, new_AGEMA_signal_12420, mcs1_mcs_mat1_0_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_10517, new_AGEMA_signal_10516, mcs1_mcs_mat1_0_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_8925, new_AGEMA_signal_8924, mcs1_mcs_mat1_0_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_11487, new_AGEMA_signal_11486, mcs1_mcs_mat1_0_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .b ({new_AGEMA_signal_9557, new_AGEMA_signal_9556, mcs1_mcs_mat1_0_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_10517, new_AGEMA_signal_10516, mcs1_mcs_mat1_0_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_9557, new_AGEMA_signal_9556, mcs1_mcs_mat1_0_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437]}), .c ({new_AGEMA_signal_8195, new_AGEMA_signal_8194, mcs1_mcs_mat1_0_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_8925, new_AGEMA_signal_8924, mcs1_mcs_mat1_0_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_10519, new_AGEMA_signal_10518, mcs1_mcs_mat1_0_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_8927, new_AGEMA_signal_8926, mcs1_mcs_mat1_0_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_11489, new_AGEMA_signal_11488, mcs1_mcs_mat1_0_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, mcs1_mcs_mat1_0_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_11491, new_AGEMA_signal_11490, mcs1_mcs_mat1_0_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12423, new_AGEMA_signal_12422, mcs1_mcs_mat1_0_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_10519, new_AGEMA_signal_10518, mcs1_mcs_mat1_0_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_11491, new_AGEMA_signal_11490, mcs1_mcs_mat1_0_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12425, new_AGEMA_signal_12424, mcs1_mcs_mat1_0_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_8927, new_AGEMA_signal_8926, mcs1_mcs_mat1_0_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_10521, new_AGEMA_signal_10520, mcs1_mcs_mat1_0_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_11491, new_AGEMA_signal_11490, mcs1_mcs_mat1_0_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({new_AGEMA_signal_8197, new_AGEMA_signal_8196, mcs1_mcs_mat1_0_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_8927, new_AGEMA_signal_8926, mcs1_mcs_mat1_0_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_9559, new_AGEMA_signal_9558, mcs1_mcs_mat1_0_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .c ({new_AGEMA_signal_10519, new_AGEMA_signal_10518, mcs1_mcs_mat1_0_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_8929, new_AGEMA_signal_8928, mcs1_mcs_mat1_0_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7685, new_AGEMA_signal_7684, mcs1_mcs_mat1_0_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_9559, new_AGEMA_signal_9558, mcs1_mcs_mat1_0_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_10521, new_AGEMA_signal_10520, mcs1_mcs_mat1_0_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, mcs1_mcs_mat1_0_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_11493, new_AGEMA_signal_11492, mcs1_mcs_mat1_0_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_8929, new_AGEMA_signal_8928, mcs1_mcs_mat1_0_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, mcs1_mcs_mat1_0_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({new_AGEMA_signal_9563, new_AGEMA_signal_9562, mcs1_mcs_mat1_0_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_10521, new_AGEMA_signal_10520, mcs1_mcs_mat1_0_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443]}), .c ({new_AGEMA_signal_9563, new_AGEMA_signal_9562, mcs1_mcs_mat1_0_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_8197, new_AGEMA_signal_8196, mcs1_mcs_mat1_0_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449]}), .c ({new_AGEMA_signal_8929, new_AGEMA_signal_8928, mcs1_mcs_mat1_0_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_11497, new_AGEMA_signal_11496, mcs1_mcs_mat1_0_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_12427, new_AGEMA_signal_12426, mcs1_mcs_mat1_0_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({new_AGEMA_signal_10523, new_AGEMA_signal_10522, mcs1_mcs_mat1_0_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_11495, new_AGEMA_signal_11494, mcs1_mcs_mat1_0_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_12429, new_AGEMA_signal_12428, mcs1_mcs_mat1_0_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_8931, new_AGEMA_signal_8930, mcs1_mcs_mat1_0_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_13043, new_AGEMA_signal_13042, mcs1_mcs_mat1_0_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_11497, new_AGEMA_signal_11496, mcs1_mcs_mat1_0_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .c ({new_AGEMA_signal_12429, new_AGEMA_signal_12428, mcs1_mcs_mat1_0_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_8199, new_AGEMA_signal_8198, mcs1_mcs_mat1_0_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_10523, new_AGEMA_signal_10522, mcs1_mcs_mat1_0_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_11497, new_AGEMA_signal_11496, mcs1_mcs_mat1_0_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_7687, new_AGEMA_signal_7686, mcs1_mcs_mat1_0_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, mcs1_mcs_mat1_0_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_10523, new_AGEMA_signal_10522, mcs1_mcs_mat1_0_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, mcs1_mcs_mat1_0_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455]}), .c ({new_AGEMA_signal_8199, new_AGEMA_signal_8198, mcs1_mcs_mat1_0_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_8931, new_AGEMA_signal_8930, mcs1_mcs_mat1_0_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_14017, new_AGEMA_signal_14016, mcs1_mcs_mat1_0_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_13045, new_AGEMA_signal_13044, mcs1_mcs_mat1_0_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_14435, new_AGEMA_signal_14434, mcs1_mcs_mat1_0_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_11499, new_AGEMA_signal_11498, mcs1_mcs_mat1_0_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_13537, new_AGEMA_signal_13536, mcs1_mcs_mat1_0_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_14013, new_AGEMA_signal_14012, mcs1_mcs_mat1_0_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({new_AGEMA_signal_13539, new_AGEMA_signal_13538, mcs1_mcs_mat1_0_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_14015, new_AGEMA_signal_14014, mcs1_mcs_mat1_0_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461]}), .c ({new_AGEMA_signal_13539, new_AGEMA_signal_13538, mcs1_mcs_mat1_0_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_11499, new_AGEMA_signal_11498, mcs1_mcs_mat1_0_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467]}), .c ({new_AGEMA_signal_13045, new_AGEMA_signal_13044, mcs1_mcs_mat1_0_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_8203, new_AGEMA_signal_8202, mcs1_mcs_mat1_0_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_8933, new_AGEMA_signal_8932, mcs1_mcs_mat1_0_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_9569, new_AGEMA_signal_9568, mcs1_mcs_mat1_0_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_8205, new_AGEMA_signal_8204, mcs1_mcs_mat1_0_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_9571, new_AGEMA_signal_9570, mcs1_mcs_mat1_0_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_10529, new_AGEMA_signal_10528, mcs1_mcs_mat1_0_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_10531, new_AGEMA_signal_10530, mcs1_mcs_mat1_0_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, mcs1_mcs_mat1_0_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_11501, new_AGEMA_signal_11500, mcs1_mcs_mat1_0_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_9575, new_AGEMA_signal_9574, mcs1_mcs_mat1_0_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_10531, new_AGEMA_signal_10530, mcs1_mcs_mat1_0_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_9575, new_AGEMA_signal_9574, mcs1_mcs_mat1_0_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473]}), .c ({new_AGEMA_signal_8205, new_AGEMA_signal_8204, mcs1_mcs_mat1_0_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_8933, new_AGEMA_signal_8932, mcs1_mcs_mat1_0_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, mcs1_mcs_mat1_0_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_10533, new_AGEMA_signal_10532, mcs1_mcs_mat1_0_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_11503, new_AGEMA_signal_11502, mcs1_mcs_mat1_0_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_11505, new_AGEMA_signal_11504, mcs1_mcs_mat1_0_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_9577, new_AGEMA_signal_9576, mcs1_mcs_mat1_0_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_12431, new_AGEMA_signal_12430, mcs1_mcs_mat1_0_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_8935, new_AGEMA_signal_8934, mcs1_mcs_mat1_0_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_9577, new_AGEMA_signal_9576, mcs1_mcs_mat1_0_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({new_AGEMA_signal_11505, new_AGEMA_signal_11504, mcs1_mcs_mat1_0_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_12433, new_AGEMA_signal_12432, mcs1_mcs_mat1_0_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_7691, new_AGEMA_signal_7690, mcs1_mcs_mat1_0_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_10533, new_AGEMA_signal_10532, mcs1_mcs_mat1_0_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_11505, new_AGEMA_signal_11504, mcs1_mcs_mat1_0_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_8207, new_AGEMA_signal_8206, mcs1_mcs_mat1_0_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_9583, new_AGEMA_signal_9582, mcs1_mcs_mat1_0_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_10533, new_AGEMA_signal_10532, mcs1_mcs_mat1_0_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_9581, new_AGEMA_signal_9580, mcs1_mcs_mat1_0_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_10535, new_AGEMA_signal_10534, mcs1_mcs_mat1_0_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_11507, new_AGEMA_signal_11506, mcs1_mcs_mat1_0_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, mcs1_mcs_mat1_0_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8207, new_AGEMA_signal_8206, mcs1_mcs_mat1_0_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_10535, new_AGEMA_signal_10534, mcs1_mcs_mat1_0_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_8935, new_AGEMA_signal_8934, mcs1_mcs_mat1_0_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, mcs1_mcs_mat1_0_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479]}), .c ({new_AGEMA_signal_9583, new_AGEMA_signal_9582, mcs1_mcs_mat1_0_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_8207, new_AGEMA_signal_8206, mcs1_mcs_mat1_0_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485]}), .c ({new_AGEMA_signal_8935, new_AGEMA_signal_8934, mcs1_mcs_mat1_0_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_13049, new_AGEMA_signal_13048, mcs1_mcs_mat1_0_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_13541, new_AGEMA_signal_13540, mcs1_mcs_mat1_0_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_14927, new_AGEMA_signal_14926, mcs1_mcs_mat1_0_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_11509, new_AGEMA_signal_11508, mcs1_mcs_mat1_0_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_15519, new_AGEMA_signal_15518, mcs1_mcs_mat1_0_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_14439, new_AGEMA_signal_14438, mcs1_mcs_mat1_0_mcs_out[47]}), .b ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_14927, new_AGEMA_signal_14926, mcs1_mcs_mat1_0_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_14019, new_AGEMA_signal_14018, mcs1_mcs_mat1_0_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .c ({new_AGEMA_signal_14439, new_AGEMA_signal_14438, mcs1_mcs_mat1_0_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_10539, new_AGEMA_signal_10538, mcs1_mcs_mat1_0_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_13543, new_AGEMA_signal_13542, mcs1_mcs_mat1_0_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_14019, new_AGEMA_signal_14018, mcs1_mcs_mat1_0_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_13543, new_AGEMA_signal_13542, mcs1_mcs_mat1_0_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491]}), .c ({new_AGEMA_signal_11509, new_AGEMA_signal_11508, mcs1_mcs_mat1_0_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_13049, new_AGEMA_signal_13048, mcs1_mcs_mat1_0_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_10541, new_AGEMA_signal_10540, mcs1_mcs_mat1_0_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_8937, new_AGEMA_signal_8936, mcs1_mcs_mat1_0_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_11511, new_AGEMA_signal_11510, mcs1_mcs_mat1_0_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_9587, new_AGEMA_signal_9586, mcs1_mcs_mat1_0_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8209, new_AGEMA_signal_8208, mcs1_mcs_mat1_0_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_10541, new_AGEMA_signal_10540, mcs1_mcs_mat1_0_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_10543, new_AGEMA_signal_10542, mcs1_mcs_mat1_0_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, mcs1_mcs_mat1_0_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_11513, new_AGEMA_signal_11512, mcs1_mcs_mat1_0_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_10545, new_AGEMA_signal_10544, mcs1_mcs_mat1_0_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_7693, new_AGEMA_signal_7692, mcs1_mcs_mat1_0_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_11515, new_AGEMA_signal_11514, mcs1_mcs_mat1_0_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_9587, new_AGEMA_signal_9586, mcs1_mcs_mat1_0_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8939, new_AGEMA_signal_8938, mcs1_mcs_mat1_0_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_10545, new_AGEMA_signal_10544, mcs1_mcs_mat1_0_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_9589, new_AGEMA_signal_9588, mcs1_mcs_mat1_0_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_8939, new_AGEMA_signal_8938, mcs1_mcs_mat1_0_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_10547, new_AGEMA_signal_10546, mcs1_mcs_mat1_0_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497]}), .c ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, mcs1_mcs_mat1_0_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_8209, new_AGEMA_signal_8208, mcs1_mcs_mat1_0_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503]}), .c ({new_AGEMA_signal_8939, new_AGEMA_signal_8938, mcs1_mcs_mat1_0_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_11517, new_AGEMA_signal_11516, mcs1_mcs_mat1_0_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_7695, new_AGEMA_signal_7694, mcs1_mcs_mat1_0_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_12435, new_AGEMA_signal_12434, mcs1_mcs_mat1_0_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_8943, new_AGEMA_signal_8942, mcs1_mcs_mat1_0_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_8941, new_AGEMA_signal_8940, mcs1_mcs_mat1_0_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_9593, new_AGEMA_signal_9592, mcs1_mcs_mat1_0_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({new_AGEMA_signal_11517, new_AGEMA_signal_11516, mcs1_mcs_mat1_0_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_12437, new_AGEMA_signal_12436, mcs1_mcs_mat1_0_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_9595, new_AGEMA_signal_9594, mcs1_mcs_mat1_0_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_10549, new_AGEMA_signal_10548, mcs1_mcs_mat1_0_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_11517, new_AGEMA_signal_11516, mcs1_mcs_mat1_0_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, mcs1_mcs_mat1_0_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_8945, new_AGEMA_signal_8944, mcs1_mcs_mat1_0_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_10549, new_AGEMA_signal_10548, mcs1_mcs_mat1_0_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, mcs1_mcs_mat1_0_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_8943, new_AGEMA_signal_8942, mcs1_mcs_mat1_0_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_10551, new_AGEMA_signal_10550, mcs1_mcs_mat1_0_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_8763, new_AGEMA_signal_8762, mcs1_mcs_mat1_0_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_8943, new_AGEMA_signal_8942, mcs1_mcs_mat1_0_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({new_AGEMA_signal_8211, new_AGEMA_signal_8210, mcs1_mcs_mat1_0_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_8763, new_AGEMA_signal_8762, mcs1_mcs_mat1_0_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, mcs1_mcs_mat1_0_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509]}), .c ({new_AGEMA_signal_8211, new_AGEMA_signal_8210, mcs1_mcs_mat1_0_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_8945, new_AGEMA_signal_8944, mcs1_mcs_mat1_0_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_9599, new_AGEMA_signal_9598, mcs1_mcs_mat1_0_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_8947, new_AGEMA_signal_8946, mcs1_mcs_mat1_0_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_10553, new_AGEMA_signal_10552, mcs1_mcs_mat1_0_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_8213, new_AGEMA_signal_8212, mcs1_mcs_mat1_0_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_8765, new_AGEMA_signal_8764, mcs1_mcs_mat1_0_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_12439, new_AGEMA_signal_12438, mcs1_mcs_mat1_0_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_9601, new_AGEMA_signal_9600, mcs1_mcs_mat1_0_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_13051, new_AGEMA_signal_13050, mcs1_mcs_mat1_0_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515]}), .c ({new_AGEMA_signal_9601, new_AGEMA_signal_9600, mcs1_mcs_mat1_0_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_8213, new_AGEMA_signal_8212, mcs1_mcs_mat1_0_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521]}), .c ({new_AGEMA_signal_8947, new_AGEMA_signal_8946, mcs1_mcs_mat1_0_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_14441, new_AGEMA_signal_14440, mcs1_mcs_mat1_0_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_14021, new_AGEMA_signal_14020, mcs1_mcs_mat1_0_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_14929, new_AGEMA_signal_14928, mcs1_mcs_mat1_0_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_11523, new_AGEMA_signal_11522, mcs1_mcs_mat1_0_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_14023, new_AGEMA_signal_14022, mcs1_mcs_mat1_0_mcs_out[29]}), .c ({new_AGEMA_signal_14441, new_AGEMA_signal_14440, mcs1_mcs_mat1_0_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_11521, new_AGEMA_signal_11520, mcs1_mcs_mat1_0_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_14021, new_AGEMA_signal_14020, mcs1_mcs_mat1_0_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_14443, new_AGEMA_signal_14442, mcs1_mcs_mat1_0_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_13549, new_AGEMA_signal_13548, mcs1_mcs_mat1_0_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .c ({new_AGEMA_signal_14021, new_AGEMA_signal_14020, mcs1_mcs_mat1_0_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_14445, new_AGEMA_signal_14444, mcs1_mcs_mat1_0_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_13545, new_AGEMA_signal_13544, mcs1_mcs_mat1_0_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_14931, new_AGEMA_signal_14930, mcs1_mcs_mat1_0_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_14025, new_AGEMA_signal_14024, mcs1_mcs_mat1_0_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_13547, new_AGEMA_signal_13546, mcs1_mcs_mat1_0_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_14445, new_AGEMA_signal_14444, mcs1_mcs_mat1_0_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_13053, new_AGEMA_signal_13052, mcs1_mcs_mat1_0_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_13547, new_AGEMA_signal_13546, mcs1_mcs_mat1_0_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_13549, new_AGEMA_signal_13548, mcs1_mcs_mat1_0_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_11523, new_AGEMA_signal_11522, mcs1_mcs_mat1_0_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_14025, new_AGEMA_signal_14024, mcs1_mcs_mat1_0_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_13549, new_AGEMA_signal_13548, mcs1_mcs_mat1_0_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527]}), .c ({new_AGEMA_signal_11523, new_AGEMA_signal_11522, mcs1_mcs_mat1_0_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_13053, new_AGEMA_signal_13052, mcs1_mcs_mat1_0_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, mcs1_mcs_mat1_0_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_10559, new_AGEMA_signal_10558, mcs1_mcs_mat1_0_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_8949, new_AGEMA_signal_8948, mcs1_mcs_mat1_0_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8215, new_AGEMA_signal_8214, mcs1_mcs_mat1_0_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, mcs1_mcs_mat1_0_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_10561, new_AGEMA_signal_10560, mcs1_mcs_mat1_0_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_11525, new_AGEMA_signal_11524, mcs1_mcs_mat1_0_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_9607, new_AGEMA_signal_9606, mcs1_mcs_mat1_0_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8215, new_AGEMA_signal_8214, mcs1_mcs_mat1_0_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_10561, new_AGEMA_signal_10560, mcs1_mcs_mat1_0_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_11527, new_AGEMA_signal_11526, mcs1_mcs_mat1_0_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .c ({new_AGEMA_signal_12441, new_AGEMA_signal_12440, mcs1_mcs_mat1_0_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_9607, new_AGEMA_signal_9606, mcs1_mcs_mat1_0_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_10563, new_AGEMA_signal_10562, mcs1_mcs_mat1_0_mcs_out[24]}), .c ({new_AGEMA_signal_11527, new_AGEMA_signal_11526, mcs1_mcs_mat1_0_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_9605, new_AGEMA_signal_9604, mcs1_mcs_mat1_0_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .c ({new_AGEMA_signal_10563, new_AGEMA_signal_10562, mcs1_mcs_mat1_0_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_8949, new_AGEMA_signal_8948, mcs1_mcs_mat1_0_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7699, new_AGEMA_signal_7698, mcs1_mcs_mat1_0_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_9605, new_AGEMA_signal_9604, mcs1_mcs_mat1_0_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533]}), .c ({new_AGEMA_signal_9607, new_AGEMA_signal_9606, mcs1_mcs_mat1_0_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_8215, new_AGEMA_signal_8214, mcs1_mcs_mat1_0_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1541], Fresh[1540], Fresh[1539]}), .c ({new_AGEMA_signal_8949, new_AGEMA_signal_8948, mcs1_mcs_mat1_0_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, mcs1_mcs_mat1_0_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .c ({new_AGEMA_signal_10565, new_AGEMA_signal_10564, mcs1_mcs_mat1_0_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_8951, new_AGEMA_signal_8950, mcs1_mcs_mat1_0_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8217, new_AGEMA_signal_8216, mcs1_mcs_mat1_0_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, mcs1_mcs_mat1_0_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_10567, new_AGEMA_signal_10566, mcs1_mcs_mat1_0_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .c ({new_AGEMA_signal_11529, new_AGEMA_signal_11528, mcs1_mcs_mat1_0_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_9613, new_AGEMA_signal_9612, mcs1_mcs_mat1_0_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8217, new_AGEMA_signal_8216, mcs1_mcs_mat1_0_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_10567, new_AGEMA_signal_10566, mcs1_mcs_mat1_0_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_11531, new_AGEMA_signal_11530, mcs1_mcs_mat1_0_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_12443, new_AGEMA_signal_12442, mcs1_mcs_mat1_0_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_9613, new_AGEMA_signal_9612, mcs1_mcs_mat1_0_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_10569, new_AGEMA_signal_10568, mcs1_mcs_mat1_0_mcs_out[20]}), .c ({new_AGEMA_signal_11531, new_AGEMA_signal_11530, mcs1_mcs_mat1_0_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_9611, new_AGEMA_signal_9610, mcs1_mcs_mat1_0_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_10569, new_AGEMA_signal_10568, mcs1_mcs_mat1_0_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_8951, new_AGEMA_signal_8950, mcs1_mcs_mat1_0_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7701, new_AGEMA_signal_7700, mcs1_mcs_mat1_0_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_9611, new_AGEMA_signal_9610, mcs1_mcs_mat1_0_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({new_AGEMA_signal_9613, new_AGEMA_signal_9612, mcs1_mcs_mat1_0_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1547], Fresh[1546], Fresh[1545]}), .c ({new_AGEMA_signal_8217, new_AGEMA_signal_8216, mcs1_mcs_mat1_0_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_8951, new_AGEMA_signal_8950, mcs1_mcs_mat1_0_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, mcs1_mcs_mat1_0_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, mcs1_mcs_mat1_0_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_10571, new_AGEMA_signal_10570, mcs1_mcs_mat1_0_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_10573, new_AGEMA_signal_10572, mcs1_mcs_mat1_0_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_7703, new_AGEMA_signal_7702, mcs1_mcs_mat1_0_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_11533, new_AGEMA_signal_11532, mcs1_mcs_mat1_0_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_11535, new_AGEMA_signal_11534, mcs1_mcs_mat1_0_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_8219, new_AGEMA_signal_8218, mcs1_mcs_mat1_0_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_12445, new_AGEMA_signal_12444, mcs1_mcs_mat1_0_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_10573, new_AGEMA_signal_10572, mcs1_mcs_mat1_0_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_11535, new_AGEMA_signal_11534, mcs1_mcs_mat1_0_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_9617, new_AGEMA_signal_9616, mcs1_mcs_mat1_0_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .c ({new_AGEMA_signal_10573, new_AGEMA_signal_10572, mcs1_mcs_mat1_0_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_8953, new_AGEMA_signal_8952, mcs1_mcs_mat1_0_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_8955, new_AGEMA_signal_8954, mcs1_mcs_mat1_0_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_9617, new_AGEMA_signal_9616, mcs1_mcs_mat1_0_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_9619, new_AGEMA_signal_9618, mcs1_mcs_mat1_0_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_8219, new_AGEMA_signal_8218, mcs1_mcs_mat1_0_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_10575, new_AGEMA_signal_10574, mcs1_mcs_mat1_0_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1553], Fresh[1552], Fresh[1551]}), .c ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, mcs1_mcs_mat1_0_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({new_AGEMA_signal_8219, new_AGEMA_signal_8218, mcs1_mcs_mat1_0_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1559], Fresh[1558], Fresh[1557]}), .c ({new_AGEMA_signal_8955, new_AGEMA_signal_8954, mcs1_mcs_mat1_0_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_14451, new_AGEMA_signal_14450, mcs1_mcs_mat1_0_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_12447, new_AGEMA_signal_12446, mcs1_mcs_mat1_0_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_14933, new_AGEMA_signal_14932, mcs1_mcs_mat1_0_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_14031, new_AGEMA_signal_14030, mcs1_mcs_mat1_0_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_14027, new_AGEMA_signal_14026, mcs1_mcs_mat1_0_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_14447, new_AGEMA_signal_14446, mcs1_mcs_mat1_0_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_13553, new_AGEMA_signal_13552, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_11537, new_AGEMA_signal_11536, mcs1_mcs_mat1_0_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_14027, new_AGEMA_signal_14026, mcs1_mcs_mat1_0_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_12447, new_AGEMA_signal_12446, mcs1_mcs_mat1_0_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_14029, new_AGEMA_signal_14028, mcs1_mcs_mat1_0_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_14449, new_AGEMA_signal_14448, mcs1_mcs_mat1_0_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_13551, new_AGEMA_signal_13550, mcs1_mcs_mat1_0_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_13553, new_AGEMA_signal_13552, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_14029, new_AGEMA_signal_14028, mcs1_mcs_mat1_0_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_10577, new_AGEMA_signal_10576, mcs1_mcs_mat1_0_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_11537, new_AGEMA_signal_11536, mcs1_mcs_mat1_0_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_12447, new_AGEMA_signal_12446, mcs1_mcs_mat1_0_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_14935, new_AGEMA_signal_14934, mcs1_mcs_mat1_0_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_15521, new_AGEMA_signal_15520, mcs1_mcs_mat1_0_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_14451, new_AGEMA_signal_14450, mcs1_mcs_mat1_0_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_13553, new_AGEMA_signal_13552, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_14935, new_AGEMA_signal_14934, mcs1_mcs_mat1_0_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_14031, new_AGEMA_signal_14030, mcs1_mcs_mat1_0_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_14451, new_AGEMA_signal_14450, mcs1_mcs_mat1_0_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_13551, new_AGEMA_signal_13550, mcs1_mcs_mat1_0_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_14031, new_AGEMA_signal_14030, mcs1_mcs_mat1_0_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, shiftr_out[124]}), .b ({new_AGEMA_signal_13055, new_AGEMA_signal_13054, mcs1_mcs_mat1_0_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_13551, new_AGEMA_signal_13550, mcs1_mcs_mat1_0_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12983, new_AGEMA_signal_12982, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_13553, new_AGEMA_signal_13552, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1565], Fresh[1564], Fresh[1563]}), .c ({new_AGEMA_signal_11537, new_AGEMA_signal_11536, mcs1_mcs_mat1_0_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({new_AGEMA_signal_13055, new_AGEMA_signal_13054, mcs1_mcs_mat1_0_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_8767, new_AGEMA_signal_8766, mcs1_mcs_mat1_0_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .c ({new_AGEMA_signal_8957, new_AGEMA_signal_8956, mcs1_mcs_mat1_0_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_10581, new_AGEMA_signal_10580, mcs1_mcs_mat1_0_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_11539, new_AGEMA_signal_11538, mcs1_mcs_mat1_0_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_9623, new_AGEMA_signal_9622, mcs1_mcs_mat1_0_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_10579, new_AGEMA_signal_10578, mcs1_mcs_mat1_0_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_8959, new_AGEMA_signal_8958, mcs1_mcs_mat1_0_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_8767, new_AGEMA_signal_8766, mcs1_mcs_mat1_0_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_9623, new_AGEMA_signal_9622, mcs1_mcs_mat1_0_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_7705, new_AGEMA_signal_7704, mcs1_mcs_mat1_0_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8221, new_AGEMA_signal_8220, mcs1_mcs_mat1_0_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_8767, new_AGEMA_signal_8766, mcs1_mcs_mat1_0_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_11541, new_AGEMA_signal_11540, mcs1_mcs_mat1_0_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, shiftr_out[92]}), .c ({new_AGEMA_signal_12449, new_AGEMA_signal_12448, mcs1_mcs_mat1_0_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_7705, new_AGEMA_signal_7704, mcs1_mcs_mat1_0_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_10581, new_AGEMA_signal_10580, mcs1_mcs_mat1_0_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_11541, new_AGEMA_signal_11540, mcs1_mcs_mat1_0_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_9625, new_AGEMA_signal_9624, mcs1_mcs_mat1_0_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_8959, new_AGEMA_signal_8958, mcs1_mcs_mat1_0_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_10581, new_AGEMA_signal_10580, mcs1_mcs_mat1_0_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8867, new_AGEMA_signal_8866, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1571], Fresh[1570], Fresh[1569]}), .c ({new_AGEMA_signal_9625, new_AGEMA_signal_9624, mcs1_mcs_mat1_0_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7643, new_AGEMA_signal_7642, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_8221, new_AGEMA_signal_8220, mcs1_mcs_mat1_0_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8735, new_AGEMA_signal_8734, shiftr_out[95]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1577], Fresh[1576], Fresh[1575]}), .c ({new_AGEMA_signal_8959, new_AGEMA_signal_8958, mcs1_mcs_mat1_0_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_13057, new_AGEMA_signal_13056, mcs1_mcs_mat1_0_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_8963, new_AGEMA_signal_8962, mcs1_mcs_mat1_0_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_13555, new_AGEMA_signal_13554, mcs1_mcs_mat1_0_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_12451, new_AGEMA_signal_12450, mcs1_mcs_mat1_0_mcs_out[7]}), .b ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .c ({new_AGEMA_signal_13057, new_AGEMA_signal_13056, mcs1_mcs_mat1_0_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_11543, new_AGEMA_signal_11542, mcs1_mcs_mat1_0_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .c ({new_AGEMA_signal_12451, new_AGEMA_signal_12450, mcs1_mcs_mat1_0_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_10583, new_AGEMA_signal_10582, mcs1_mcs_mat1_0_mcs_out[6]}), .b ({new_AGEMA_signal_8225, new_AGEMA_signal_8224, mcs1_mcs_mat1_0_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_11543, new_AGEMA_signal_11542, mcs1_mcs_mat1_0_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_8223, new_AGEMA_signal_8222, mcs1_mcs_mat1_0_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, mcs1_mcs_mat1_0_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_10583, new_AGEMA_signal_10582, mcs1_mcs_mat1_0_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8879, new_AGEMA_signal_8878, shiftr_out[61]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, mcs1_mcs_mat1_0_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7655, new_AGEMA_signal_7654, shiftr_out[62]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1583], Fresh[1582], Fresh[1581]}), .c ({new_AGEMA_signal_8225, new_AGEMA_signal_8224, mcs1_mcs_mat1_0_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8747, new_AGEMA_signal_8746, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_8963, new_AGEMA_signal_8962, mcs1_mcs_mat1_0_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_8965, new_AGEMA_signal_8964, mcs1_mcs_mat1_0_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_9629, new_AGEMA_signal_9628, mcs1_mcs_mat1_0_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_10587, new_AGEMA_signal_10586, mcs1_mcs_mat1_0_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .b ({new_AGEMA_signal_8967, new_AGEMA_signal_8966, mcs1_mcs_mat1_0_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_9629, new_AGEMA_signal_9628, mcs1_mcs_mat1_0_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_10589, new_AGEMA_signal_10588, mcs1_mcs_mat1_0_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_8227, new_AGEMA_signal_8226, mcs1_mcs_mat1_0_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_11545, new_AGEMA_signal_11544, mcs1_mcs_mat1_0_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_10591, new_AGEMA_signal_10590, mcs1_mcs_mat1_0_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, mcs1_mcs_mat1_0_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_11547, new_AGEMA_signal_11546, mcs1_mcs_mat1_0_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_9635, new_AGEMA_signal_9634, mcs1_mcs_mat1_0_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_7709, new_AGEMA_signal_7708, mcs1_mcs_mat1_0_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_10591, new_AGEMA_signal_10590, mcs1_mcs_mat1_0_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8891, new_AGEMA_signal_8890, shiftr_out[29]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1589], Fresh[1588], Fresh[1587]}), .c ({new_AGEMA_signal_9635, new_AGEMA_signal_9634, mcs1_mcs_mat1_0_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7667, new_AGEMA_signal_7666, shiftr_out[30]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({new_AGEMA_signal_8227, new_AGEMA_signal_8226, mcs1_mcs_mat1_0_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8759, new_AGEMA_signal_8758, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1595], Fresh[1594], Fresh[1593]}), .c ({new_AGEMA_signal_8967, new_AGEMA_signal_8966, mcs1_mcs_mat1_0_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U96 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, mcs1_mcs_mat1_1_n128}), .b ({new_AGEMA_signal_12453, new_AGEMA_signal_12452, mcs1_mcs_mat1_1_n127}), .c ({temp_next_s2[89], temp_next_s1[89], temp_next_s0[89]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U95 ( .a ({new_AGEMA_signal_11633, new_AGEMA_signal_11632, mcs1_mcs_mat1_1_mcs_out[41]}), .b ({new_AGEMA_signal_9707, new_AGEMA_signal_9706, mcs1_mcs_mat1_1_mcs_out[45]}), .c ({new_AGEMA_signal_12453, new_AGEMA_signal_12452, mcs1_mcs_mat1_1_n127}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U94 ( .a ({new_AGEMA_signal_12519, new_AGEMA_signal_12518, mcs1_mcs_mat1_1_mcs_out[33]}), .b ({new_AGEMA_signal_12517, new_AGEMA_signal_12516, mcs1_mcs_mat1_1_mcs_out[37]}), .c ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, mcs1_mcs_mat1_1_n128}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U93 ( .a ({new_AGEMA_signal_16021, new_AGEMA_signal_16020, mcs1_mcs_mat1_1_n126}), .b ({new_AGEMA_signal_13559, new_AGEMA_signal_13558, mcs1_mcs_mat1_1_n125}), .c ({temp_next_s2[88], temp_next_s1[88], temp_next_s0[88]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U92 ( .a ({new_AGEMA_signal_10667, new_AGEMA_signal_10666, mcs1_mcs_mat1_1_mcs_out[40]}), .b ({new_AGEMA_signal_13099, new_AGEMA_signal_13098, mcs1_mcs_mat1_1_mcs_out[44]}), .c ({new_AGEMA_signal_13559, new_AGEMA_signal_13558, mcs1_mcs_mat1_1_n125}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U91 ( .a ({new_AGEMA_signal_15549, new_AGEMA_signal_15548, mcs1_mcs_mat1_1_mcs_out[32]}), .b ({new_AGEMA_signal_10671, new_AGEMA_signal_10670, mcs1_mcs_mat1_1_mcs_out[36]}), .c ({new_AGEMA_signal_16021, new_AGEMA_signal_16020, mcs1_mcs_mat1_1_n126}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U90 ( .a ({new_AGEMA_signal_14453, new_AGEMA_signal_14452, mcs1_mcs_mat1_1_n124}), .b ({new_AGEMA_signal_13061, new_AGEMA_signal_13060, mcs1_mcs_mat1_1_n123}), .c ({temp_next_s2[59], temp_next_s1[59], temp_next_s0[59]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U89 ( .a ({new_AGEMA_signal_10681, new_AGEMA_signal_10680, mcs1_mcs_mat1_1_mcs_out[27]}), .b ({new_AGEMA_signal_12521, new_AGEMA_signal_12520, mcs1_mcs_mat1_1_mcs_out[31]}), .c ({new_AGEMA_signal_13061, new_AGEMA_signal_13060, mcs1_mcs_mat1_1_n123}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U88 ( .a ({new_AGEMA_signal_14067, new_AGEMA_signal_14066, mcs1_mcs_mat1_1_mcs_out[19]}), .b ({new_AGEMA_signal_10687, new_AGEMA_signal_10686, mcs1_mcs_mat1_1_mcs_out[23]}), .c ({new_AGEMA_signal_14453, new_AGEMA_signal_14452, mcs1_mcs_mat1_1_n124}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U87 ( .a ({new_AGEMA_signal_14939, new_AGEMA_signal_14938, mcs1_mcs_mat1_1_n122}), .b ({new_AGEMA_signal_12455, new_AGEMA_signal_12454, mcs1_mcs_mat1_1_n121}), .c ({temp_next_s2[58], temp_next_s1[58], temp_next_s0[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U86 ( .a ({new_AGEMA_signal_11645, new_AGEMA_signal_11644, mcs1_mcs_mat1_1_mcs_out[26]}), .b ({new_AGEMA_signal_11641, new_AGEMA_signal_11640, mcs1_mcs_mat1_1_mcs_out[30]}), .c ({new_AGEMA_signal_12455, new_AGEMA_signal_12454, mcs1_mcs_mat1_1_n121}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U85 ( .a ({new_AGEMA_signal_14495, new_AGEMA_signal_14494, mcs1_mcs_mat1_1_mcs_out[18]}), .b ({new_AGEMA_signal_11649, new_AGEMA_signal_11648, mcs1_mcs_mat1_1_mcs_out[22]}), .c ({new_AGEMA_signal_14939, new_AGEMA_signal_14938, mcs1_mcs_mat1_1_n122}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U84 ( .a ({new_AGEMA_signal_15525, new_AGEMA_signal_15524, mcs1_mcs_mat1_1_n120}), .b ({new_AGEMA_signal_13063, new_AGEMA_signal_13062, mcs1_mcs_mat1_1_n119}), .c ({temp_next_s2[57], temp_next_s1[57], temp_next_s0[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U83 ( .a ({new_AGEMA_signal_12525, new_AGEMA_signal_12524, mcs1_mcs_mat1_1_mcs_out[25]}), .b ({new_AGEMA_signal_10677, new_AGEMA_signal_10676, mcs1_mcs_mat1_1_mcs_out[29]}), .c ({new_AGEMA_signal_13063, new_AGEMA_signal_13062, mcs1_mcs_mat1_1_n119}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U82 ( .a ({new_AGEMA_signal_14983, new_AGEMA_signal_14982, mcs1_mcs_mat1_1_mcs_out[17]}), .b ({new_AGEMA_signal_12527, new_AGEMA_signal_12526, mcs1_mcs_mat1_1_mcs_out[21]}), .c ({new_AGEMA_signal_15525, new_AGEMA_signal_15524, mcs1_mcs_mat1_1_n120}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U81 ( .a ({new_AGEMA_signal_14455, new_AGEMA_signal_14454, mcs1_mcs_mat1_1_n118}), .b ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, mcs1_mcs_mat1_1_n117}), .c ({temp_next_s2[56], temp_next_s1[56], temp_next_s0[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U80 ( .a ({new_AGEMA_signal_10685, new_AGEMA_signal_10684, mcs1_mcs_mat1_1_mcs_out[24]}), .b ({new_AGEMA_signal_12523, new_AGEMA_signal_12522, mcs1_mcs_mat1_1_mcs_out[28]}), .c ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, mcs1_mcs_mat1_1_n117}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U79 ( .a ({new_AGEMA_signal_14071, new_AGEMA_signal_14070, mcs1_mcs_mat1_1_mcs_out[16]}), .b ({new_AGEMA_signal_10691, new_AGEMA_signal_10690, mcs1_mcs_mat1_1_mcs_out[20]}), .c ({new_AGEMA_signal_14455, new_AGEMA_signal_14454, mcs1_mcs_mat1_1_n118}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U78 ( .a ({new_AGEMA_signal_13067, new_AGEMA_signal_13066, mcs1_mcs_mat1_1_n116}), .b ({new_AGEMA_signal_14457, new_AGEMA_signal_14456, mcs1_mcs_mat1_1_n115}), .c ({temp_next_s2[27], temp_next_s1[27], temp_next_s0[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U77 ( .a ({new_AGEMA_signal_14073, new_AGEMA_signal_14072, mcs1_mcs_mat1_1_mcs_out[3]}), .b ({new_AGEMA_signal_12535, new_AGEMA_signal_12534, mcs1_mcs_mat1_1_mcs_out[7]}), .c ({new_AGEMA_signal_14457, new_AGEMA_signal_14456, mcs1_mcs_mat1_1_n115}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U76 ( .a ({new_AGEMA_signal_9037, new_AGEMA_signal_9036, mcs1_mcs_mat1_1_mcs_out[11]}), .b ({new_AGEMA_signal_12529, new_AGEMA_signal_12528, mcs1_mcs_mat1_1_mcs_out[15]}), .c ({new_AGEMA_signal_13067, new_AGEMA_signal_13066, mcs1_mcs_mat1_1_n116}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U75 ( .a ({new_AGEMA_signal_14945, new_AGEMA_signal_14944, mcs1_mcs_mat1_1_n114}), .b ({new_AGEMA_signal_13069, new_AGEMA_signal_13068, mcs1_mcs_mat1_1_n113}), .c ({new_AGEMA_signal_15527, new_AGEMA_signal_15526, mcs_out[251]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U74 ( .a ({new_AGEMA_signal_12477, new_AGEMA_signal_12476, mcs1_mcs_mat1_1_mcs_out[123]}), .b ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_13069, new_AGEMA_signal_13068, mcs1_mcs_mat1_1_n113}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U73 ( .a ({new_AGEMA_signal_14481, new_AGEMA_signal_14480, mcs1_mcs_mat1_1_mcs_out[115]}), .b ({new_AGEMA_signal_12481, new_AGEMA_signal_12480, mcs1_mcs_mat1_1_mcs_out[119]}), .c ({new_AGEMA_signal_14945, new_AGEMA_signal_14944, mcs1_mcs_mat1_1_n114}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U72 ( .a ({new_AGEMA_signal_14459, new_AGEMA_signal_14458, mcs1_mcs_mat1_1_n112}), .b ({new_AGEMA_signal_10593, new_AGEMA_signal_10592, mcs1_mcs_mat1_1_n111}), .c ({new_AGEMA_signal_14947, new_AGEMA_signal_14946, mcs_out[250]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U71 ( .a ({new_AGEMA_signal_9637, new_AGEMA_signal_9636, mcs1_mcs_mat1_1_mcs_out[122]}), .b ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_10593, new_AGEMA_signal_10592, mcs1_mcs_mat1_1_n111}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U70 ( .a ({new_AGEMA_signal_14043, new_AGEMA_signal_14042, mcs1_mcs_mat1_1_mcs_out[114]}), .b ({new_AGEMA_signal_12483, new_AGEMA_signal_12482, mcs1_mcs_mat1_1_mcs_out[118]}), .c ({new_AGEMA_signal_14459, new_AGEMA_signal_14458, mcs1_mcs_mat1_1_n112}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U69 ( .a ({new_AGEMA_signal_12457, new_AGEMA_signal_12456, mcs1_mcs_mat1_1_n110}), .b ({new_AGEMA_signal_14461, new_AGEMA_signal_14460, mcs1_mcs_mat1_1_n109}), .c ({temp_next_s2[26], temp_next_s1[26], temp_next_s0[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U68 ( .a ({new_AGEMA_signal_14075, new_AGEMA_signal_14074, mcs1_mcs_mat1_1_mcs_out[2]}), .b ({new_AGEMA_signal_10705, new_AGEMA_signal_10704, mcs1_mcs_mat1_1_mcs_out[6]}), .c ({new_AGEMA_signal_14461, new_AGEMA_signal_14460, mcs1_mcs_mat1_1_n109}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U67 ( .a ({new_AGEMA_signal_11661, new_AGEMA_signal_11660, mcs1_mcs_mat1_1_mcs_out[10]}), .b ({new_AGEMA_signal_11655, new_AGEMA_signal_11654, mcs1_mcs_mat1_1_mcs_out[14]}), .c ({new_AGEMA_signal_12457, new_AGEMA_signal_12456, mcs1_mcs_mat1_1_n110}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U66 ( .a ({new_AGEMA_signal_14033, new_AGEMA_signal_14032, mcs1_mcs_mat1_1_n108}), .b ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, mcs1_mcs_mat1_1_n107}), .c ({new_AGEMA_signal_14463, new_AGEMA_signal_14462, mcs_out[249]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U65 ( .a ({new_AGEMA_signal_12479, new_AGEMA_signal_12478, mcs1_mcs_mat1_1_mcs_out[121]}), .b ({new_AGEMA_signal_8969, new_AGEMA_signal_8968, mcs1_mcs_mat1_1_mcs_out[125]}), .c ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, mcs1_mcs_mat1_1_n107}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U64 ( .a ({new_AGEMA_signal_13567, new_AGEMA_signal_13566, mcs1_mcs_mat1_1_mcs_out[113]}), .b ({new_AGEMA_signal_11567, new_AGEMA_signal_11566, mcs1_mcs_mat1_1_mcs_out[117]}), .c ({new_AGEMA_signal_14033, new_AGEMA_signal_14032, mcs1_mcs_mat1_1_n108}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U63 ( .a ({new_AGEMA_signal_15529, new_AGEMA_signal_15528, mcs1_mcs_mat1_1_n106}), .b ({new_AGEMA_signal_12459, new_AGEMA_signal_12458, mcs1_mcs_mat1_1_n105}), .c ({new_AGEMA_signal_16025, new_AGEMA_signal_16024, mcs_out[248]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U62 ( .a ({new_AGEMA_signal_11561, new_AGEMA_signal_11560, mcs1_mcs_mat1_1_mcs_out[120]}), .b ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_12459, new_AGEMA_signal_12458, mcs1_mcs_mat1_1_n105}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U61 ( .a ({new_AGEMA_signal_14973, new_AGEMA_signal_14972, mcs1_mcs_mat1_1_mcs_out[112]}), .b ({new_AGEMA_signal_10605, new_AGEMA_signal_10604, mcs1_mcs_mat1_1_mcs_out[116]}), .c ({new_AGEMA_signal_15529, new_AGEMA_signal_15528, mcs1_mcs_mat1_1_n106}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U60 ( .a ({new_AGEMA_signal_12461, new_AGEMA_signal_12460, mcs1_mcs_mat1_1_n104}), .b ({new_AGEMA_signal_15531, new_AGEMA_signal_15530, mcs1_mcs_mat1_1_n103}), .c ({new_AGEMA_signal_16027, new_AGEMA_signal_16026, mcs_out[219]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U59 ( .a ({new_AGEMA_signal_12485, new_AGEMA_signal_12484, mcs1_mcs_mat1_1_mcs_out[111]}), .b ({new_AGEMA_signal_14975, new_AGEMA_signal_14974, mcs1_mcs_mat1_1_mcs_out[99]}), .c ({new_AGEMA_signal_15531, new_AGEMA_signal_15530, mcs1_mcs_mat1_1_n103}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U58 ( .a ({new_AGEMA_signal_11585, new_AGEMA_signal_11584, mcs1_mcs_mat1_1_mcs_out[103]}), .b ({new_AGEMA_signal_11577, new_AGEMA_signal_11576, mcs1_mcs_mat1_1_mcs_out[107]}), .c ({new_AGEMA_signal_12461, new_AGEMA_signal_12460, mcs1_mcs_mat1_1_n104}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U57 ( .a ({new_AGEMA_signal_12463, new_AGEMA_signal_12462, mcs1_mcs_mat1_1_n102}), .b ({new_AGEMA_signal_14465, new_AGEMA_signal_14464, mcs1_mcs_mat1_1_n101}), .c ({new_AGEMA_signal_14951, new_AGEMA_signal_14950, mcs_out[218]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U56 ( .a ({new_AGEMA_signal_12487, new_AGEMA_signal_12486, mcs1_mcs_mat1_1_mcs_out[110]}), .b ({new_AGEMA_signal_14049, new_AGEMA_signal_14048, mcs1_mcs_mat1_1_mcs_out[98]}), .c ({new_AGEMA_signal_14465, new_AGEMA_signal_14464, mcs1_mcs_mat1_1_n101}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U55 ( .a ({new_AGEMA_signal_9655, new_AGEMA_signal_9654, mcs1_mcs_mat1_1_mcs_out[102]}), .b ({new_AGEMA_signal_11579, new_AGEMA_signal_11578, mcs1_mcs_mat1_1_mcs_out[106]}), .c ({new_AGEMA_signal_12463, new_AGEMA_signal_12462, mcs1_mcs_mat1_1_n102}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U54 ( .a ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, mcs1_mcs_mat1_1_n100}), .b ({new_AGEMA_signal_13561, new_AGEMA_signal_13560, mcs1_mcs_mat1_1_n99}), .c ({new_AGEMA_signal_14035, new_AGEMA_signal_14034, mcs_out[217]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U53 ( .a ({new_AGEMA_signal_12489, new_AGEMA_signal_12488, mcs1_mcs_mat1_1_mcs_out[109]}), .b ({new_AGEMA_signal_13091, new_AGEMA_signal_13090, mcs1_mcs_mat1_1_mcs_out[97]}), .c ({new_AGEMA_signal_13561, new_AGEMA_signal_13560, mcs1_mcs_mat1_1_n99}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U52 ( .a ({new_AGEMA_signal_10619, new_AGEMA_signal_10618, mcs1_mcs_mat1_1_mcs_out[101]}), .b ({new_AGEMA_signal_11581, new_AGEMA_signal_11580, mcs1_mcs_mat1_1_mcs_out[105]}), .c ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, mcs1_mcs_mat1_1_n100}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U51 ( .a ({new_AGEMA_signal_13073, new_AGEMA_signal_13072, mcs1_mcs_mat1_1_n98}), .b ({new_AGEMA_signal_16363, new_AGEMA_signal_16362, mcs1_mcs_mat1_1_n97}), .c ({new_AGEMA_signal_16465, new_AGEMA_signal_16464, mcs_out[216]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U50 ( .a ({new_AGEMA_signal_12491, new_AGEMA_signal_12490, mcs1_mcs_mat1_1_mcs_out[108]}), .b ({new_AGEMA_signal_16033, new_AGEMA_signal_16032, mcs1_mcs_mat1_1_mcs_out[96]}), .c ({new_AGEMA_signal_16363, new_AGEMA_signal_16362, mcs1_mcs_mat1_1_n97}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U49 ( .a ({new_AGEMA_signal_11587, new_AGEMA_signal_11586, mcs1_mcs_mat1_1_mcs_out[100]}), .b ({new_AGEMA_signal_12493, new_AGEMA_signal_12492, mcs1_mcs_mat1_1_mcs_out[104]}), .c ({new_AGEMA_signal_13073, new_AGEMA_signal_13072, mcs1_mcs_mat1_1_n98}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U48 ( .a ({new_AGEMA_signal_14467, new_AGEMA_signal_14466, mcs1_mcs_mat1_1_n96}), .b ({new_AGEMA_signal_12467, new_AGEMA_signal_12466, mcs1_mcs_mat1_1_n95}), .c ({new_AGEMA_signal_14953, new_AGEMA_signal_14952, mcs_out[187]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U47 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_11593, new_AGEMA_signal_11592, mcs1_mcs_mat1_1_mcs_out[95]}), .c ({new_AGEMA_signal_12467, new_AGEMA_signal_12466, mcs1_mcs_mat1_1_n95}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U46 ( .a ({new_AGEMA_signal_14051, new_AGEMA_signal_14050, mcs1_mcs_mat1_1_mcs_out[83]}), .b ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, mcs1_mcs_mat1_1_mcs_out[87]}), .c ({new_AGEMA_signal_14467, new_AGEMA_signal_14466, mcs1_mcs_mat1_1_n96}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U45 ( .a ({new_AGEMA_signal_14469, new_AGEMA_signal_14468, mcs1_mcs_mat1_1_n94}), .b ({new_AGEMA_signal_10595, new_AGEMA_signal_10594, mcs1_mcs_mat1_1_n93}), .c ({new_AGEMA_signal_14955, new_AGEMA_signal_14954, mcs_out[186]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U43 ( .a ({new_AGEMA_signal_14053, new_AGEMA_signal_14052, mcs1_mcs_mat1_1_mcs_out[82]}), .b ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_14469, new_AGEMA_signal_14468, mcs1_mcs_mat1_1_n94}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U42 ( .a ({new_AGEMA_signal_14471, new_AGEMA_signal_14470, mcs1_mcs_mat1_1_n92}), .b ({new_AGEMA_signal_10597, new_AGEMA_signal_10596, mcs1_mcs_mat1_1_n91}), .c ({new_AGEMA_signal_14957, new_AGEMA_signal_14956, mcs_out[185]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U41 ( .a ({new_AGEMA_signal_8999, new_AGEMA_signal_8998, mcs1_mcs_mat1_1_mcs_out[89]}), .b ({new_AGEMA_signal_9665, new_AGEMA_signal_9664, mcs1_mcs_mat1_1_mcs_out[93]}), .c ({new_AGEMA_signal_10597, new_AGEMA_signal_10596, mcs1_mcs_mat1_1_n91}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U40 ( .a ({new_AGEMA_signal_14055, new_AGEMA_signal_14054, mcs1_mcs_mat1_1_mcs_out[81]}), .b ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_14471, new_AGEMA_signal_14470, mcs1_mcs_mat1_1_n92}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U39 ( .a ({new_AGEMA_signal_14959, new_AGEMA_signal_14958, mcs1_mcs_mat1_1_n90}), .b ({new_AGEMA_signal_13075, new_AGEMA_signal_13074, mcs1_mcs_mat1_1_n89}), .c ({new_AGEMA_signal_15533, new_AGEMA_signal_15532, mcs_out[184]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U38 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_12495, new_AGEMA_signal_12494, mcs1_mcs_mat1_1_mcs_out[92]}), .c ({new_AGEMA_signal_13075, new_AGEMA_signal_13074, mcs1_mcs_mat1_1_n89}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U37 ( .a ({new_AGEMA_signal_14487, new_AGEMA_signal_14486, mcs1_mcs_mat1_1_mcs_out[80]}), .b ({new_AGEMA_signal_10627, new_AGEMA_signal_10626, mcs1_mcs_mat1_1_mcs_out[84]}), .c ({new_AGEMA_signal_14959, new_AGEMA_signal_14958, mcs1_mcs_mat1_1_n90}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U36 ( .a ({new_AGEMA_signal_14961, new_AGEMA_signal_14960, mcs1_mcs_mat1_1_n88}), .b ({new_AGEMA_signal_11549, new_AGEMA_signal_11548, mcs1_mcs_mat1_1_n87}), .c ({temp_next_s2[25], temp_next_s1[25], temp_next_s0[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U35 ( .a ({new_AGEMA_signal_9041, new_AGEMA_signal_9040, mcs1_mcs_mat1_1_mcs_out[5]}), .b ({new_AGEMA_signal_10701, new_AGEMA_signal_10700, mcs1_mcs_mat1_1_mcs_out[9]}), .c ({new_AGEMA_signal_11549, new_AGEMA_signal_11548, mcs1_mcs_mat1_1_n87}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U34 ( .a ({new_AGEMA_signal_11657, new_AGEMA_signal_11656, mcs1_mcs_mat1_1_mcs_out[13]}), .b ({new_AGEMA_signal_14499, new_AGEMA_signal_14498, mcs1_mcs_mat1_1_mcs_out[1]}), .c ({new_AGEMA_signal_14961, new_AGEMA_signal_14960, mcs1_mcs_mat1_1_n88}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U33 ( .a ({new_AGEMA_signal_15537, new_AGEMA_signal_15536, mcs1_mcs_mat1_1_n86}), .b ({new_AGEMA_signal_12469, new_AGEMA_signal_12468, mcs1_mcs_mat1_1_n85}), .c ({new_AGEMA_signal_16029, new_AGEMA_signal_16028, mcs_out[155]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U32 ( .a ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, mcs1_mcs_mat1_1_mcs_out[75]}), .b ({new_AGEMA_signal_11599, new_AGEMA_signal_11598, mcs1_mcs_mat1_1_mcs_out[79]}), .c ({new_AGEMA_signal_12469, new_AGEMA_signal_12468, mcs1_mcs_mat1_1_n85}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U31 ( .a ({new_AGEMA_signal_14977, new_AGEMA_signal_14976, mcs1_mcs_mat1_1_mcs_out[67]}), .b ({new_AGEMA_signal_11607, new_AGEMA_signal_11606, mcs1_mcs_mat1_1_mcs_out[71]}), .c ({new_AGEMA_signal_15537, new_AGEMA_signal_15536, mcs1_mcs_mat1_1_n86}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U30 ( .a ({new_AGEMA_signal_14963, new_AGEMA_signal_14962, mcs1_mcs_mat1_1_n84}), .b ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, mcs1_mcs_mat1_1_n83}), .c ({new_AGEMA_signal_15539, new_AGEMA_signal_15538, mcs_out[154]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U29 ( .a ({new_AGEMA_signal_12499, new_AGEMA_signal_12498, mcs1_mcs_mat1_1_mcs_out[74]}), .b ({new_AGEMA_signal_8243, new_AGEMA_signal_8242, mcs1_mcs_mat1_1_mcs_out[78]}), .c ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, mcs1_mcs_mat1_1_n83}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U28 ( .a ({new_AGEMA_signal_14489, new_AGEMA_signal_14488, mcs1_mcs_mat1_1_mcs_out[66]}), .b ({new_AGEMA_signal_12503, new_AGEMA_signal_12502, mcs1_mcs_mat1_1_mcs_out[70]}), .c ({new_AGEMA_signal_14963, new_AGEMA_signal_14962, mcs1_mcs_mat1_1_n84}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U27 ( .a ({new_AGEMA_signal_14037, new_AGEMA_signal_14036, mcs1_mcs_mat1_1_n82}), .b ({new_AGEMA_signal_11551, new_AGEMA_signal_11550, mcs1_mcs_mat1_1_n81}), .c ({new_AGEMA_signal_14473, new_AGEMA_signal_14472, mcs_out[153]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U26 ( .a ({new_AGEMA_signal_10633, new_AGEMA_signal_10632, mcs1_mcs_mat1_1_mcs_out[73]}), .b ({new_AGEMA_signal_9671, new_AGEMA_signal_9670, mcs1_mcs_mat1_1_mcs_out[77]}), .c ({new_AGEMA_signal_11551, new_AGEMA_signal_11550, mcs1_mcs_mat1_1_n81}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U25 ( .a ({new_AGEMA_signal_13583, new_AGEMA_signal_13582, mcs1_mcs_mat1_1_mcs_out[65]}), .b ({new_AGEMA_signal_12505, new_AGEMA_signal_12504, mcs1_mcs_mat1_1_mcs_out[69]}), .c ({new_AGEMA_signal_14037, new_AGEMA_signal_14036, mcs1_mcs_mat1_1_n82}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U24 ( .a ({new_AGEMA_signal_16031, new_AGEMA_signal_16030, mcs1_mcs_mat1_1_n80}), .b ({new_AGEMA_signal_13079, new_AGEMA_signal_13078, mcs1_mcs_mat1_1_n79}), .c ({new_AGEMA_signal_16365, new_AGEMA_signal_16364, mcs_out[152]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U23 ( .a ({new_AGEMA_signal_12501, new_AGEMA_signal_12500, mcs1_mcs_mat1_1_mcs_out[72]}), .b ({new_AGEMA_signal_12497, new_AGEMA_signal_12496, mcs1_mcs_mat1_1_mcs_out[76]}), .c ({new_AGEMA_signal_13079, new_AGEMA_signal_13078, mcs1_mcs_mat1_1_n79}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U22 ( .a ({new_AGEMA_signal_15547, new_AGEMA_signal_15546, mcs1_mcs_mat1_1_mcs_out[64]}), .b ({new_AGEMA_signal_11611, new_AGEMA_signal_11610, mcs1_mcs_mat1_1_mcs_out[68]}), .c ({new_AGEMA_signal_16031, new_AGEMA_signal_16030, mcs1_mcs_mat1_1_n80}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U21 ( .a ({new_AGEMA_signal_14039, new_AGEMA_signal_14038, mcs1_mcs_mat1_1_n78}), .b ({new_AGEMA_signal_12471, new_AGEMA_signal_12470, mcs1_mcs_mat1_1_n77}), .c ({temp_next_s2[123], temp_next_s1[123], temp_next_s0[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U20 ( .a ({new_AGEMA_signal_10649, new_AGEMA_signal_10648, mcs1_mcs_mat1_1_mcs_out[59]}), .b ({new_AGEMA_signal_11615, new_AGEMA_signal_11614, mcs1_mcs_mat1_1_mcs_out[63]}), .c ({new_AGEMA_signal_12471, new_AGEMA_signal_12470, mcs1_mcs_mat1_1_n77}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U19 ( .a ({new_AGEMA_signal_13587, new_AGEMA_signal_13586, mcs1_mcs_mat1_1_mcs_out[51]}), .b ({new_AGEMA_signal_11621, new_AGEMA_signal_11620, mcs1_mcs_mat1_1_mcs_out[55]}), .c ({new_AGEMA_signal_14039, new_AGEMA_signal_14038, mcs1_mcs_mat1_1_n78}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U18 ( .a ({new_AGEMA_signal_13081, new_AGEMA_signal_13080, mcs1_mcs_mat1_1_n76}), .b ({new_AGEMA_signal_11553, new_AGEMA_signal_11552, mcs1_mcs_mat1_1_n75}), .c ({temp_next_s2[122], temp_next_s1[122], temp_next_s0[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U17 ( .a ({new_AGEMA_signal_9691, new_AGEMA_signal_9690, mcs1_mcs_mat1_1_mcs_out[58]}), .b ({new_AGEMA_signal_10643, new_AGEMA_signal_10642, mcs1_mcs_mat1_1_mcs_out[62]}), .c ({new_AGEMA_signal_11553, new_AGEMA_signal_11552, mcs1_mcs_mat1_1_n75}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U16 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_12509, new_AGEMA_signal_12508, mcs1_mcs_mat1_1_mcs_out[54]}), .c ({new_AGEMA_signal_13081, new_AGEMA_signal_13080, mcs1_mcs_mat1_1_n76}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U15 ( .a ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, mcs1_mcs_mat1_1_n74}), .b ({new_AGEMA_signal_11555, new_AGEMA_signal_11554, mcs1_mcs_mat1_1_n73}), .c ({temp_next_s2[121], temp_next_s1[121], temp_next_s0[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U14 ( .a ({new_AGEMA_signal_10651, new_AGEMA_signal_10650, mcs1_mcs_mat1_1_mcs_out[57]}), .b ({new_AGEMA_signal_10645, new_AGEMA_signal_10644, mcs1_mcs_mat1_1_mcs_out[61]}), .c ({new_AGEMA_signal_11555, new_AGEMA_signal_11554, mcs1_mcs_mat1_1_n73}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U13 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_12511, new_AGEMA_signal_12510, mcs1_mcs_mat1_1_mcs_out[53]}), .c ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, mcs1_mcs_mat1_1_n74}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U12 ( .a ({new_AGEMA_signal_14477, new_AGEMA_signal_14476, mcs1_mcs_mat1_1_n72}), .b ({new_AGEMA_signal_13085, new_AGEMA_signal_13084, mcs1_mcs_mat1_1_n71}), .c ({temp_next_s2[120], temp_next_s1[120], temp_next_s0[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U11 ( .a ({new_AGEMA_signal_11619, new_AGEMA_signal_11618, mcs1_mcs_mat1_1_mcs_out[56]}), .b ({new_AGEMA_signal_12507, new_AGEMA_signal_12506, mcs1_mcs_mat1_1_mcs_out[60]}), .c ({new_AGEMA_signal_13085, new_AGEMA_signal_13084, mcs1_mcs_mat1_1_n71}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U10 ( .a ({new_AGEMA_signal_14061, new_AGEMA_signal_14060, mcs1_mcs_mat1_1_mcs_out[48]}), .b ({new_AGEMA_signal_11625, new_AGEMA_signal_11624, mcs1_mcs_mat1_1_mcs_out[52]}), .c ({new_AGEMA_signal_14477, new_AGEMA_signal_14476, mcs1_mcs_mat1_1_n72}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U9 ( .a ({new_AGEMA_signal_14967, new_AGEMA_signal_14966, mcs1_mcs_mat1_1_n70}), .b ({new_AGEMA_signal_12473, new_AGEMA_signal_12472, mcs1_mcs_mat1_1_n69}), .c ({temp_next_s2[91], temp_next_s1[91], temp_next_s0[91]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U8 ( .a ({new_AGEMA_signal_11629, new_AGEMA_signal_11628, mcs1_mcs_mat1_1_mcs_out[43]}), .b ({new_AGEMA_signal_11627, new_AGEMA_signal_11626, mcs1_mcs_mat1_1_mcs_out[47]}), .c ({new_AGEMA_signal_12473, new_AGEMA_signal_12472, mcs1_mcs_mat1_1_n69}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U7 ( .a ({new_AGEMA_signal_14493, new_AGEMA_signal_14492, mcs1_mcs_mat1_1_mcs_out[35]}), .b ({new_AGEMA_signal_12515, new_AGEMA_signal_12514, mcs1_mcs_mat1_1_mcs_out[39]}), .c ({new_AGEMA_signal_14967, new_AGEMA_signal_14966, mcs1_mcs_mat1_1_n70}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U6 ( .a ({new_AGEMA_signal_14479, new_AGEMA_signal_14478, mcs1_mcs_mat1_1_n68}), .b ({new_AGEMA_signal_12475, new_AGEMA_signal_12474, mcs1_mcs_mat1_1_n67}), .c ({temp_next_s2[90], temp_next_s1[90], temp_next_s0[90]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U5 ( .a ({new_AGEMA_signal_11631, new_AGEMA_signal_11630, mcs1_mcs_mat1_1_mcs_out[42]}), .b ({new_AGEMA_signal_9015, new_AGEMA_signal_9014, mcs1_mcs_mat1_1_mcs_out[46]}), .c ({new_AGEMA_signal_12475, new_AGEMA_signal_12474, mcs1_mcs_mat1_1_n67}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U4 ( .a ({new_AGEMA_signal_14063, new_AGEMA_signal_14062, mcs1_mcs_mat1_1_mcs_out[34]}), .b ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, mcs1_mcs_mat1_1_mcs_out[38]}), .c ({new_AGEMA_signal_14479, new_AGEMA_signal_14478, mcs1_mcs_mat1_1_n68}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U3 ( .a ({new_AGEMA_signal_14971, new_AGEMA_signal_14970, mcs1_mcs_mat1_1_n66}), .b ({new_AGEMA_signal_14041, new_AGEMA_signal_14040, mcs1_mcs_mat1_1_n65}), .c ({temp_next_s2[24], temp_next_s1[24], temp_next_s0[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U2 ( .a ({new_AGEMA_signal_13601, new_AGEMA_signal_13600, mcs1_mcs_mat1_1_mcs_out[4]}), .b ({new_AGEMA_signal_12533, new_AGEMA_signal_12532, mcs1_mcs_mat1_1_mcs_out[8]}), .c ({new_AGEMA_signal_14041, new_AGEMA_signal_14040, mcs1_mcs_mat1_1_n65}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_U1 ( .a ({new_AGEMA_signal_14501, new_AGEMA_signal_14500, mcs1_mcs_mat1_1_mcs_out[0]}), .b ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, mcs1_mcs_mat1_1_mcs_out[12]}), .c ({new_AGEMA_signal_14971, new_AGEMA_signal_14970, mcs1_mcs_mat1_1_n66}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_11557, new_AGEMA_signal_11556, mcs1_mcs_mat1_1_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_12477, new_AGEMA_signal_12476, mcs1_mcs_mat1_1_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_10599, new_AGEMA_signal_10598, mcs1_mcs_mat1_1_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_7711, new_AGEMA_signal_7710, mcs1_mcs_mat1_1_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_11557, new_AGEMA_signal_11556, mcs1_mcs_mat1_1_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_8229, new_AGEMA_signal_8228, mcs1_mcs_mat1_1_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_8971, new_AGEMA_signal_8970, mcs1_mcs_mat1_1_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_9637, new_AGEMA_signal_9636, mcs1_mcs_mat1_1_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_8231, new_AGEMA_signal_8230, mcs1_mcs_mat1_1_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .c ({new_AGEMA_signal_8971, new_AGEMA_signal_8970, mcs1_mcs_mat1_1_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_11559, new_AGEMA_signal_11558, mcs1_mcs_mat1_1_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .c ({new_AGEMA_signal_12479, new_AGEMA_signal_12478, mcs1_mcs_mat1_1_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_10599, new_AGEMA_signal_10598, mcs1_mcs_mat1_1_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_11559, new_AGEMA_signal_11558, mcs1_mcs_mat1_1_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, mcs1_mcs_mat1_1_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_8973, new_AGEMA_signal_8972, mcs1_mcs_mat1_1_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_10599, new_AGEMA_signal_10598, mcs1_mcs_mat1_1_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_10601, new_AGEMA_signal_10600, mcs1_mcs_mat1_1_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_11561, new_AGEMA_signal_11560, mcs1_mcs_mat1_1_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, mcs1_mcs_mat1_1_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_8231, new_AGEMA_signal_8230, mcs1_mcs_mat1_1_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_10601, new_AGEMA_signal_10600, mcs1_mcs_mat1_1_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, mcs1_mcs_mat1_1_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1601], Fresh[1600], Fresh[1599]}), .c ({new_AGEMA_signal_8231, new_AGEMA_signal_8230, mcs1_mcs_mat1_1_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({new_AGEMA_signal_8973, new_AGEMA_signal_8972, mcs1_mcs_mat1_1_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_11563, new_AGEMA_signal_11562, mcs1_mcs_mat1_1_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .c ({new_AGEMA_signal_12481, new_AGEMA_signal_12480, mcs1_mcs_mat1_1_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_10603, new_AGEMA_signal_10602, mcs1_mcs_mat1_1_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_8979, new_AGEMA_signal_8978, mcs1_mcs_mat1_1_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_11563, new_AGEMA_signal_11562, mcs1_mcs_mat1_1_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_11565, new_AGEMA_signal_11564, mcs1_mcs_mat1_1_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_9643, new_AGEMA_signal_9642, mcs1_mcs_mat1_1_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_12483, new_AGEMA_signal_12482, mcs1_mcs_mat1_1_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_10603, new_AGEMA_signal_10602, mcs1_mcs_mat1_1_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .c ({new_AGEMA_signal_11565, new_AGEMA_signal_11564, mcs1_mcs_mat1_1_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_10603, new_AGEMA_signal_10602, mcs1_mcs_mat1_1_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9641, new_AGEMA_signal_9640, mcs1_mcs_mat1_1_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_11567, new_AGEMA_signal_11566, mcs1_mcs_mat1_1_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, mcs1_mcs_mat1_1_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_8233, new_AGEMA_signal_8232, mcs1_mcs_mat1_1_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_10603, new_AGEMA_signal_10602, mcs1_mcs_mat1_1_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_8977, new_AGEMA_signal_8976, mcs1_mcs_mat1_1_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_9643, new_AGEMA_signal_9642, mcs1_mcs_mat1_1_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_10605, new_AGEMA_signal_10604, mcs1_mcs_mat1_1_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_7713, new_AGEMA_signal_7712, mcs1_mcs_mat1_1_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_8979, new_AGEMA_signal_8978, mcs1_mcs_mat1_1_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_9643, new_AGEMA_signal_9642, mcs1_mcs_mat1_1_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_8233, new_AGEMA_signal_8232, mcs1_mcs_mat1_1_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_8977, new_AGEMA_signal_8976, mcs1_mcs_mat1_1_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1607], Fresh[1606], Fresh[1605]}), .c ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, mcs1_mcs_mat1_1_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_8233, new_AGEMA_signal_8232, mcs1_mcs_mat1_1_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1613], Fresh[1612], Fresh[1611]}), .c ({new_AGEMA_signal_8979, new_AGEMA_signal_8978, mcs1_mcs_mat1_1_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_14045, new_AGEMA_signal_14044, mcs1_mcs_mat1_1_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_11569, new_AGEMA_signal_11568, mcs1_mcs_mat1_1_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_14481, new_AGEMA_signal_14480, mcs1_mcs_mat1_1_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_13087, new_AGEMA_signal_13086, mcs1_mcs_mat1_1_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, mcs1_mcs_mat1_1_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_13567, new_AGEMA_signal_13566, mcs1_mcs_mat1_1_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_14047, new_AGEMA_signal_14046, mcs1_mcs_mat1_1_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_14483, new_AGEMA_signal_14482, mcs1_mcs_mat1_1_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_14973, new_AGEMA_signal_14972, mcs1_mcs_mat1_1_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_14045, new_AGEMA_signal_14044, mcs1_mcs_mat1_1_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_14483, new_AGEMA_signal_14482, mcs1_mcs_mat1_1_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_10607, new_AGEMA_signal_10606, mcs1_mcs_mat1_1_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_13571, new_AGEMA_signal_13570, mcs1_mcs_mat1_1_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_14045, new_AGEMA_signal_14044, mcs1_mcs_mat1_1_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_11571, new_AGEMA_signal_11570, mcs1_mcs_mat1_1_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_13569, new_AGEMA_signal_13568, mcs1_mcs_mat1_1_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_14047, new_AGEMA_signal_14046, mcs1_mcs_mat1_1_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({new_AGEMA_signal_13571, new_AGEMA_signal_13570, mcs1_mcs_mat1_1_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1619], Fresh[1618], Fresh[1617]}), .c ({new_AGEMA_signal_11571, new_AGEMA_signal_11570, mcs1_mcs_mat1_1_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, mcs1_mcs_mat1_1_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({new_AGEMA_signal_11573, new_AGEMA_signal_11572, mcs1_mcs_mat1_1_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12485, new_AGEMA_signal_12484, mcs1_mcs_mat1_1_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({new_AGEMA_signal_11575, new_AGEMA_signal_11574, mcs1_mcs_mat1_1_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12487, new_AGEMA_signal_12486, mcs1_mcs_mat1_1_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_8981, new_AGEMA_signal_8980, mcs1_mcs_mat1_1_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_11573, new_AGEMA_signal_11572, mcs1_mcs_mat1_1_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12489, new_AGEMA_signal_12488, mcs1_mcs_mat1_1_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_8235, new_AGEMA_signal_8234, mcs1_mcs_mat1_1_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_10609, new_AGEMA_signal_10608, mcs1_mcs_mat1_1_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_11573, new_AGEMA_signal_11572, mcs1_mcs_mat1_1_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_9647, new_AGEMA_signal_9646, mcs1_mcs_mat1_1_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_11575, new_AGEMA_signal_11574, mcs1_mcs_mat1_1_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12491, new_AGEMA_signal_12490, mcs1_mcs_mat1_1_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_10611, new_AGEMA_signal_10610, mcs1_mcs_mat1_1_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_11575, new_AGEMA_signal_11574, mcs1_mcs_mat1_1_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_8981, new_AGEMA_signal_8980, mcs1_mcs_mat1_1_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_9649, new_AGEMA_signal_9648, mcs1_mcs_mat1_1_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_10611, new_AGEMA_signal_10610, mcs1_mcs_mat1_1_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1625], Fresh[1624], Fresh[1623]}), .c ({new_AGEMA_signal_9649, new_AGEMA_signal_9648, mcs1_mcs_mat1_1_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({new_AGEMA_signal_8235, new_AGEMA_signal_8234, mcs1_mcs_mat1_1_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1631], Fresh[1630], Fresh[1629]}), .c ({new_AGEMA_signal_8981, new_AGEMA_signal_8980, mcs1_mcs_mat1_1_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_10615, new_AGEMA_signal_10614, mcs1_mcs_mat1_1_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_10613, new_AGEMA_signal_10612, mcs1_mcs_mat1_1_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_11577, new_AGEMA_signal_11576, mcs1_mcs_mat1_1_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_10613, new_AGEMA_signal_10612, mcs1_mcs_mat1_1_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_8983, new_AGEMA_signal_8982, mcs1_mcs_mat1_1_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_11579, new_AGEMA_signal_11578, mcs1_mcs_mat1_1_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_8237, new_AGEMA_signal_8236, mcs1_mcs_mat1_1_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .c ({new_AGEMA_signal_8983, new_AGEMA_signal_8982, mcs1_mcs_mat1_1_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_10613, new_AGEMA_signal_10612, mcs1_mcs_mat1_1_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_11581, new_AGEMA_signal_11580, mcs1_mcs_mat1_1_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_9653, new_AGEMA_signal_9652, mcs1_mcs_mat1_1_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_7717, new_AGEMA_signal_7716, mcs1_mcs_mat1_1_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_10613, new_AGEMA_signal_10612, mcs1_mcs_mat1_1_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_11583, new_AGEMA_signal_11582, mcs1_mcs_mat1_1_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_12493, new_AGEMA_signal_12492, mcs1_mcs_mat1_1_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_10615, new_AGEMA_signal_10614, mcs1_mcs_mat1_1_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_9653, new_AGEMA_signal_9652, mcs1_mcs_mat1_1_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_11583, new_AGEMA_signal_11582, mcs1_mcs_mat1_1_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, mcs1_mcs_mat1_1_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .c ({new_AGEMA_signal_10615, new_AGEMA_signal_10614, mcs1_mcs_mat1_1_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_8237, new_AGEMA_signal_8236, mcs1_mcs_mat1_1_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_8985, new_AGEMA_signal_8984, mcs1_mcs_mat1_1_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, mcs1_mcs_mat1_1_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({new_AGEMA_signal_9653, new_AGEMA_signal_9652, mcs1_mcs_mat1_1_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1637], Fresh[1636], Fresh[1635]}), .c ({new_AGEMA_signal_8237, new_AGEMA_signal_8236, mcs1_mcs_mat1_1_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({new_AGEMA_signal_8985, new_AGEMA_signal_8984, mcs1_mcs_mat1_1_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_8987, new_AGEMA_signal_8986, mcs1_mcs_mat1_1_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_10617, new_AGEMA_signal_10616, mcs1_mcs_mat1_1_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_11585, new_AGEMA_signal_11584, mcs1_mcs_mat1_1_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_9661, new_AGEMA_signal_9660, mcs1_mcs_mat1_1_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_10617, new_AGEMA_signal_10616, mcs1_mcs_mat1_1_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, mcs1_mcs_mat1_1_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_8989, new_AGEMA_signal_8988, mcs1_mcs_mat1_1_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_10619, new_AGEMA_signal_10618, mcs1_mcs_mat1_1_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_9659, new_AGEMA_signal_9658, mcs1_mcs_mat1_1_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_10621, new_AGEMA_signal_10620, mcs1_mcs_mat1_1_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_11587, new_AGEMA_signal_11586, mcs1_mcs_mat1_1_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, mcs1_mcs_mat1_1_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_9661, new_AGEMA_signal_9660, mcs1_mcs_mat1_1_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_10621, new_AGEMA_signal_10620, mcs1_mcs_mat1_1_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_8239, new_AGEMA_signal_8238, mcs1_mcs_mat1_1_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .c ({new_AGEMA_signal_9659, new_AGEMA_signal_9658, mcs1_mcs_mat1_1_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1643], Fresh[1642], Fresh[1641]}), .c ({new_AGEMA_signal_9661, new_AGEMA_signal_9660, mcs1_mcs_mat1_1_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({new_AGEMA_signal_8239, new_AGEMA_signal_8238, mcs1_mcs_mat1_1_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1649], Fresh[1648], Fresh[1647]}), .c ({new_AGEMA_signal_8989, new_AGEMA_signal_8988, mcs1_mcs_mat1_1_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_15545, new_AGEMA_signal_15544, mcs1_mcs_mat1_1_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_13093, new_AGEMA_signal_13092, mcs1_mcs_mat1_1_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_16033, new_AGEMA_signal_16032, mcs1_mcs_mat1_1_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_14975, new_AGEMA_signal_14974, mcs1_mcs_mat1_1_mcs_out[99]}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .c ({new_AGEMA_signal_15545, new_AGEMA_signal_15544, mcs1_mcs_mat1_1_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_14485, new_AGEMA_signal_14484, mcs1_mcs_mat1_1_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .c ({new_AGEMA_signal_14975, new_AGEMA_signal_14974, mcs1_mcs_mat1_1_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_14049, new_AGEMA_signal_14048, mcs1_mcs_mat1_1_mcs_out[98]}), .b ({new_AGEMA_signal_11591, new_AGEMA_signal_11590, mcs1_mcs_mat1_1_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_14485, new_AGEMA_signal_14484, mcs1_mcs_mat1_1_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_11589, new_AGEMA_signal_11588, mcs1_mcs_mat1_1_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_13573, new_AGEMA_signal_13572, mcs1_mcs_mat1_1_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_14049, new_AGEMA_signal_14048, mcs1_mcs_mat1_1_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({new_AGEMA_signal_13573, new_AGEMA_signal_13572, mcs1_mcs_mat1_1_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1655], Fresh[1654], Fresh[1653]}), .c ({new_AGEMA_signal_11591, new_AGEMA_signal_11590, mcs1_mcs_mat1_1_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({new_AGEMA_signal_13093, new_AGEMA_signal_13092, mcs1_mcs_mat1_1_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_10625, new_AGEMA_signal_10624, mcs1_mcs_mat1_1_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_11593, new_AGEMA_signal_11592, mcs1_mcs_mat1_1_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_8993, new_AGEMA_signal_8992, mcs1_mcs_mat1_1_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_8995, new_AGEMA_signal_8994, mcs1_mcs_mat1_1_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_9665, new_AGEMA_signal_9664, mcs1_mcs_mat1_1_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_11595, new_AGEMA_signal_11594, mcs1_mcs_mat1_1_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_8241, new_AGEMA_signal_8240, mcs1_mcs_mat1_1_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_12495, new_AGEMA_signal_12494, mcs1_mcs_mat1_1_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_10625, new_AGEMA_signal_10624, mcs1_mcs_mat1_1_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_11595, new_AGEMA_signal_11594, mcs1_mcs_mat1_1_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_7721, new_AGEMA_signal_7720, mcs1_mcs_mat1_1_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_9667, new_AGEMA_signal_9666, mcs1_mcs_mat1_1_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_10625, new_AGEMA_signal_10624, mcs1_mcs_mat1_1_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1661], Fresh[1660], Fresh[1659]}), .c ({new_AGEMA_signal_9667, new_AGEMA_signal_9666, mcs1_mcs_mat1_1_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({new_AGEMA_signal_8241, new_AGEMA_signal_8240, mcs1_mcs_mat1_1_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1667], Fresh[1666], Fresh[1665]}), .c ({new_AGEMA_signal_8995, new_AGEMA_signal_8994, mcs1_mcs_mat1_1_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_13579, new_AGEMA_signal_13578, mcs1_mcs_mat1_1_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_13581, new_AGEMA_signal_13580, mcs1_mcs_mat1_1_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_14051, new_AGEMA_signal_14050, mcs1_mcs_mat1_1_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_13575, new_AGEMA_signal_13574, mcs1_mcs_mat1_1_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_10629, new_AGEMA_signal_10628, mcs1_mcs_mat1_1_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_14053, new_AGEMA_signal_14052, mcs1_mcs_mat1_1_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, mcs1_mcs_mat1_1_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_13575, new_AGEMA_signal_13574, mcs1_mcs_mat1_1_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_13577, new_AGEMA_signal_13576, mcs1_mcs_mat1_1_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_14055, new_AGEMA_signal_14054, mcs1_mcs_mat1_1_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_11597, new_AGEMA_signal_11596, mcs1_mcs_mat1_1_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, mcs1_mcs_mat1_1_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_13577, new_AGEMA_signal_13576, mcs1_mcs_mat1_1_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_14057, new_AGEMA_signal_14056, mcs1_mcs_mat1_1_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .c ({new_AGEMA_signal_14487, new_AGEMA_signal_14486, mcs1_mcs_mat1_1_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_13579, new_AGEMA_signal_13578, mcs1_mcs_mat1_1_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_11597, new_AGEMA_signal_11596, mcs1_mcs_mat1_1_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_14057, new_AGEMA_signal_14056, mcs1_mcs_mat1_1_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({new_AGEMA_signal_13581, new_AGEMA_signal_13580, mcs1_mcs_mat1_1_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1673], Fresh[1672], Fresh[1671]}), .c ({new_AGEMA_signal_11597, new_AGEMA_signal_11596, mcs1_mcs_mat1_1_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, mcs1_mcs_mat1_1_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_10631, new_AGEMA_signal_10630, mcs1_mcs_mat1_1_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_11599, new_AGEMA_signal_11598, mcs1_mcs_mat1_1_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_9001, new_AGEMA_signal_9000, mcs1_mcs_mat1_1_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_9671, new_AGEMA_signal_9670, mcs1_mcs_mat1_1_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_11601, new_AGEMA_signal_11600, mcs1_mcs_mat1_1_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_8245, new_AGEMA_signal_8244, mcs1_mcs_mat1_1_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_12497, new_AGEMA_signal_12496, mcs1_mcs_mat1_1_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_10631, new_AGEMA_signal_10630, mcs1_mcs_mat1_1_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .c ({new_AGEMA_signal_11601, new_AGEMA_signal_11600, mcs1_mcs_mat1_1_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_7723, new_AGEMA_signal_7722, mcs1_mcs_mat1_1_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_9673, new_AGEMA_signal_9672, mcs1_mcs_mat1_1_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_10631, new_AGEMA_signal_10630, mcs1_mcs_mat1_1_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1679], Fresh[1678], Fresh[1677]}), .c ({new_AGEMA_signal_9673, new_AGEMA_signal_9672, mcs1_mcs_mat1_1_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({new_AGEMA_signal_8245, new_AGEMA_signal_8244, mcs1_mcs_mat1_1_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1685], Fresh[1684], Fresh[1683]}), .c ({new_AGEMA_signal_9001, new_AGEMA_signal_9000, mcs1_mcs_mat1_1_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_11603, new_AGEMA_signal_11602, mcs1_mcs_mat1_1_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_12499, new_AGEMA_signal_12498, mcs1_mcs_mat1_1_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_10635, new_AGEMA_signal_10634, mcs1_mcs_mat1_1_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9677, new_AGEMA_signal_9676, mcs1_mcs_mat1_1_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_11603, new_AGEMA_signal_11602, mcs1_mcs_mat1_1_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_8769, new_AGEMA_signal_8768, mcs1_mcs_mat1_1_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, mcs1_mcs_mat1_1_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_9677, new_AGEMA_signal_9676, mcs1_mcs_mat1_1_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_8769, new_AGEMA_signal_8768, mcs1_mcs_mat1_1_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_10633, new_AGEMA_signal_10632, mcs1_mcs_mat1_1_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_8247, new_AGEMA_signal_8246, mcs1_mcs_mat1_1_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_8249, new_AGEMA_signal_8248, mcs1_mcs_mat1_1_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_8769, new_AGEMA_signal_8768, mcs1_mcs_mat1_1_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_9003, new_AGEMA_signal_9002, mcs1_mcs_mat1_1_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .c ({new_AGEMA_signal_9677, new_AGEMA_signal_9676, mcs1_mcs_mat1_1_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_11605, new_AGEMA_signal_11604, mcs1_mcs_mat1_1_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_8247, new_AGEMA_signal_8246, mcs1_mcs_mat1_1_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_12501, new_AGEMA_signal_12500, mcs1_mcs_mat1_1_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_10635, new_AGEMA_signal_10634, mcs1_mcs_mat1_1_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9003, new_AGEMA_signal_9002, mcs1_mcs_mat1_1_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_11605, new_AGEMA_signal_11604, mcs1_mcs_mat1_1_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .b ({new_AGEMA_signal_9679, new_AGEMA_signal_9678, mcs1_mcs_mat1_1_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_10635, new_AGEMA_signal_10634, mcs1_mcs_mat1_1_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({new_AGEMA_signal_9679, new_AGEMA_signal_9678, mcs1_mcs_mat1_1_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1691], Fresh[1690], Fresh[1689]}), .c ({new_AGEMA_signal_8249, new_AGEMA_signal_8248, mcs1_mcs_mat1_1_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({new_AGEMA_signal_9003, new_AGEMA_signal_9002, mcs1_mcs_mat1_1_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_10637, new_AGEMA_signal_10636, mcs1_mcs_mat1_1_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_9005, new_AGEMA_signal_9004, mcs1_mcs_mat1_1_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_11607, new_AGEMA_signal_11606, mcs1_mcs_mat1_1_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_9683, new_AGEMA_signal_9682, mcs1_mcs_mat1_1_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_11609, new_AGEMA_signal_11608, mcs1_mcs_mat1_1_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12503, new_AGEMA_signal_12502, mcs1_mcs_mat1_1_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_10637, new_AGEMA_signal_10636, mcs1_mcs_mat1_1_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_11609, new_AGEMA_signal_11608, mcs1_mcs_mat1_1_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12505, new_AGEMA_signal_12504, mcs1_mcs_mat1_1_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_9005, new_AGEMA_signal_9004, mcs1_mcs_mat1_1_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_10639, new_AGEMA_signal_10638, mcs1_mcs_mat1_1_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_11609, new_AGEMA_signal_11608, mcs1_mcs_mat1_1_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({new_AGEMA_signal_8251, new_AGEMA_signal_8250, mcs1_mcs_mat1_1_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_9005, new_AGEMA_signal_9004, mcs1_mcs_mat1_1_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, mcs1_mcs_mat1_1_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .c ({new_AGEMA_signal_10637, new_AGEMA_signal_10636, mcs1_mcs_mat1_1_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_9007, new_AGEMA_signal_9006, mcs1_mcs_mat1_1_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7727, new_AGEMA_signal_7726, mcs1_mcs_mat1_1_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, mcs1_mcs_mat1_1_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_10639, new_AGEMA_signal_10638, mcs1_mcs_mat1_1_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_9683, new_AGEMA_signal_9682, mcs1_mcs_mat1_1_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_11611, new_AGEMA_signal_11610, mcs1_mcs_mat1_1_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_9007, new_AGEMA_signal_9006, mcs1_mcs_mat1_1_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_9683, new_AGEMA_signal_9682, mcs1_mcs_mat1_1_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({new_AGEMA_signal_9685, new_AGEMA_signal_9684, mcs1_mcs_mat1_1_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_10639, new_AGEMA_signal_10638, mcs1_mcs_mat1_1_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1697], Fresh[1696], Fresh[1695]}), .c ({new_AGEMA_signal_9685, new_AGEMA_signal_9684, mcs1_mcs_mat1_1_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({new_AGEMA_signal_8251, new_AGEMA_signal_8250, mcs1_mcs_mat1_1_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1703], Fresh[1702], Fresh[1701]}), .c ({new_AGEMA_signal_9007, new_AGEMA_signal_9006, mcs1_mcs_mat1_1_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_14491, new_AGEMA_signal_14490, mcs1_mcs_mat1_1_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_14977, new_AGEMA_signal_14976, mcs1_mcs_mat1_1_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({new_AGEMA_signal_14059, new_AGEMA_signal_14058, mcs1_mcs_mat1_1_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_14489, new_AGEMA_signal_14488, mcs1_mcs_mat1_1_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_14979, new_AGEMA_signal_14978, mcs1_mcs_mat1_1_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_13097, new_AGEMA_signal_13096, mcs1_mcs_mat1_1_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_15547, new_AGEMA_signal_15546, mcs1_mcs_mat1_1_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_14491, new_AGEMA_signal_14490, mcs1_mcs_mat1_1_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .c ({new_AGEMA_signal_14979, new_AGEMA_signal_14978, mcs1_mcs_mat1_1_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_11613, new_AGEMA_signal_11612, mcs1_mcs_mat1_1_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_14059, new_AGEMA_signal_14058, mcs1_mcs_mat1_1_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_14491, new_AGEMA_signal_14490, mcs1_mcs_mat1_1_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_10641, new_AGEMA_signal_10640, mcs1_mcs_mat1_1_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_13585, new_AGEMA_signal_13584, mcs1_mcs_mat1_1_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_14059, new_AGEMA_signal_14058, mcs1_mcs_mat1_1_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({new_AGEMA_signal_13585, new_AGEMA_signal_13584, mcs1_mcs_mat1_1_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1709], Fresh[1708], Fresh[1707]}), .c ({new_AGEMA_signal_11613, new_AGEMA_signal_11612, mcs1_mcs_mat1_1_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({new_AGEMA_signal_13097, new_AGEMA_signal_13096, mcs1_mcs_mat1_1_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_10647, new_AGEMA_signal_10646, mcs1_mcs_mat1_1_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_9009, new_AGEMA_signal_9008, mcs1_mcs_mat1_1_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_11615, new_AGEMA_signal_11614, mcs1_mcs_mat1_1_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_8253, new_AGEMA_signal_8252, mcs1_mcs_mat1_1_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, mcs1_mcs_mat1_1_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_10643, new_AGEMA_signal_10642, mcs1_mcs_mat1_1_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({new_AGEMA_signal_9689, new_AGEMA_signal_9688, mcs1_mcs_mat1_1_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_10645, new_AGEMA_signal_10644, mcs1_mcs_mat1_1_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1715], Fresh[1714], Fresh[1713]}), .c ({new_AGEMA_signal_9689, new_AGEMA_signal_9688, mcs1_mcs_mat1_1_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({new_AGEMA_signal_8253, new_AGEMA_signal_8252, mcs1_mcs_mat1_1_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1721], Fresh[1720], Fresh[1719]}), .c ({new_AGEMA_signal_9009, new_AGEMA_signal_9008, mcs1_mcs_mat1_1_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_8257, new_AGEMA_signal_8256, mcs1_mcs_mat1_1_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_9011, new_AGEMA_signal_9010, mcs1_mcs_mat1_1_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_9691, new_AGEMA_signal_9690, mcs1_mcs_mat1_1_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_8259, new_AGEMA_signal_8258, mcs1_mcs_mat1_1_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, mcs1_mcs_mat1_1_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_10651, new_AGEMA_signal_10650, mcs1_mcs_mat1_1_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_10653, new_AGEMA_signal_10652, mcs1_mcs_mat1_1_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_9695, new_AGEMA_signal_9694, mcs1_mcs_mat1_1_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_11619, new_AGEMA_signal_11618, mcs1_mcs_mat1_1_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_9697, new_AGEMA_signal_9696, mcs1_mcs_mat1_1_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_10653, new_AGEMA_signal_10652, mcs1_mcs_mat1_1_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({new_AGEMA_signal_9697, new_AGEMA_signal_9696, mcs1_mcs_mat1_1_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1727], Fresh[1726], Fresh[1725]}), .c ({new_AGEMA_signal_8259, new_AGEMA_signal_8258, mcs1_mcs_mat1_1_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({new_AGEMA_signal_9011, new_AGEMA_signal_9010, mcs1_mcs_mat1_1_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_9701, new_AGEMA_signal_9700, mcs1_mcs_mat1_1_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_10655, new_AGEMA_signal_10654, mcs1_mcs_mat1_1_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_11621, new_AGEMA_signal_11620, mcs1_mcs_mat1_1_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_11623, new_AGEMA_signal_11622, mcs1_mcs_mat1_1_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, mcs1_mcs_mat1_1_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_12509, new_AGEMA_signal_12508, mcs1_mcs_mat1_1_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_9013, new_AGEMA_signal_9012, mcs1_mcs_mat1_1_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, mcs1_mcs_mat1_1_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({new_AGEMA_signal_11623, new_AGEMA_signal_11622, mcs1_mcs_mat1_1_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_12511, new_AGEMA_signal_12510, mcs1_mcs_mat1_1_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_7733, new_AGEMA_signal_7732, mcs1_mcs_mat1_1_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_10655, new_AGEMA_signal_10654, mcs1_mcs_mat1_1_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_11623, new_AGEMA_signal_11622, mcs1_mcs_mat1_1_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_8261, new_AGEMA_signal_8260, mcs1_mcs_mat1_1_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, mcs1_mcs_mat1_1_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_10655, new_AGEMA_signal_10654, mcs1_mcs_mat1_1_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_9703, new_AGEMA_signal_9702, mcs1_mcs_mat1_1_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_10657, new_AGEMA_signal_10656, mcs1_mcs_mat1_1_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_11625, new_AGEMA_signal_11624, mcs1_mcs_mat1_1_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_9701, new_AGEMA_signal_9700, mcs1_mcs_mat1_1_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8261, new_AGEMA_signal_8260, mcs1_mcs_mat1_1_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_10657, new_AGEMA_signal_10656, mcs1_mcs_mat1_1_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_9013, new_AGEMA_signal_9012, mcs1_mcs_mat1_1_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_9701, new_AGEMA_signal_9700, mcs1_mcs_mat1_1_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1733], Fresh[1732], Fresh[1731]}), .c ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, mcs1_mcs_mat1_1_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({new_AGEMA_signal_8261, new_AGEMA_signal_8260, mcs1_mcs_mat1_1_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1739], Fresh[1738], Fresh[1737]}), .c ({new_AGEMA_signal_9013, new_AGEMA_signal_9012, mcs1_mcs_mat1_1_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_9017, new_AGEMA_signal_9016, mcs1_mcs_mat1_1_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_9707, new_AGEMA_signal_9706, mcs1_mcs_mat1_1_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_12513, new_AGEMA_signal_12512, mcs1_mcs_mat1_1_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_8263, new_AGEMA_signal_8262, mcs1_mcs_mat1_1_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_13099, new_AGEMA_signal_13098, mcs1_mcs_mat1_1_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_11627, new_AGEMA_signal_11626, mcs1_mcs_mat1_1_mcs_out[47]}), .b ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_12513, new_AGEMA_signal_12512, mcs1_mcs_mat1_1_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_10659, new_AGEMA_signal_10658, mcs1_mcs_mat1_1_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .c ({new_AGEMA_signal_11627, new_AGEMA_signal_11626, mcs1_mcs_mat1_1_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_7735, new_AGEMA_signal_7734, mcs1_mcs_mat1_1_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_9709, new_AGEMA_signal_9708, mcs1_mcs_mat1_1_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_10659, new_AGEMA_signal_10658, mcs1_mcs_mat1_1_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({new_AGEMA_signal_9709, new_AGEMA_signal_9708, mcs1_mcs_mat1_1_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1745], Fresh[1744], Fresh[1743]}), .c ({new_AGEMA_signal_8263, new_AGEMA_signal_8262, mcs1_mcs_mat1_1_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({new_AGEMA_signal_9017, new_AGEMA_signal_9016, mcs1_mcs_mat1_1_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_10661, new_AGEMA_signal_10660, mcs1_mcs_mat1_1_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_9019, new_AGEMA_signal_9018, mcs1_mcs_mat1_1_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_11629, new_AGEMA_signal_11628, mcs1_mcs_mat1_1_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, mcs1_mcs_mat1_1_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8265, new_AGEMA_signal_8264, mcs1_mcs_mat1_1_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_10661, new_AGEMA_signal_10660, mcs1_mcs_mat1_1_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_10663, new_AGEMA_signal_10662, mcs1_mcs_mat1_1_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_9715, new_AGEMA_signal_9714, mcs1_mcs_mat1_1_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_11631, new_AGEMA_signal_11630, mcs1_mcs_mat1_1_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_10665, new_AGEMA_signal_10664, mcs1_mcs_mat1_1_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_7737, new_AGEMA_signal_7736, mcs1_mcs_mat1_1_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_11633, new_AGEMA_signal_11632, mcs1_mcs_mat1_1_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, mcs1_mcs_mat1_1_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9021, new_AGEMA_signal_9020, mcs1_mcs_mat1_1_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_10665, new_AGEMA_signal_10664, mcs1_mcs_mat1_1_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_9713, new_AGEMA_signal_9712, mcs1_mcs_mat1_1_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_9021, new_AGEMA_signal_9020, mcs1_mcs_mat1_1_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_10667, new_AGEMA_signal_10666, mcs1_mcs_mat1_1_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1751], Fresh[1750], Fresh[1749]}), .c ({new_AGEMA_signal_9715, new_AGEMA_signal_9714, mcs1_mcs_mat1_1_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({new_AGEMA_signal_8265, new_AGEMA_signal_8264, mcs1_mcs_mat1_1_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1757], Fresh[1756], Fresh[1755]}), .c ({new_AGEMA_signal_9021, new_AGEMA_signal_9020, mcs1_mcs_mat1_1_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_11635, new_AGEMA_signal_11634, mcs1_mcs_mat1_1_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_7739, new_AGEMA_signal_7738, mcs1_mcs_mat1_1_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_12515, new_AGEMA_signal_12514, mcs1_mcs_mat1_1_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_9025, new_AGEMA_signal_9024, mcs1_mcs_mat1_1_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_9023, new_AGEMA_signal_9022, mcs1_mcs_mat1_1_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, mcs1_mcs_mat1_1_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({new_AGEMA_signal_11635, new_AGEMA_signal_11634, mcs1_mcs_mat1_1_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_12517, new_AGEMA_signal_12516, mcs1_mcs_mat1_1_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_9719, new_AGEMA_signal_9718, mcs1_mcs_mat1_1_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_10669, new_AGEMA_signal_10668, mcs1_mcs_mat1_1_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_11635, new_AGEMA_signal_11634, mcs1_mcs_mat1_1_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_9721, new_AGEMA_signal_9720, mcs1_mcs_mat1_1_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9027, new_AGEMA_signal_9026, mcs1_mcs_mat1_1_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_10669, new_AGEMA_signal_10668, mcs1_mcs_mat1_1_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_9721, new_AGEMA_signal_9720, mcs1_mcs_mat1_1_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9025, new_AGEMA_signal_9024, mcs1_mcs_mat1_1_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_10671, new_AGEMA_signal_10670, mcs1_mcs_mat1_1_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_8771, new_AGEMA_signal_8770, mcs1_mcs_mat1_1_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_9025, new_AGEMA_signal_9024, mcs1_mcs_mat1_1_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({new_AGEMA_signal_8267, new_AGEMA_signal_8266, mcs1_mcs_mat1_1_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_8771, new_AGEMA_signal_8770, mcs1_mcs_mat1_1_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({new_AGEMA_signal_9721, new_AGEMA_signal_9720, mcs1_mcs_mat1_1_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1763], Fresh[1762], Fresh[1761]}), .c ({new_AGEMA_signal_8267, new_AGEMA_signal_8266, mcs1_mcs_mat1_1_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({new_AGEMA_signal_9027, new_AGEMA_signal_9026, mcs1_mcs_mat1_1_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_13589, new_AGEMA_signal_13588, mcs1_mcs_mat1_1_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, mcs1_mcs_mat1_1_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_14063, new_AGEMA_signal_14062, mcs1_mcs_mat1_1_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_11637, new_AGEMA_signal_11636, mcs1_mcs_mat1_1_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_12519, new_AGEMA_signal_12518, mcs1_mcs_mat1_1_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_14981, new_AGEMA_signal_14980, mcs1_mcs_mat1_1_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_13591, new_AGEMA_signal_13590, mcs1_mcs_mat1_1_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_15549, new_AGEMA_signal_15548, mcs1_mcs_mat1_1_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1769], Fresh[1768], Fresh[1767]}), .c ({new_AGEMA_signal_13591, new_AGEMA_signal_13590, mcs1_mcs_mat1_1_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({new_AGEMA_signal_11637, new_AGEMA_signal_11636, mcs1_mcs_mat1_1_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1775], Fresh[1774], Fresh[1773]}), .c ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, mcs1_mcs_mat1_1_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_11639, new_AGEMA_signal_11638, mcs1_mcs_mat1_1_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_10675, new_AGEMA_signal_10674, mcs1_mcs_mat1_1_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_12521, new_AGEMA_signal_12520, mcs1_mcs_mat1_1_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_8271, new_AGEMA_signal_8270, mcs1_mcs_mat1_1_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_10677, new_AGEMA_signal_10676, mcs1_mcs_mat1_1_mcs_out[29]}), .c ({new_AGEMA_signal_11639, new_AGEMA_signal_11638, mcs1_mcs_mat1_1_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_8269, new_AGEMA_signal_8268, mcs1_mcs_mat1_1_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_10675, new_AGEMA_signal_10674, mcs1_mcs_mat1_1_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_11641, new_AGEMA_signal_11640, mcs1_mcs_mat1_1_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_9727, new_AGEMA_signal_9726, mcs1_mcs_mat1_1_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .c ({new_AGEMA_signal_10675, new_AGEMA_signal_10674, mcs1_mcs_mat1_1_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_11643, new_AGEMA_signal_11642, mcs1_mcs_mat1_1_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, mcs1_mcs_mat1_1_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_12523, new_AGEMA_signal_12522, mcs1_mcs_mat1_1_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_10679, new_AGEMA_signal_10678, mcs1_mcs_mat1_1_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_9725, new_AGEMA_signal_9724, mcs1_mcs_mat1_1_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_11643, new_AGEMA_signal_11642, mcs1_mcs_mat1_1_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_9029, new_AGEMA_signal_9028, mcs1_mcs_mat1_1_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_9725, new_AGEMA_signal_9724, mcs1_mcs_mat1_1_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_9727, new_AGEMA_signal_9726, mcs1_mcs_mat1_1_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8271, new_AGEMA_signal_8270, mcs1_mcs_mat1_1_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_10679, new_AGEMA_signal_10678, mcs1_mcs_mat1_1_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({new_AGEMA_signal_9727, new_AGEMA_signal_9726, mcs1_mcs_mat1_1_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1781], Fresh[1780], Fresh[1779]}), .c ({new_AGEMA_signal_8271, new_AGEMA_signal_8270, mcs1_mcs_mat1_1_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({new_AGEMA_signal_9029, new_AGEMA_signal_9028, mcs1_mcs_mat1_1_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_9729, new_AGEMA_signal_9728, mcs1_mcs_mat1_1_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_10681, new_AGEMA_signal_10680, mcs1_mcs_mat1_1_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_9031, new_AGEMA_signal_9030, mcs1_mcs_mat1_1_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8273, new_AGEMA_signal_8272, mcs1_mcs_mat1_1_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_9729, new_AGEMA_signal_9728, mcs1_mcs_mat1_1_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_10683, new_AGEMA_signal_10682, mcs1_mcs_mat1_1_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_11645, new_AGEMA_signal_11644, mcs1_mcs_mat1_1_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_9733, new_AGEMA_signal_9732, mcs1_mcs_mat1_1_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8273, new_AGEMA_signal_8272, mcs1_mcs_mat1_1_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_10683, new_AGEMA_signal_10682, mcs1_mcs_mat1_1_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_11647, new_AGEMA_signal_11646, mcs1_mcs_mat1_1_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .c ({new_AGEMA_signal_12525, new_AGEMA_signal_12524, mcs1_mcs_mat1_1_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_9733, new_AGEMA_signal_9732, mcs1_mcs_mat1_1_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_10685, new_AGEMA_signal_10684, mcs1_mcs_mat1_1_mcs_out[24]}), .c ({new_AGEMA_signal_11647, new_AGEMA_signal_11646, mcs1_mcs_mat1_1_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_9731, new_AGEMA_signal_9730, mcs1_mcs_mat1_1_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .c ({new_AGEMA_signal_10685, new_AGEMA_signal_10684, mcs1_mcs_mat1_1_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_9031, new_AGEMA_signal_9030, mcs1_mcs_mat1_1_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7743, new_AGEMA_signal_7742, mcs1_mcs_mat1_1_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_9731, new_AGEMA_signal_9730, mcs1_mcs_mat1_1_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1787], Fresh[1786], Fresh[1785]}), .c ({new_AGEMA_signal_9733, new_AGEMA_signal_9732, mcs1_mcs_mat1_1_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({new_AGEMA_signal_8273, new_AGEMA_signal_8272, mcs1_mcs_mat1_1_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1793], Fresh[1792], Fresh[1791]}), .c ({new_AGEMA_signal_9031, new_AGEMA_signal_9030, mcs1_mcs_mat1_1_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_9735, new_AGEMA_signal_9734, mcs1_mcs_mat1_1_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .c ({new_AGEMA_signal_10687, new_AGEMA_signal_10686, mcs1_mcs_mat1_1_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_9033, new_AGEMA_signal_9032, mcs1_mcs_mat1_1_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8275, new_AGEMA_signal_8274, mcs1_mcs_mat1_1_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_9735, new_AGEMA_signal_9734, mcs1_mcs_mat1_1_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_10689, new_AGEMA_signal_10688, mcs1_mcs_mat1_1_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .c ({new_AGEMA_signal_11649, new_AGEMA_signal_11648, mcs1_mcs_mat1_1_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_9739, new_AGEMA_signal_9738, mcs1_mcs_mat1_1_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8275, new_AGEMA_signal_8274, mcs1_mcs_mat1_1_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_10689, new_AGEMA_signal_10688, mcs1_mcs_mat1_1_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_11651, new_AGEMA_signal_11650, mcs1_mcs_mat1_1_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_7517, new_AGEMA_signal_7516, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_12527, new_AGEMA_signal_12526, mcs1_mcs_mat1_1_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_9739, new_AGEMA_signal_9738, mcs1_mcs_mat1_1_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_10691, new_AGEMA_signal_10690, mcs1_mcs_mat1_1_mcs_out[20]}), .c ({new_AGEMA_signal_11651, new_AGEMA_signal_11650, mcs1_mcs_mat1_1_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_9737, new_AGEMA_signal_9736, mcs1_mcs_mat1_1_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_10691, new_AGEMA_signal_10690, mcs1_mcs_mat1_1_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_9033, new_AGEMA_signal_9032, mcs1_mcs_mat1_1_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7745, new_AGEMA_signal_7744, mcs1_mcs_mat1_1_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_9737, new_AGEMA_signal_9736, mcs1_mcs_mat1_1_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({new_AGEMA_signal_9739, new_AGEMA_signal_9738, mcs1_mcs_mat1_1_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1799], Fresh[1798], Fresh[1797]}), .c ({new_AGEMA_signal_8275, new_AGEMA_signal_8274, mcs1_mcs_mat1_1_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({new_AGEMA_signal_9033, new_AGEMA_signal_9032, mcs1_mcs_mat1_1_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_13593, new_AGEMA_signal_13592, mcs1_mcs_mat1_1_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_13599, new_AGEMA_signal_13598, mcs1_mcs_mat1_1_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_14067, new_AGEMA_signal_14066, mcs1_mcs_mat1_1_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_14069, new_AGEMA_signal_14068, mcs1_mcs_mat1_1_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_10693, new_AGEMA_signal_10692, mcs1_mcs_mat1_1_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_14495, new_AGEMA_signal_14494, mcs1_mcs_mat1_1_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_14497, new_AGEMA_signal_14496, mcs1_mcs_mat1_1_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_11653, new_AGEMA_signal_11652, mcs1_mcs_mat1_1_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_14983, new_AGEMA_signal_14982, mcs1_mcs_mat1_1_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_14069, new_AGEMA_signal_14068, mcs1_mcs_mat1_1_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_14497, new_AGEMA_signal_14496, mcs1_mcs_mat1_1_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_13595, new_AGEMA_signal_13594, mcs1_mcs_mat1_1_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .c ({new_AGEMA_signal_14069, new_AGEMA_signal_14068, mcs1_mcs_mat1_1_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_13103, new_AGEMA_signal_13102, mcs1_mcs_mat1_1_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_13105, new_AGEMA_signal_13104, mcs1_mcs_mat1_1_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_13595, new_AGEMA_signal_13594, mcs1_mcs_mat1_1_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_13597, new_AGEMA_signal_13596, mcs1_mcs_mat1_1_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_11653, new_AGEMA_signal_11652, mcs1_mcs_mat1_1_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_14071, new_AGEMA_signal_14070, mcs1_mcs_mat1_1_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1805], Fresh[1804], Fresh[1803]}), .c ({new_AGEMA_signal_13599, new_AGEMA_signal_13598, mcs1_mcs_mat1_1_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({new_AGEMA_signal_11653, new_AGEMA_signal_11652, mcs1_mcs_mat1_1_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1811], Fresh[1810], Fresh[1809]}), .c ({new_AGEMA_signal_13105, new_AGEMA_signal_13104, mcs1_mcs_mat1_1_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_11659, new_AGEMA_signal_11658, mcs1_mcs_mat1_1_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_8773, new_AGEMA_signal_8772, mcs1_mcs_mat1_1_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_12529, new_AGEMA_signal_12528, mcs1_mcs_mat1_1_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_10699, new_AGEMA_signal_10698, mcs1_mcs_mat1_1_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_10695, new_AGEMA_signal_10694, mcs1_mcs_mat1_1_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_11655, new_AGEMA_signal_11654, mcs1_mcs_mat1_1_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_9743, new_AGEMA_signal_9742, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_8277, new_AGEMA_signal_8276, mcs1_mcs_mat1_1_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_10695, new_AGEMA_signal_10694, mcs1_mcs_mat1_1_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_8773, new_AGEMA_signal_8772, mcs1_mcs_mat1_1_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_10697, new_AGEMA_signal_10696, mcs1_mcs_mat1_1_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_11657, new_AGEMA_signal_11656, mcs1_mcs_mat1_1_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_9741, new_AGEMA_signal_9740, mcs1_mcs_mat1_1_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_9743, new_AGEMA_signal_9742, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_10697, new_AGEMA_signal_10696, mcs1_mcs_mat1_1_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_7747, new_AGEMA_signal_7746, mcs1_mcs_mat1_1_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_8277, new_AGEMA_signal_8276, mcs1_mcs_mat1_1_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8773, new_AGEMA_signal_8772, mcs1_mcs_mat1_1_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, mcs1_mcs_mat1_1_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, mcs1_mcs_mat1_1_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_11659, new_AGEMA_signal_11658, mcs1_mcs_mat1_1_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_9743, new_AGEMA_signal_9742, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, mcs1_mcs_mat1_1_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_10699, new_AGEMA_signal_10698, mcs1_mcs_mat1_1_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_11659, new_AGEMA_signal_11658, mcs1_mcs_mat1_1_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_9741, new_AGEMA_signal_9740, mcs1_mcs_mat1_1_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_10699, new_AGEMA_signal_10698, mcs1_mcs_mat1_1_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, shiftr_out[120]}), .b ({new_AGEMA_signal_9035, new_AGEMA_signal_9034, mcs1_mcs_mat1_1_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_9741, new_AGEMA_signal_9740, mcs1_mcs_mat1_1_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8855, new_AGEMA_signal_8854, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({new_AGEMA_signal_9743, new_AGEMA_signal_9742, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7631, new_AGEMA_signal_7630, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1817], Fresh[1816], Fresh[1815]}), .c ({new_AGEMA_signal_8277, new_AGEMA_signal_8276, mcs1_mcs_mat1_1_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8723, new_AGEMA_signal_8722, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({new_AGEMA_signal_9035, new_AGEMA_signal_9034, mcs1_mcs_mat1_1_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, mcs1_mcs_mat1_1_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .c ({new_AGEMA_signal_9037, new_AGEMA_signal_9036, mcs1_mcs_mat1_1_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_10703, new_AGEMA_signal_10702, mcs1_mcs_mat1_1_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_11661, new_AGEMA_signal_11660, mcs1_mcs_mat1_1_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_9745, new_AGEMA_signal_9744, mcs1_mcs_mat1_1_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_10701, new_AGEMA_signal_10700, mcs1_mcs_mat1_1_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_9039, new_AGEMA_signal_9038, mcs1_mcs_mat1_1_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, mcs1_mcs_mat1_1_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_9745, new_AGEMA_signal_9744, mcs1_mcs_mat1_1_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_7749, new_AGEMA_signal_7748, mcs1_mcs_mat1_1_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8279, new_AGEMA_signal_8278, mcs1_mcs_mat1_1_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, mcs1_mcs_mat1_1_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_11663, new_AGEMA_signal_11662, mcs1_mcs_mat1_1_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_7505, new_AGEMA_signal_7504, shiftr_out[88]}), .c ({new_AGEMA_signal_12533, new_AGEMA_signal_12532, mcs1_mcs_mat1_1_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_7749, new_AGEMA_signal_7748, mcs1_mcs_mat1_1_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_10703, new_AGEMA_signal_10702, mcs1_mcs_mat1_1_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_11663, new_AGEMA_signal_11662, mcs1_mcs_mat1_1_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_9747, new_AGEMA_signal_9746, mcs1_mcs_mat1_1_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_9039, new_AGEMA_signal_9038, mcs1_mcs_mat1_1_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_10703, new_AGEMA_signal_10702, mcs1_mcs_mat1_1_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1823], Fresh[1822], Fresh[1821]}), .c ({new_AGEMA_signal_9747, new_AGEMA_signal_9746, mcs1_mcs_mat1_1_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({new_AGEMA_signal_8279, new_AGEMA_signal_8278, mcs1_mcs_mat1_1_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, shiftr_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1829], Fresh[1828], Fresh[1827]}), .c ({new_AGEMA_signal_9039, new_AGEMA_signal_9038, mcs1_mcs_mat1_1_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_13109, new_AGEMA_signal_13108, mcs1_mcs_mat1_1_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_9043, new_AGEMA_signal_9042, mcs1_mcs_mat1_1_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_13601, new_AGEMA_signal_13600, mcs1_mcs_mat1_1_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_12535, new_AGEMA_signal_12534, mcs1_mcs_mat1_1_mcs_out[7]}), .b ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .c ({new_AGEMA_signal_13109, new_AGEMA_signal_13108, mcs1_mcs_mat1_1_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_11665, new_AGEMA_signal_11664, mcs1_mcs_mat1_1_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .c ({new_AGEMA_signal_12535, new_AGEMA_signal_12534, mcs1_mcs_mat1_1_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_10705, new_AGEMA_signal_10704, mcs1_mcs_mat1_1_mcs_out[6]}), .b ({new_AGEMA_signal_8283, new_AGEMA_signal_8282, mcs1_mcs_mat1_1_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_11665, new_AGEMA_signal_11664, mcs1_mcs_mat1_1_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_8281, new_AGEMA_signal_8280, mcs1_mcs_mat1_1_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_9749, new_AGEMA_signal_9748, mcs1_mcs_mat1_1_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_10705, new_AGEMA_signal_10704, mcs1_mcs_mat1_1_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, shiftr_out[57]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({new_AGEMA_signal_9749, new_AGEMA_signal_9748, mcs1_mcs_mat1_1_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, shiftr_out[58]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1835], Fresh[1834], Fresh[1833]}), .c ({new_AGEMA_signal_8283, new_AGEMA_signal_8282, mcs1_mcs_mat1_1_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({new_AGEMA_signal_9043, new_AGEMA_signal_9042, mcs1_mcs_mat1_1_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_13111, new_AGEMA_signal_13110, mcs1_mcs_mat1_1_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_13603, new_AGEMA_signal_13602, mcs1_mcs_mat1_1_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_14075, new_AGEMA_signal_14074, mcs1_mcs_mat1_1_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .b ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, mcs1_mcs_mat1_1_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_13603, new_AGEMA_signal_13602, mcs1_mcs_mat1_1_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_14077, new_AGEMA_signal_14076, mcs1_mcs_mat1_1_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_11667, new_AGEMA_signal_11666, mcs1_mcs_mat1_1_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_14499, new_AGEMA_signal_14498, mcs1_mcs_mat1_1_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_14079, new_AGEMA_signal_14078, mcs1_mcs_mat1_1_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_13607, new_AGEMA_signal_13606, mcs1_mcs_mat1_1_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_14501, new_AGEMA_signal_14500, mcs1_mcs_mat1_1_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_13609, new_AGEMA_signal_13608, mcs1_mcs_mat1_1_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_10707, new_AGEMA_signal_10706, mcs1_mcs_mat1_1_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_14079, new_AGEMA_signal_14078, mcs1_mcs_mat1_1_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12995, new_AGEMA_signal_12994, shiftr_out[25]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1841], Fresh[1840], Fresh[1839]}), .c ({new_AGEMA_signal_13609, new_AGEMA_signal_13608, mcs1_mcs_mat1_1_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, shiftr_out[26]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({new_AGEMA_signal_11667, new_AGEMA_signal_11666, mcs1_mcs_mat1_1_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1847], Fresh[1846], Fresh[1845]}), .c ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, mcs1_mcs_mat1_1_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U96 ( .a ({new_AGEMA_signal_15551, new_AGEMA_signal_15550, mcs1_mcs_mat1_2_n128}), .b ({new_AGEMA_signal_12537, new_AGEMA_signal_12536, mcs1_mcs_mat1_2_n127}), .c ({temp_next_s2[85], temp_next_s1[85], temp_next_s0[85]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U95 ( .a ({new_AGEMA_signal_11739, new_AGEMA_signal_11738, mcs1_mcs_mat1_2_mcs_out[41]}), .b ({new_AGEMA_signal_9813, new_AGEMA_signal_9812, mcs1_mcs_mat1_2_mcs_out[45]}), .c ({new_AGEMA_signal_12537, new_AGEMA_signal_12536, mcs1_mcs_mat1_2_n127}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U94 ( .a ({new_AGEMA_signal_8779, new_AGEMA_signal_8778, mcs1_mcs_mat1_2_mcs_out[33]}), .b ({new_AGEMA_signal_15029, new_AGEMA_signal_15028, mcs1_mcs_mat1_2_mcs_out[37]}), .c ({new_AGEMA_signal_15551, new_AGEMA_signal_15550, mcs1_mcs_mat1_2_n128}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U93 ( .a ({new_AGEMA_signal_14503, new_AGEMA_signal_14502, mcs1_mcs_mat1_2_n126}), .b ({new_AGEMA_signal_13611, new_AGEMA_signal_13610, mcs1_mcs_mat1_2_n125}), .c ({temp_next_s2[84], temp_next_s1[84], temp_next_s0[84]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U92 ( .a ({new_AGEMA_signal_10783, new_AGEMA_signal_10782, mcs1_mcs_mat1_2_mcs_out[40]}), .b ({new_AGEMA_signal_13163, new_AGEMA_signal_13162, mcs1_mcs_mat1_2_mcs_out[44]}), .c ({new_AGEMA_signal_13611, new_AGEMA_signal_13610, mcs1_mcs_mat1_2_n125}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U91 ( .a ({new_AGEMA_signal_13171, new_AGEMA_signal_13170, mcs1_mcs_mat1_2_mcs_out[32]}), .b ({new_AGEMA_signal_14113, new_AGEMA_signal_14112, mcs1_mcs_mat1_2_mcs_out[36]}), .c ({new_AGEMA_signal_14503, new_AGEMA_signal_14502, mcs1_mcs_mat1_2_n126}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U90 ( .a ({new_AGEMA_signal_14505, new_AGEMA_signal_14504, mcs1_mcs_mat1_2_n124}), .b ({new_AGEMA_signal_13115, new_AGEMA_signal_13114, mcs1_mcs_mat1_2_n123}), .c ({temp_next_s2[55], temp_next_s1[55], temp_next_s0[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U89 ( .a ({new_AGEMA_signal_10797, new_AGEMA_signal_10796, mcs1_mcs_mat1_2_mcs_out[27]}), .b ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, mcs1_mcs_mat1_2_mcs_out[31]}), .c ({new_AGEMA_signal_13115, new_AGEMA_signal_13114, mcs1_mcs_mat1_2_n123}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U88 ( .a ({new_AGEMA_signal_10805, new_AGEMA_signal_10804, mcs1_mcs_mat1_2_mcs_out[19]}), .b ({new_AGEMA_signal_14115, new_AGEMA_signal_14114, mcs1_mcs_mat1_2_mcs_out[23]}), .c ({new_AGEMA_signal_14505, new_AGEMA_signal_14504, mcs1_mcs_mat1_2_n124}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U87 ( .a ({new_AGEMA_signal_14989, new_AGEMA_signal_14988, mcs1_mcs_mat1_2_n122}), .b ({new_AGEMA_signal_12539, new_AGEMA_signal_12538, mcs1_mcs_mat1_2_n121}), .c ({temp_next_s2[54], temp_next_s1[54], temp_next_s0[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U86 ( .a ({new_AGEMA_signal_11751, new_AGEMA_signal_11750, mcs1_mcs_mat1_2_mcs_out[26]}), .b ({new_AGEMA_signal_11747, new_AGEMA_signal_11746, mcs1_mcs_mat1_2_mcs_out[30]}), .c ({new_AGEMA_signal_12539, new_AGEMA_signal_12538, mcs1_mcs_mat1_2_n121}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U85 ( .a ({new_AGEMA_signal_11757, new_AGEMA_signal_11756, mcs1_mcs_mat1_2_mcs_out[18]}), .b ({new_AGEMA_signal_14547, new_AGEMA_signal_14546, mcs1_mcs_mat1_2_mcs_out[22]}), .c ({new_AGEMA_signal_14989, new_AGEMA_signal_14988, mcs1_mcs_mat1_2_n122}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U84 ( .a ({new_AGEMA_signal_15555, new_AGEMA_signal_15554, mcs1_mcs_mat1_2_n120}), .b ({new_AGEMA_signal_13117, new_AGEMA_signal_13116, mcs1_mcs_mat1_2_n119}), .c ({temp_next_s2[53], temp_next_s1[53], temp_next_s0[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U83 ( .a ({new_AGEMA_signal_12601, new_AGEMA_signal_12600, mcs1_mcs_mat1_2_mcs_out[25]}), .b ({new_AGEMA_signal_10793, new_AGEMA_signal_10792, mcs1_mcs_mat1_2_mcs_out[29]}), .c ({new_AGEMA_signal_13117, new_AGEMA_signal_13116, mcs1_mcs_mat1_2_n119}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U82 ( .a ({new_AGEMA_signal_12603, new_AGEMA_signal_12602, mcs1_mcs_mat1_2_mcs_out[17]}), .b ({new_AGEMA_signal_15031, new_AGEMA_signal_15030, mcs1_mcs_mat1_2_mcs_out[21]}), .c ({new_AGEMA_signal_15555, new_AGEMA_signal_15554, mcs1_mcs_mat1_2_n120}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U81 ( .a ({new_AGEMA_signal_14507, new_AGEMA_signal_14506, mcs1_mcs_mat1_2_n118}), .b ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, mcs1_mcs_mat1_2_n117}), .c ({temp_next_s2[52], temp_next_s1[52], temp_next_s0[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U80 ( .a ({new_AGEMA_signal_10801, new_AGEMA_signal_10800, mcs1_mcs_mat1_2_mcs_out[24]}), .b ({new_AGEMA_signal_12599, new_AGEMA_signal_12598, mcs1_mcs_mat1_2_mcs_out[28]}), .c ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, mcs1_mcs_mat1_2_n117}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U79 ( .a ({new_AGEMA_signal_10809, new_AGEMA_signal_10808, mcs1_mcs_mat1_2_mcs_out[16]}), .b ({new_AGEMA_signal_14119, new_AGEMA_signal_14118, mcs1_mcs_mat1_2_mcs_out[20]}), .c ({new_AGEMA_signal_14507, new_AGEMA_signal_14506, mcs1_mcs_mat1_2_n118}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U78 ( .a ({new_AGEMA_signal_13121, new_AGEMA_signal_13120, mcs1_mcs_mat1_2_n116}), .b ({new_AGEMA_signal_15557, new_AGEMA_signal_15556, mcs1_mcs_mat1_2_n115}), .c ({temp_next_s2[23], temp_next_s1[23], temp_next_s0[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U77 ( .a ({new_AGEMA_signal_10823, new_AGEMA_signal_10822, mcs1_mcs_mat1_2_mcs_out[3]}), .b ({new_AGEMA_signal_15033, new_AGEMA_signal_15032, mcs1_mcs_mat1_2_mcs_out[7]}), .c ({new_AGEMA_signal_15557, new_AGEMA_signal_15556, mcs1_mcs_mat1_2_n115}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U76 ( .a ({new_AGEMA_signal_9107, new_AGEMA_signal_9106, mcs1_mcs_mat1_2_mcs_out[11]}), .b ({new_AGEMA_signal_12605, new_AGEMA_signal_12604, mcs1_mcs_mat1_2_mcs_out[15]}), .c ({new_AGEMA_signal_13121, new_AGEMA_signal_13120, mcs1_mcs_mat1_2_n116}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U75 ( .a ({new_AGEMA_signal_15559, new_AGEMA_signal_15558, mcs1_mcs_mat1_2_n114}), .b ({new_AGEMA_signal_13123, new_AGEMA_signal_13122, mcs1_mcs_mat1_2_n113}), .c ({new_AGEMA_signal_16041, new_AGEMA_signal_16040, mcs_out[247]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U74 ( .a ({new_AGEMA_signal_12559, new_AGEMA_signal_12558, mcs1_mcs_mat1_2_mcs_out[123]}), .b ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_13123, new_AGEMA_signal_13122, mcs1_mcs_mat1_2_n113}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U73 ( .a ({new_AGEMA_signal_11685, new_AGEMA_signal_11684, mcs1_mcs_mat1_2_mcs_out[115]}), .b ({new_AGEMA_signal_15015, new_AGEMA_signal_15014, mcs1_mcs_mat1_2_mcs_out[119]}), .c ({new_AGEMA_signal_15559, new_AGEMA_signal_15558, mcs1_mcs_mat1_2_n114}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U72 ( .a ({new_AGEMA_signal_15561, new_AGEMA_signal_15560, mcs1_mcs_mat1_2_n112}), .b ({new_AGEMA_signal_10709, new_AGEMA_signal_10708, mcs1_mcs_mat1_2_n111}), .c ({new_AGEMA_signal_16043, new_AGEMA_signal_16042, mcs_out[246]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U71 ( .a ({new_AGEMA_signal_9751, new_AGEMA_signal_9750, mcs1_mcs_mat1_2_mcs_out[122]}), .b ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_10709, new_AGEMA_signal_10708, mcs1_mcs_mat1_2_n111}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U70 ( .a ({new_AGEMA_signal_10721, new_AGEMA_signal_10720, mcs1_mcs_mat1_2_mcs_out[114]}), .b ({new_AGEMA_signal_15017, new_AGEMA_signal_15016, mcs1_mcs_mat1_2_mcs_out[118]}), .c ({new_AGEMA_signal_15561, new_AGEMA_signal_15560, mcs1_mcs_mat1_2_n112}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U69 ( .a ({new_AGEMA_signal_12541, new_AGEMA_signal_12540, mcs1_mcs_mat1_2_n110}), .b ({new_AGEMA_signal_14509, new_AGEMA_signal_14508, mcs1_mcs_mat1_2_n109}), .c ({temp_next_s2[22], temp_next_s1[22], temp_next_s0[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U68 ( .a ({new_AGEMA_signal_10825, new_AGEMA_signal_10824, mcs1_mcs_mat1_2_mcs_out[2]}), .b ({new_AGEMA_signal_14121, new_AGEMA_signal_14120, mcs1_mcs_mat1_2_mcs_out[6]}), .c ({new_AGEMA_signal_14509, new_AGEMA_signal_14508, mcs1_mcs_mat1_2_n109}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U67 ( .a ({new_AGEMA_signal_11767, new_AGEMA_signal_11766, mcs1_mcs_mat1_2_mcs_out[10]}), .b ({new_AGEMA_signal_11761, new_AGEMA_signal_11760, mcs1_mcs_mat1_2_mcs_out[14]}), .c ({new_AGEMA_signal_12541, new_AGEMA_signal_12540, mcs1_mcs_mat1_2_n110}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U66 ( .a ({new_AGEMA_signal_14995, new_AGEMA_signal_14994, mcs1_mcs_mat1_2_n108}), .b ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, mcs1_mcs_mat1_2_n107}), .c ({new_AGEMA_signal_15563, new_AGEMA_signal_15562, mcs_out[245]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U65 ( .a ({new_AGEMA_signal_12561, new_AGEMA_signal_12560, mcs1_mcs_mat1_2_mcs_out[121]}), .b ({new_AGEMA_signal_9045, new_AGEMA_signal_9044, mcs1_mcs_mat1_2_mcs_out[125]}), .c ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, mcs1_mcs_mat1_2_n107}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U64 ( .a ({new_AGEMA_signal_9755, new_AGEMA_signal_9754, mcs1_mcs_mat1_2_mcs_out[113]}), .b ({new_AGEMA_signal_14527, new_AGEMA_signal_14526, mcs1_mcs_mat1_2_mcs_out[117]}), .c ({new_AGEMA_signal_14995, new_AGEMA_signal_14994, mcs1_mcs_mat1_2_n108}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U63 ( .a ({new_AGEMA_signal_14511, new_AGEMA_signal_14510, mcs1_mcs_mat1_2_n106}), .b ({new_AGEMA_signal_12543, new_AGEMA_signal_12542, mcs1_mcs_mat1_2_n105}), .c ({new_AGEMA_signal_14997, new_AGEMA_signal_14996, mcs_out[244]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U62 ( .a ({new_AGEMA_signal_11681, new_AGEMA_signal_11680, mcs1_mcs_mat1_2_mcs_out[120]}), .b ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_12543, new_AGEMA_signal_12542, mcs1_mcs_mat1_2_n105}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U61 ( .a ({new_AGEMA_signal_12563, new_AGEMA_signal_12562, mcs1_mcs_mat1_2_mcs_out[112]}), .b ({new_AGEMA_signal_14093, new_AGEMA_signal_14092, mcs1_mcs_mat1_2_mcs_out[116]}), .c ({new_AGEMA_signal_14511, new_AGEMA_signal_14510, mcs1_mcs_mat1_2_n106}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U60 ( .a ({new_AGEMA_signal_14999, new_AGEMA_signal_14998, mcs1_mcs_mat1_2_n104}), .b ({new_AGEMA_signal_13127, new_AGEMA_signal_13126, mcs1_mcs_mat1_2_n103}), .c ({new_AGEMA_signal_15565, new_AGEMA_signal_15564, mcs_out[215]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U59 ( .a ({new_AGEMA_signal_12565, new_AGEMA_signal_12564, mcs1_mcs_mat1_2_mcs_out[111]}), .b ({new_AGEMA_signal_12575, new_AGEMA_signal_12574, mcs1_mcs_mat1_2_mcs_out[99]}), .c ({new_AGEMA_signal_13127, new_AGEMA_signal_13126, mcs1_mcs_mat1_2_n103}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U58 ( .a ({new_AGEMA_signal_14529, new_AGEMA_signal_14528, mcs1_mcs_mat1_2_mcs_out[103]}), .b ({new_AGEMA_signal_11693, new_AGEMA_signal_11692, mcs1_mcs_mat1_2_mcs_out[107]}), .c ({new_AGEMA_signal_14999, new_AGEMA_signal_14998, mcs1_mcs_mat1_2_n104}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U57 ( .a ({new_AGEMA_signal_14081, new_AGEMA_signal_14080, mcs1_mcs_mat1_2_n102}), .b ({new_AGEMA_signal_13129, new_AGEMA_signal_13128, mcs1_mcs_mat1_2_n101}), .c ({new_AGEMA_signal_14513, new_AGEMA_signal_14512, mcs_out[214]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U56 ( .a ({new_AGEMA_signal_12567, new_AGEMA_signal_12566, mcs1_mcs_mat1_2_mcs_out[110]}), .b ({new_AGEMA_signal_10737, new_AGEMA_signal_10736, mcs1_mcs_mat1_2_mcs_out[98]}), .c ({new_AGEMA_signal_13129, new_AGEMA_signal_13128, mcs1_mcs_mat1_2_n101}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U55 ( .a ({new_AGEMA_signal_13625, new_AGEMA_signal_13624, mcs1_mcs_mat1_2_mcs_out[102]}), .b ({new_AGEMA_signal_11695, new_AGEMA_signal_11694, mcs1_mcs_mat1_2_mcs_out[106]}), .c ({new_AGEMA_signal_14081, new_AGEMA_signal_14080, mcs1_mcs_mat1_2_n102}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U54 ( .a ({new_AGEMA_signal_14515, new_AGEMA_signal_14514, mcs1_mcs_mat1_2_n100}), .b ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, mcs1_mcs_mat1_2_n99}), .c ({new_AGEMA_signal_15001, new_AGEMA_signal_15000, mcs_out[213]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U53 ( .a ({new_AGEMA_signal_12569, new_AGEMA_signal_12568, mcs1_mcs_mat1_2_mcs_out[109]}), .b ({new_AGEMA_signal_9061, new_AGEMA_signal_9060, mcs1_mcs_mat1_2_mcs_out[97]}), .c ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, mcs1_mcs_mat1_2_n99}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U52 ( .a ({new_AGEMA_signal_14097, new_AGEMA_signal_14096, mcs1_mcs_mat1_2_mcs_out[101]}), .b ({new_AGEMA_signal_11697, new_AGEMA_signal_11696, mcs1_mcs_mat1_2_mcs_out[105]}), .c ({new_AGEMA_signal_14515, new_AGEMA_signal_14514, mcs1_mcs_mat1_2_n100}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U51 ( .a ({new_AGEMA_signal_15003, new_AGEMA_signal_15002, mcs1_mcs_mat1_2_n98}), .b ({new_AGEMA_signal_14083, new_AGEMA_signal_14082, mcs1_mcs_mat1_2_n97}), .c ({new_AGEMA_signal_15567, new_AGEMA_signal_15566, mcs_out[212]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U50 ( .a ({new_AGEMA_signal_12571, new_AGEMA_signal_12570, mcs1_mcs_mat1_2_mcs_out[108]}), .b ({new_AGEMA_signal_13633, new_AGEMA_signal_13632, mcs1_mcs_mat1_2_mcs_out[96]}), .c ({new_AGEMA_signal_14083, new_AGEMA_signal_14082, mcs1_mcs_mat1_2_n97}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U49 ( .a ({new_AGEMA_signal_14531, new_AGEMA_signal_14530, mcs1_mcs_mat1_2_mcs_out[100]}), .b ({new_AGEMA_signal_12573, new_AGEMA_signal_12572, mcs1_mcs_mat1_2_mcs_out[104]}), .c ({new_AGEMA_signal_15003, new_AGEMA_signal_15002, mcs1_mcs_mat1_2_n98}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U48 ( .a ({new_AGEMA_signal_14085, new_AGEMA_signal_14084, mcs1_mcs_mat1_2_n96}), .b ({new_AGEMA_signal_12545, new_AGEMA_signal_12544, mcs1_mcs_mat1_2_n95}), .c ({new_AGEMA_signal_14517, new_AGEMA_signal_14516, mcs_out[183]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U47 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_11705, new_AGEMA_signal_11704, mcs1_mcs_mat1_2_mcs_out[95]}), .c ({new_AGEMA_signal_12545, new_AGEMA_signal_12544, mcs1_mcs_mat1_2_n95}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U46 ( .a ({new_AGEMA_signal_10741, new_AGEMA_signal_10740, mcs1_mcs_mat1_2_mcs_out[83]}), .b ({new_AGEMA_signal_13635, new_AGEMA_signal_13634, mcs1_mcs_mat1_2_mcs_out[87]}), .c ({new_AGEMA_signal_14085, new_AGEMA_signal_14084, mcs1_mcs_mat1_2_n96}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U45 ( .a ({new_AGEMA_signal_11669, new_AGEMA_signal_11668, mcs1_mcs_mat1_2_n94}), .b ({new_AGEMA_signal_10711, new_AGEMA_signal_10710, mcs1_mcs_mat1_2_n93}), .c ({new_AGEMA_signal_12547, new_AGEMA_signal_12546, mcs_out[182]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U43 ( .a ({new_AGEMA_signal_10743, new_AGEMA_signal_10742, mcs1_mcs_mat1_2_mcs_out[82]}), .b ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_11669, new_AGEMA_signal_11668, mcs1_mcs_mat1_2_n94}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U42 ( .a ({new_AGEMA_signal_13133, new_AGEMA_signal_13132, mcs1_mcs_mat1_2_n92}), .b ({new_AGEMA_signal_10713, new_AGEMA_signal_10712, mcs1_mcs_mat1_2_n91}), .c ({new_AGEMA_signal_13613, new_AGEMA_signal_13612, mcs_out[181]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U41 ( .a ({new_AGEMA_signal_9073, new_AGEMA_signal_9072, mcs1_mcs_mat1_2_mcs_out[89]}), .b ({new_AGEMA_signal_9773, new_AGEMA_signal_9772, mcs1_mcs_mat1_2_mcs_out[93]}), .c ({new_AGEMA_signal_10713, new_AGEMA_signal_10712, mcs1_mcs_mat1_2_n91}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U40 ( .a ({new_AGEMA_signal_10745, new_AGEMA_signal_10744, mcs1_mcs_mat1_2_mcs_out[81]}), .b ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_13133, new_AGEMA_signal_13132, mcs1_mcs_mat1_2_n92}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U39 ( .a ({new_AGEMA_signal_14519, new_AGEMA_signal_14518, mcs1_mcs_mat1_2_n90}), .b ({new_AGEMA_signal_13135, new_AGEMA_signal_13134, mcs1_mcs_mat1_2_n89}), .c ({new_AGEMA_signal_15005, new_AGEMA_signal_15004, mcs_out[180]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U38 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_12577, new_AGEMA_signal_12576, mcs1_mcs_mat1_2_mcs_out[92]}), .c ({new_AGEMA_signal_13135, new_AGEMA_signal_13134, mcs1_mcs_mat1_2_n89}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U37 ( .a ({new_AGEMA_signal_11709, new_AGEMA_signal_11708, mcs1_mcs_mat1_2_mcs_out[80]}), .b ({new_AGEMA_signal_14101, new_AGEMA_signal_14100, mcs1_mcs_mat1_2_mcs_out[84]}), .c ({new_AGEMA_signal_14519, new_AGEMA_signal_14518, mcs1_mcs_mat1_2_n90}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U36 ( .a ({new_AGEMA_signal_12549, new_AGEMA_signal_12548, mcs1_mcs_mat1_2_n88}), .b ({new_AGEMA_signal_13615, new_AGEMA_signal_13614, mcs1_mcs_mat1_2_n87}), .c ({temp_next_s2[21], temp_next_s1[21], temp_next_s0[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U35 ( .a ({new_AGEMA_signal_13177, new_AGEMA_signal_13176, mcs1_mcs_mat1_2_mcs_out[5]}), .b ({new_AGEMA_signal_10817, new_AGEMA_signal_10816, mcs1_mcs_mat1_2_mcs_out[9]}), .c ({new_AGEMA_signal_13615, new_AGEMA_signal_13614, mcs1_mcs_mat1_2_n87}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U34 ( .a ({new_AGEMA_signal_11763, new_AGEMA_signal_11762, mcs1_mcs_mat1_2_mcs_out[13]}), .b ({new_AGEMA_signal_11775, new_AGEMA_signal_11774, mcs1_mcs_mat1_2_mcs_out[1]}), .c ({new_AGEMA_signal_12549, new_AGEMA_signal_12548, mcs1_mcs_mat1_2_n88}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U33 ( .a ({new_AGEMA_signal_15007, new_AGEMA_signal_15006, mcs1_mcs_mat1_2_n86}), .b ({new_AGEMA_signal_12551, new_AGEMA_signal_12550, mcs1_mcs_mat1_2_n85}), .c ({new_AGEMA_signal_15569, new_AGEMA_signal_15568, mcs_out[151]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U32 ( .a ({new_AGEMA_signal_9789, new_AGEMA_signal_9788, mcs1_mcs_mat1_2_mcs_out[75]}), .b ({new_AGEMA_signal_11711, new_AGEMA_signal_11710, mcs1_mcs_mat1_2_mcs_out[79]}), .c ({new_AGEMA_signal_12551, new_AGEMA_signal_12550, mcs1_mcs_mat1_2_n85}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U31 ( .a ({new_AGEMA_signal_12585, new_AGEMA_signal_12584, mcs1_mcs_mat1_2_mcs_out[67]}), .b ({new_AGEMA_signal_14533, new_AGEMA_signal_14532, mcs1_mcs_mat1_2_mcs_out[71]}), .c ({new_AGEMA_signal_15007, new_AGEMA_signal_15006, mcs1_mcs_mat1_2_n86}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U30 ( .a ({new_AGEMA_signal_15571, new_AGEMA_signal_15570, mcs1_mcs_mat1_2_n84}), .b ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, mcs1_mcs_mat1_2_n83}), .c ({new_AGEMA_signal_16045, new_AGEMA_signal_16044, mcs_out[150]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U29 ( .a ({new_AGEMA_signal_12581, new_AGEMA_signal_12580, mcs1_mcs_mat1_2_mcs_out[74]}), .b ({new_AGEMA_signal_8305, new_AGEMA_signal_8304, mcs1_mcs_mat1_2_mcs_out[78]}), .c ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, mcs1_mcs_mat1_2_n83}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U28 ( .a ({new_AGEMA_signal_11721, new_AGEMA_signal_11720, mcs1_mcs_mat1_2_mcs_out[66]}), .b ({new_AGEMA_signal_15019, new_AGEMA_signal_15018, mcs1_mcs_mat1_2_mcs_out[70]}), .c ({new_AGEMA_signal_15571, new_AGEMA_signal_15570, mcs1_mcs_mat1_2_n84}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U27 ( .a ({new_AGEMA_signal_15573, new_AGEMA_signal_15572, mcs1_mcs_mat1_2_n82}), .b ({new_AGEMA_signal_11671, new_AGEMA_signal_11670, mcs1_mcs_mat1_2_n81}), .c ({new_AGEMA_signal_16047, new_AGEMA_signal_16046, mcs_out[149]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U26 ( .a ({new_AGEMA_signal_10751, new_AGEMA_signal_10750, mcs1_mcs_mat1_2_mcs_out[73]}), .b ({new_AGEMA_signal_9785, new_AGEMA_signal_9784, mcs1_mcs_mat1_2_mcs_out[77]}), .c ({new_AGEMA_signal_11671, new_AGEMA_signal_11670, mcs1_mcs_mat1_2_n81}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U25 ( .a ({new_AGEMA_signal_9795, new_AGEMA_signal_9794, mcs1_mcs_mat1_2_mcs_out[65]}), .b ({new_AGEMA_signal_15021, new_AGEMA_signal_15020, mcs1_mcs_mat1_2_mcs_out[69]}), .c ({new_AGEMA_signal_15573, new_AGEMA_signal_15572, mcs1_mcs_mat1_2_n82}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U24 ( .a ({new_AGEMA_signal_15009, new_AGEMA_signal_15008, mcs1_mcs_mat1_2_n80}), .b ({new_AGEMA_signal_13139, new_AGEMA_signal_13138, mcs1_mcs_mat1_2_n79}), .c ({new_AGEMA_signal_15575, new_AGEMA_signal_15574, mcs_out[148]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U23 ( .a ({new_AGEMA_signal_12583, new_AGEMA_signal_12582, mcs1_mcs_mat1_2_mcs_out[72]}), .b ({new_AGEMA_signal_12579, new_AGEMA_signal_12578, mcs1_mcs_mat1_2_mcs_out[76]}), .c ({new_AGEMA_signal_13139, new_AGEMA_signal_13138, mcs1_mcs_mat1_2_n79}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U22 ( .a ({new_AGEMA_signal_13159, new_AGEMA_signal_13158, mcs1_mcs_mat1_2_mcs_out[64]}), .b ({new_AGEMA_signal_14537, new_AGEMA_signal_14536, mcs1_mcs_mat1_2_mcs_out[68]}), .c ({new_AGEMA_signal_15009, new_AGEMA_signal_15008, mcs1_mcs_mat1_2_n80}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U21 ( .a ({new_AGEMA_signal_15011, new_AGEMA_signal_15010, mcs1_mcs_mat1_2_n78}), .b ({new_AGEMA_signal_12553, new_AGEMA_signal_12552, mcs1_mcs_mat1_2_n77}), .c ({temp_next_s2[119], temp_next_s1[119], temp_next_s0[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U20 ( .a ({new_AGEMA_signal_10765, new_AGEMA_signal_10764, mcs1_mcs_mat1_2_mcs_out[59]}), .b ({new_AGEMA_signal_11725, new_AGEMA_signal_11724, mcs1_mcs_mat1_2_mcs_out[63]}), .c ({new_AGEMA_signal_12553, new_AGEMA_signal_12552, mcs1_mcs_mat1_2_n77}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U19 ( .a ({new_AGEMA_signal_9811, new_AGEMA_signal_9810, mcs1_mcs_mat1_2_mcs_out[51]}), .b ({new_AGEMA_signal_14539, new_AGEMA_signal_14538, mcs1_mcs_mat1_2_mcs_out[55]}), .c ({new_AGEMA_signal_15011, new_AGEMA_signal_15010, mcs1_mcs_mat1_2_n78}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U18 ( .a ({new_AGEMA_signal_15579, new_AGEMA_signal_15578, mcs1_mcs_mat1_2_n76}), .b ({new_AGEMA_signal_11673, new_AGEMA_signal_11672, mcs1_mcs_mat1_2_n75}), .c ({temp_next_s2[118], temp_next_s1[118], temp_next_s0[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U17 ( .a ({new_AGEMA_signal_9803, new_AGEMA_signal_9802, mcs1_mcs_mat1_2_mcs_out[58]}), .b ({new_AGEMA_signal_10759, new_AGEMA_signal_10758, mcs1_mcs_mat1_2_mcs_out[62]}), .c ({new_AGEMA_signal_11673, new_AGEMA_signal_11672, mcs1_mcs_mat1_2_n75}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U16 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_15023, new_AGEMA_signal_15022, mcs1_mcs_mat1_2_mcs_out[54]}), .c ({new_AGEMA_signal_15579, new_AGEMA_signal_15578, mcs1_mcs_mat1_2_n76}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U15 ( .a ({new_AGEMA_signal_15581, new_AGEMA_signal_15580, mcs1_mcs_mat1_2_n74}), .b ({new_AGEMA_signal_11675, new_AGEMA_signal_11674, mcs1_mcs_mat1_2_n73}), .c ({temp_next_s2[117], temp_next_s1[117], temp_next_s0[117]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U14 ( .a ({new_AGEMA_signal_10767, new_AGEMA_signal_10766, mcs1_mcs_mat1_2_mcs_out[57]}), .b ({new_AGEMA_signal_10761, new_AGEMA_signal_10760, mcs1_mcs_mat1_2_mcs_out[61]}), .c ({new_AGEMA_signal_11675, new_AGEMA_signal_11674, mcs1_mcs_mat1_2_n73}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U13 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_15025, new_AGEMA_signal_15024, mcs1_mcs_mat1_2_mcs_out[53]}), .c ({new_AGEMA_signal_15581, new_AGEMA_signal_15580, mcs1_mcs_mat1_2_n74}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U12 ( .a ({new_AGEMA_signal_15013, new_AGEMA_signal_15012, mcs1_mcs_mat1_2_n72}), .b ({new_AGEMA_signal_13141, new_AGEMA_signal_13140, mcs1_mcs_mat1_2_n71}), .c ({temp_next_s2[116], temp_next_s1[116], temp_next_s0[116]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U11 ( .a ({new_AGEMA_signal_11729, new_AGEMA_signal_11728, mcs1_mcs_mat1_2_mcs_out[56]}), .b ({new_AGEMA_signal_12589, new_AGEMA_signal_12588, mcs1_mcs_mat1_2_mcs_out[60]}), .c ({new_AGEMA_signal_13141, new_AGEMA_signal_13140, mcs1_mcs_mat1_2_n71}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U10 ( .a ({new_AGEMA_signal_10773, new_AGEMA_signal_10772, mcs1_mcs_mat1_2_mcs_out[48]}), .b ({new_AGEMA_signal_14543, new_AGEMA_signal_14542, mcs1_mcs_mat1_2_mcs_out[52]}), .c ({new_AGEMA_signal_15013, new_AGEMA_signal_15012, mcs1_mcs_mat1_2_n72}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U9 ( .a ({new_AGEMA_signal_15585, new_AGEMA_signal_15584, mcs1_mcs_mat1_2_n70}), .b ({new_AGEMA_signal_12555, new_AGEMA_signal_12554, mcs1_mcs_mat1_2_n69}), .c ({temp_next_s2[87], temp_next_s1[87], temp_next_s0[87]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U8 ( .a ({new_AGEMA_signal_11735, new_AGEMA_signal_11734, mcs1_mcs_mat1_2_mcs_out[43]}), .b ({new_AGEMA_signal_11733, new_AGEMA_signal_11732, mcs1_mcs_mat1_2_mcs_out[47]}), .c ({new_AGEMA_signal_12555, new_AGEMA_signal_12554, mcs1_mcs_mat1_2_n69}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U7 ( .a ({new_AGEMA_signal_11743, new_AGEMA_signal_11742, mcs1_mcs_mat1_2_mcs_out[35]}), .b ({new_AGEMA_signal_15027, new_AGEMA_signal_15026, mcs1_mcs_mat1_2_mcs_out[39]}), .c ({new_AGEMA_signal_15585, new_AGEMA_signal_15584, mcs1_mcs_mat1_2_n70}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U6 ( .a ({new_AGEMA_signal_14089, new_AGEMA_signal_14088, mcs1_mcs_mat1_2_n68}), .b ({new_AGEMA_signal_12557, new_AGEMA_signal_12556, mcs1_mcs_mat1_2_n67}), .c ({temp_next_s2[86], temp_next_s1[86], temp_next_s0[86]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U5 ( .a ({new_AGEMA_signal_11737, new_AGEMA_signal_11736, mcs1_mcs_mat1_2_mcs_out[42]}), .b ({new_AGEMA_signal_9087, new_AGEMA_signal_9086, mcs1_mcs_mat1_2_mcs_out[46]}), .c ({new_AGEMA_signal_12557, new_AGEMA_signal_12556, mcs1_mcs_mat1_2_n67}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U4 ( .a ({new_AGEMA_signal_10787, new_AGEMA_signal_10786, mcs1_mcs_mat1_2_mcs_out[34]}), .b ({new_AGEMA_signal_13651, new_AGEMA_signal_13650, mcs1_mcs_mat1_2_mcs_out[38]}), .c ({new_AGEMA_signal_14089, new_AGEMA_signal_14088, mcs1_mcs_mat1_2_n68}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U3 ( .a ({new_AGEMA_signal_13617, new_AGEMA_signal_13616, mcs1_mcs_mat1_2_n66}), .b ({new_AGEMA_signal_16367, new_AGEMA_signal_16366, mcs1_mcs_mat1_2_n65}), .c ({temp_next_s2[20], temp_next_s1[20], temp_next_s0[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U2 ( .a ({new_AGEMA_signal_16055, new_AGEMA_signal_16054, mcs1_mcs_mat1_2_mcs_out[4]}), .b ({new_AGEMA_signal_12609, new_AGEMA_signal_12608, mcs1_mcs_mat1_2_mcs_out[8]}), .c ({new_AGEMA_signal_16367, new_AGEMA_signal_16366, mcs1_mcs_mat1_2_n65}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_U1 ( .a ({new_AGEMA_signal_11777, new_AGEMA_signal_11776, mcs1_mcs_mat1_2_mcs_out[0]}), .b ({new_AGEMA_signal_13175, new_AGEMA_signal_13174, mcs1_mcs_mat1_2_mcs_out[12]}), .c ({new_AGEMA_signal_13617, new_AGEMA_signal_13616, mcs1_mcs_mat1_2_n66}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_11677, new_AGEMA_signal_11676, mcs1_mcs_mat1_2_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_12559, new_AGEMA_signal_12558, mcs1_mcs_mat1_2_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_10715, new_AGEMA_signal_10714, mcs1_mcs_mat1_2_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_7753, new_AGEMA_signal_7752, mcs1_mcs_mat1_2_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_11677, new_AGEMA_signal_11676, mcs1_mcs_mat1_2_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_8285, new_AGEMA_signal_8284, mcs1_mcs_mat1_2_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_9047, new_AGEMA_signal_9046, mcs1_mcs_mat1_2_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_9751, new_AGEMA_signal_9750, mcs1_mcs_mat1_2_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_8287, new_AGEMA_signal_8286, mcs1_mcs_mat1_2_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .c ({new_AGEMA_signal_9047, new_AGEMA_signal_9046, mcs1_mcs_mat1_2_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_11679, new_AGEMA_signal_11678, mcs1_mcs_mat1_2_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .c ({new_AGEMA_signal_12561, new_AGEMA_signal_12560, mcs1_mcs_mat1_2_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_10715, new_AGEMA_signal_10714, mcs1_mcs_mat1_2_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_11679, new_AGEMA_signal_11678, mcs1_mcs_mat1_2_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_9753, new_AGEMA_signal_9752, mcs1_mcs_mat1_2_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9049, new_AGEMA_signal_9048, mcs1_mcs_mat1_2_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_10715, new_AGEMA_signal_10714, mcs1_mcs_mat1_2_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_10717, new_AGEMA_signal_10716, mcs1_mcs_mat1_2_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_11681, new_AGEMA_signal_11680, mcs1_mcs_mat1_2_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_9753, new_AGEMA_signal_9752, mcs1_mcs_mat1_2_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_8287, new_AGEMA_signal_8286, mcs1_mcs_mat1_2_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_10717, new_AGEMA_signal_10716, mcs1_mcs_mat1_2_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({new_AGEMA_signal_9753, new_AGEMA_signal_9752, mcs1_mcs_mat1_2_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1853], Fresh[1852], Fresh[1851]}), .c ({new_AGEMA_signal_8287, new_AGEMA_signal_8286, mcs1_mcs_mat1_2_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({new_AGEMA_signal_9049, new_AGEMA_signal_9048, mcs1_mcs_mat1_2_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_14523, new_AGEMA_signal_14522, mcs1_mcs_mat1_2_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .c ({new_AGEMA_signal_15015, new_AGEMA_signal_15014, mcs1_mcs_mat1_2_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_14091, new_AGEMA_signal_14090, mcs1_mcs_mat1_2_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_13147, new_AGEMA_signal_13146, mcs1_mcs_mat1_2_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_14523, new_AGEMA_signal_14522, mcs1_mcs_mat1_2_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_14525, new_AGEMA_signal_14524, mcs1_mcs_mat1_2_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_13621, new_AGEMA_signal_13620, mcs1_mcs_mat1_2_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_15017, new_AGEMA_signal_15016, mcs1_mcs_mat1_2_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_14091, new_AGEMA_signal_14090, mcs1_mcs_mat1_2_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .c ({new_AGEMA_signal_14525, new_AGEMA_signal_14524, mcs1_mcs_mat1_2_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_14091, new_AGEMA_signal_14090, mcs1_mcs_mat1_2_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_13619, new_AGEMA_signal_13618, mcs1_mcs_mat1_2_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_14527, new_AGEMA_signal_14526, mcs1_mcs_mat1_2_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_13623, new_AGEMA_signal_13622, mcs1_mcs_mat1_2_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_11683, new_AGEMA_signal_11682, mcs1_mcs_mat1_2_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_14091, new_AGEMA_signal_14090, mcs1_mcs_mat1_2_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_13145, new_AGEMA_signal_13144, mcs1_mcs_mat1_2_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_13621, new_AGEMA_signal_13620, mcs1_mcs_mat1_2_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_14093, new_AGEMA_signal_14092, mcs1_mcs_mat1_2_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_10719, new_AGEMA_signal_10718, mcs1_mcs_mat1_2_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_13147, new_AGEMA_signal_13146, mcs1_mcs_mat1_2_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_13621, new_AGEMA_signal_13620, mcs1_mcs_mat1_2_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_11683, new_AGEMA_signal_11682, mcs1_mcs_mat1_2_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_13145, new_AGEMA_signal_13144, mcs1_mcs_mat1_2_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1859], Fresh[1858], Fresh[1857]}), .c ({new_AGEMA_signal_13623, new_AGEMA_signal_13622, mcs1_mcs_mat1_2_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({new_AGEMA_signal_11683, new_AGEMA_signal_11682, mcs1_mcs_mat1_2_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1865], Fresh[1864], Fresh[1863]}), .c ({new_AGEMA_signal_13147, new_AGEMA_signal_13146, mcs1_mcs_mat1_2_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_10723, new_AGEMA_signal_10722, mcs1_mcs_mat1_2_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_8289, new_AGEMA_signal_8288, mcs1_mcs_mat1_2_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_11685, new_AGEMA_signal_11684, mcs1_mcs_mat1_2_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_9051, new_AGEMA_signal_9050, mcs1_mcs_mat1_2_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_9053, new_AGEMA_signal_9052, mcs1_mcs_mat1_2_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_9755, new_AGEMA_signal_9754, mcs1_mcs_mat1_2_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_10725, new_AGEMA_signal_10724, mcs1_mcs_mat1_2_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_11687, new_AGEMA_signal_11686, mcs1_mcs_mat1_2_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_12563, new_AGEMA_signal_12562, mcs1_mcs_mat1_2_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_10723, new_AGEMA_signal_10722, mcs1_mcs_mat1_2_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_11687, new_AGEMA_signal_11686, mcs1_mcs_mat1_2_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_7755, new_AGEMA_signal_7754, mcs1_mcs_mat1_2_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9759, new_AGEMA_signal_9758, mcs1_mcs_mat1_2_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_10723, new_AGEMA_signal_10722, mcs1_mcs_mat1_2_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_8291, new_AGEMA_signal_8290, mcs1_mcs_mat1_2_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_9757, new_AGEMA_signal_9756, mcs1_mcs_mat1_2_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_10725, new_AGEMA_signal_10724, mcs1_mcs_mat1_2_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({new_AGEMA_signal_9759, new_AGEMA_signal_9758, mcs1_mcs_mat1_2_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1871], Fresh[1870], Fresh[1869]}), .c ({new_AGEMA_signal_8291, new_AGEMA_signal_8290, mcs1_mcs_mat1_2_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({new_AGEMA_signal_9053, new_AGEMA_signal_9052, mcs1_mcs_mat1_2_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({new_AGEMA_signal_11689, new_AGEMA_signal_11688, mcs1_mcs_mat1_2_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12565, new_AGEMA_signal_12564, mcs1_mcs_mat1_2_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({new_AGEMA_signal_11691, new_AGEMA_signal_11690, mcs1_mcs_mat1_2_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12567, new_AGEMA_signal_12566, mcs1_mcs_mat1_2_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_9055, new_AGEMA_signal_9054, mcs1_mcs_mat1_2_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_11689, new_AGEMA_signal_11688, mcs1_mcs_mat1_2_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12569, new_AGEMA_signal_12568, mcs1_mcs_mat1_2_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_8293, new_AGEMA_signal_8292, mcs1_mcs_mat1_2_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_10727, new_AGEMA_signal_10726, mcs1_mcs_mat1_2_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_11689, new_AGEMA_signal_11688, mcs1_mcs_mat1_2_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_9761, new_AGEMA_signal_9760, mcs1_mcs_mat1_2_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_11691, new_AGEMA_signal_11690, mcs1_mcs_mat1_2_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12571, new_AGEMA_signal_12570, mcs1_mcs_mat1_2_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_10729, new_AGEMA_signal_10728, mcs1_mcs_mat1_2_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_11691, new_AGEMA_signal_11690, mcs1_mcs_mat1_2_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_9055, new_AGEMA_signal_9054, mcs1_mcs_mat1_2_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_9763, new_AGEMA_signal_9762, mcs1_mcs_mat1_2_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_10729, new_AGEMA_signal_10728, mcs1_mcs_mat1_2_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1877], Fresh[1876], Fresh[1875]}), .c ({new_AGEMA_signal_9763, new_AGEMA_signal_9762, mcs1_mcs_mat1_2_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({new_AGEMA_signal_8293, new_AGEMA_signal_8292, mcs1_mcs_mat1_2_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1883], Fresh[1882], Fresh[1881]}), .c ({new_AGEMA_signal_9055, new_AGEMA_signal_9054, mcs1_mcs_mat1_2_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_10733, new_AGEMA_signal_10732, mcs1_mcs_mat1_2_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_10731, new_AGEMA_signal_10730, mcs1_mcs_mat1_2_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_11693, new_AGEMA_signal_11692, mcs1_mcs_mat1_2_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_10731, new_AGEMA_signal_10730, mcs1_mcs_mat1_2_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_9057, new_AGEMA_signal_9056, mcs1_mcs_mat1_2_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_11695, new_AGEMA_signal_11694, mcs1_mcs_mat1_2_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_8295, new_AGEMA_signal_8294, mcs1_mcs_mat1_2_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .c ({new_AGEMA_signal_9057, new_AGEMA_signal_9056, mcs1_mcs_mat1_2_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_10731, new_AGEMA_signal_10730, mcs1_mcs_mat1_2_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_11697, new_AGEMA_signal_11696, mcs1_mcs_mat1_2_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_9767, new_AGEMA_signal_9766, mcs1_mcs_mat1_2_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_7759, new_AGEMA_signal_7758, mcs1_mcs_mat1_2_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_10731, new_AGEMA_signal_10730, mcs1_mcs_mat1_2_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_11699, new_AGEMA_signal_11698, mcs1_mcs_mat1_2_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_12573, new_AGEMA_signal_12572, mcs1_mcs_mat1_2_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_10733, new_AGEMA_signal_10732, mcs1_mcs_mat1_2_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_9767, new_AGEMA_signal_9766, mcs1_mcs_mat1_2_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_11699, new_AGEMA_signal_11698, mcs1_mcs_mat1_2_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_9765, new_AGEMA_signal_9764, mcs1_mcs_mat1_2_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .c ({new_AGEMA_signal_10733, new_AGEMA_signal_10732, mcs1_mcs_mat1_2_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_8295, new_AGEMA_signal_8294, mcs1_mcs_mat1_2_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_9059, new_AGEMA_signal_9058, mcs1_mcs_mat1_2_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_9765, new_AGEMA_signal_9764, mcs1_mcs_mat1_2_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({new_AGEMA_signal_9767, new_AGEMA_signal_9766, mcs1_mcs_mat1_2_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1889], Fresh[1888], Fresh[1887]}), .c ({new_AGEMA_signal_8295, new_AGEMA_signal_8294, mcs1_mcs_mat1_2_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({new_AGEMA_signal_9059, new_AGEMA_signal_9058, mcs1_mcs_mat1_2_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, mcs1_mcs_mat1_2_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_14095, new_AGEMA_signal_14094, mcs1_mcs_mat1_2_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_14529, new_AGEMA_signal_14528, mcs1_mcs_mat1_2_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_13631, new_AGEMA_signal_13630, mcs1_mcs_mat1_2_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_14095, new_AGEMA_signal_14094, mcs1_mcs_mat1_2_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_13627, new_AGEMA_signal_13626, mcs1_mcs_mat1_2_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_13151, new_AGEMA_signal_13150, mcs1_mcs_mat1_2_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_14097, new_AGEMA_signal_14096, mcs1_mcs_mat1_2_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_13629, new_AGEMA_signal_13628, mcs1_mcs_mat1_2_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_14099, new_AGEMA_signal_14098, mcs1_mcs_mat1_2_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_14531, new_AGEMA_signal_14530, mcs1_mcs_mat1_2_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_10735, new_AGEMA_signal_10734, mcs1_mcs_mat1_2_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_13631, new_AGEMA_signal_13630, mcs1_mcs_mat1_2_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_14099, new_AGEMA_signal_14098, mcs1_mcs_mat1_2_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_11701, new_AGEMA_signal_11700, mcs1_mcs_mat1_2_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .c ({new_AGEMA_signal_13629, new_AGEMA_signal_13628, mcs1_mcs_mat1_2_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1895], Fresh[1894], Fresh[1893]}), .c ({new_AGEMA_signal_13631, new_AGEMA_signal_13630, mcs1_mcs_mat1_2_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({new_AGEMA_signal_11701, new_AGEMA_signal_11700, mcs1_mcs_mat1_2_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1901], Fresh[1900], Fresh[1899]}), .c ({new_AGEMA_signal_13151, new_AGEMA_signal_13150, mcs1_mcs_mat1_2_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_13153, new_AGEMA_signal_13152, mcs1_mcs_mat1_2_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_9063, new_AGEMA_signal_9062, mcs1_mcs_mat1_2_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_13633, new_AGEMA_signal_13632, mcs1_mcs_mat1_2_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_12575, new_AGEMA_signal_12574, mcs1_mcs_mat1_2_mcs_out[99]}), .b ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .c ({new_AGEMA_signal_13153, new_AGEMA_signal_13152, mcs1_mcs_mat1_2_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_11703, new_AGEMA_signal_11702, mcs1_mcs_mat1_2_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .c ({new_AGEMA_signal_12575, new_AGEMA_signal_12574, mcs1_mcs_mat1_2_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_10737, new_AGEMA_signal_10736, mcs1_mcs_mat1_2_mcs_out[98]}), .b ({new_AGEMA_signal_8299, new_AGEMA_signal_8298, mcs1_mcs_mat1_2_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_11703, new_AGEMA_signal_11702, mcs1_mcs_mat1_2_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_8297, new_AGEMA_signal_8296, mcs1_mcs_mat1_2_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_9769, new_AGEMA_signal_9768, mcs1_mcs_mat1_2_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_10737, new_AGEMA_signal_10736, mcs1_mcs_mat1_2_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({new_AGEMA_signal_9769, new_AGEMA_signal_9768, mcs1_mcs_mat1_2_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1907], Fresh[1906], Fresh[1905]}), .c ({new_AGEMA_signal_8299, new_AGEMA_signal_8298, mcs1_mcs_mat1_2_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({new_AGEMA_signal_9063, new_AGEMA_signal_9062, mcs1_mcs_mat1_2_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_10739, new_AGEMA_signal_10738, mcs1_mcs_mat1_2_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_11705, new_AGEMA_signal_11704, mcs1_mcs_mat1_2_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_9067, new_AGEMA_signal_9066, mcs1_mcs_mat1_2_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_9069, new_AGEMA_signal_9068, mcs1_mcs_mat1_2_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_9773, new_AGEMA_signal_9772, mcs1_mcs_mat1_2_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_11707, new_AGEMA_signal_11706, mcs1_mcs_mat1_2_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_8301, new_AGEMA_signal_8300, mcs1_mcs_mat1_2_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_12577, new_AGEMA_signal_12576, mcs1_mcs_mat1_2_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_10739, new_AGEMA_signal_10738, mcs1_mcs_mat1_2_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_11707, new_AGEMA_signal_11706, mcs1_mcs_mat1_2_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_7763, new_AGEMA_signal_7762, mcs1_mcs_mat1_2_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_9775, new_AGEMA_signal_9774, mcs1_mcs_mat1_2_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_10739, new_AGEMA_signal_10738, mcs1_mcs_mat1_2_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1913], Fresh[1912], Fresh[1911]}), .c ({new_AGEMA_signal_9775, new_AGEMA_signal_9774, mcs1_mcs_mat1_2_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({new_AGEMA_signal_8301, new_AGEMA_signal_8300, mcs1_mcs_mat1_2_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1919], Fresh[1918], Fresh[1917]}), .c ({new_AGEMA_signal_9069, new_AGEMA_signal_9068, mcs1_mcs_mat1_2_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_9781, new_AGEMA_signal_9780, mcs1_mcs_mat1_2_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_9783, new_AGEMA_signal_9782, mcs1_mcs_mat1_2_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_10741, new_AGEMA_signal_10740, mcs1_mcs_mat1_2_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_9777, new_AGEMA_signal_9776, mcs1_mcs_mat1_2_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_7765, new_AGEMA_signal_7764, mcs1_mcs_mat1_2_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_10743, new_AGEMA_signal_10742, mcs1_mcs_mat1_2_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_9075, new_AGEMA_signal_9074, mcs1_mcs_mat1_2_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_9777, new_AGEMA_signal_9776, mcs1_mcs_mat1_2_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_9779, new_AGEMA_signal_9778, mcs1_mcs_mat1_2_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_10745, new_AGEMA_signal_10744, mcs1_mcs_mat1_2_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_8303, new_AGEMA_signal_8302, mcs1_mcs_mat1_2_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_9075, new_AGEMA_signal_9074, mcs1_mcs_mat1_2_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_9779, new_AGEMA_signal_9778, mcs1_mcs_mat1_2_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_10747, new_AGEMA_signal_10746, mcs1_mcs_mat1_2_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .c ({new_AGEMA_signal_11709, new_AGEMA_signal_11708, mcs1_mcs_mat1_2_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_9781, new_AGEMA_signal_9780, mcs1_mcs_mat1_2_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_8303, new_AGEMA_signal_8302, mcs1_mcs_mat1_2_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_10747, new_AGEMA_signal_10746, mcs1_mcs_mat1_2_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({new_AGEMA_signal_9783, new_AGEMA_signal_9782, mcs1_mcs_mat1_2_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1925], Fresh[1924], Fresh[1923]}), .c ({new_AGEMA_signal_8303, new_AGEMA_signal_8302, mcs1_mcs_mat1_2_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({new_AGEMA_signal_9075, new_AGEMA_signal_9074, mcs1_mcs_mat1_2_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_10749, new_AGEMA_signal_10748, mcs1_mcs_mat1_2_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_11711, new_AGEMA_signal_11710, mcs1_mcs_mat1_2_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_9077, new_AGEMA_signal_9076, mcs1_mcs_mat1_2_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_9785, new_AGEMA_signal_9784, mcs1_mcs_mat1_2_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_11713, new_AGEMA_signal_11712, mcs1_mcs_mat1_2_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_8307, new_AGEMA_signal_8306, mcs1_mcs_mat1_2_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_12579, new_AGEMA_signal_12578, mcs1_mcs_mat1_2_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_10749, new_AGEMA_signal_10748, mcs1_mcs_mat1_2_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .c ({new_AGEMA_signal_11713, new_AGEMA_signal_11712, mcs1_mcs_mat1_2_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_7767, new_AGEMA_signal_7766, mcs1_mcs_mat1_2_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_9787, new_AGEMA_signal_9786, mcs1_mcs_mat1_2_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_10749, new_AGEMA_signal_10748, mcs1_mcs_mat1_2_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1931], Fresh[1930], Fresh[1929]}), .c ({new_AGEMA_signal_9787, new_AGEMA_signal_9786, mcs1_mcs_mat1_2_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({new_AGEMA_signal_8307, new_AGEMA_signal_8306, mcs1_mcs_mat1_2_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1937], Fresh[1936], Fresh[1935]}), .c ({new_AGEMA_signal_9077, new_AGEMA_signal_9076, mcs1_mcs_mat1_2_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_11715, new_AGEMA_signal_11714, mcs1_mcs_mat1_2_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_12581, new_AGEMA_signal_12580, mcs1_mcs_mat1_2_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_10753, new_AGEMA_signal_10752, mcs1_mcs_mat1_2_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9791, new_AGEMA_signal_9790, mcs1_mcs_mat1_2_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_11715, new_AGEMA_signal_11714, mcs1_mcs_mat1_2_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_8777, new_AGEMA_signal_8776, mcs1_mcs_mat1_2_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_9789, new_AGEMA_signal_9788, mcs1_mcs_mat1_2_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_9791, new_AGEMA_signal_9790, mcs1_mcs_mat1_2_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_8777, new_AGEMA_signal_8776, mcs1_mcs_mat1_2_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_10751, new_AGEMA_signal_10750, mcs1_mcs_mat1_2_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_8309, new_AGEMA_signal_8308, mcs1_mcs_mat1_2_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_8311, new_AGEMA_signal_8310, mcs1_mcs_mat1_2_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_8777, new_AGEMA_signal_8776, mcs1_mcs_mat1_2_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_9079, new_AGEMA_signal_9078, mcs1_mcs_mat1_2_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .c ({new_AGEMA_signal_9791, new_AGEMA_signal_9790, mcs1_mcs_mat1_2_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_11717, new_AGEMA_signal_11716, mcs1_mcs_mat1_2_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_8309, new_AGEMA_signal_8308, mcs1_mcs_mat1_2_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_12583, new_AGEMA_signal_12582, mcs1_mcs_mat1_2_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_10753, new_AGEMA_signal_10752, mcs1_mcs_mat1_2_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9079, new_AGEMA_signal_9078, mcs1_mcs_mat1_2_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_11717, new_AGEMA_signal_11716, mcs1_mcs_mat1_2_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .b ({new_AGEMA_signal_9793, new_AGEMA_signal_9792, mcs1_mcs_mat1_2_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_10753, new_AGEMA_signal_10752, mcs1_mcs_mat1_2_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({new_AGEMA_signal_9793, new_AGEMA_signal_9792, mcs1_mcs_mat1_2_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1943], Fresh[1942], Fresh[1941]}), .c ({new_AGEMA_signal_8311, new_AGEMA_signal_8310, mcs1_mcs_mat1_2_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({new_AGEMA_signal_9079, new_AGEMA_signal_9078, mcs1_mcs_mat1_2_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_14103, new_AGEMA_signal_14102, mcs1_mcs_mat1_2_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, mcs1_mcs_mat1_2_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_14533, new_AGEMA_signal_14532, mcs1_mcs_mat1_2_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_13639, new_AGEMA_signal_13638, mcs1_mcs_mat1_2_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_14535, new_AGEMA_signal_14534, mcs1_mcs_mat1_2_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_15019, new_AGEMA_signal_15018, mcs1_mcs_mat1_2_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_14103, new_AGEMA_signal_14102, mcs1_mcs_mat1_2_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_14535, new_AGEMA_signal_14534, mcs1_mcs_mat1_2_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_15021, new_AGEMA_signal_15020, mcs1_mcs_mat1_2_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, mcs1_mcs_mat1_2_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_14105, new_AGEMA_signal_14104, mcs1_mcs_mat1_2_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_14535, new_AGEMA_signal_14534, mcs1_mcs_mat1_2_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({new_AGEMA_signal_11719, new_AGEMA_signal_11718, mcs1_mcs_mat1_2_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, mcs1_mcs_mat1_2_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_13637, new_AGEMA_signal_13636, mcs1_mcs_mat1_2_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .c ({new_AGEMA_signal_14103, new_AGEMA_signal_14102, mcs1_mcs_mat1_2_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_13157, new_AGEMA_signal_13156, mcs1_mcs_mat1_2_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_10755, new_AGEMA_signal_10754, mcs1_mcs_mat1_2_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_13637, new_AGEMA_signal_13636, mcs1_mcs_mat1_2_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_14105, new_AGEMA_signal_14104, mcs1_mcs_mat1_2_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_13639, new_AGEMA_signal_13638, mcs1_mcs_mat1_2_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_14537, new_AGEMA_signal_14536, mcs1_mcs_mat1_2_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_13157, new_AGEMA_signal_13156, mcs1_mcs_mat1_2_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_13639, new_AGEMA_signal_13638, mcs1_mcs_mat1_2_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({new_AGEMA_signal_13641, new_AGEMA_signal_13640, mcs1_mcs_mat1_2_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_14105, new_AGEMA_signal_14104, mcs1_mcs_mat1_2_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1949], Fresh[1948], Fresh[1947]}), .c ({new_AGEMA_signal_13641, new_AGEMA_signal_13640, mcs1_mcs_mat1_2_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({new_AGEMA_signal_11719, new_AGEMA_signal_11718, mcs1_mcs_mat1_2_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1955], Fresh[1954], Fresh[1953]}), .c ({new_AGEMA_signal_13157, new_AGEMA_signal_13156, mcs1_mcs_mat1_2_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_11723, new_AGEMA_signal_11722, mcs1_mcs_mat1_2_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_12585, new_AGEMA_signal_12584, mcs1_mcs_mat1_2_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({new_AGEMA_signal_10757, new_AGEMA_signal_10756, mcs1_mcs_mat1_2_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_11721, new_AGEMA_signal_11720, mcs1_mcs_mat1_2_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_12587, new_AGEMA_signal_12586, mcs1_mcs_mat1_2_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_9081, new_AGEMA_signal_9080, mcs1_mcs_mat1_2_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_13159, new_AGEMA_signal_13158, mcs1_mcs_mat1_2_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_11723, new_AGEMA_signal_11722, mcs1_mcs_mat1_2_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .c ({new_AGEMA_signal_12587, new_AGEMA_signal_12586, mcs1_mcs_mat1_2_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_8313, new_AGEMA_signal_8312, mcs1_mcs_mat1_2_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_10757, new_AGEMA_signal_10756, mcs1_mcs_mat1_2_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_11723, new_AGEMA_signal_11722, mcs1_mcs_mat1_2_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_7771, new_AGEMA_signal_7770, mcs1_mcs_mat1_2_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_9797, new_AGEMA_signal_9796, mcs1_mcs_mat1_2_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_10757, new_AGEMA_signal_10756, mcs1_mcs_mat1_2_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({new_AGEMA_signal_9797, new_AGEMA_signal_9796, mcs1_mcs_mat1_2_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1961], Fresh[1960], Fresh[1959]}), .c ({new_AGEMA_signal_8313, new_AGEMA_signal_8312, mcs1_mcs_mat1_2_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({new_AGEMA_signal_9081, new_AGEMA_signal_9080, mcs1_mcs_mat1_2_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_10763, new_AGEMA_signal_10762, mcs1_mcs_mat1_2_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_9083, new_AGEMA_signal_9082, mcs1_mcs_mat1_2_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_11725, new_AGEMA_signal_11724, mcs1_mcs_mat1_2_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_8315, new_AGEMA_signal_8314, mcs1_mcs_mat1_2_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_9799, new_AGEMA_signal_9798, mcs1_mcs_mat1_2_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_10759, new_AGEMA_signal_10758, mcs1_mcs_mat1_2_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({new_AGEMA_signal_9801, new_AGEMA_signal_9800, mcs1_mcs_mat1_2_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_10761, new_AGEMA_signal_10760, mcs1_mcs_mat1_2_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1967], Fresh[1966], Fresh[1965]}), .c ({new_AGEMA_signal_9801, new_AGEMA_signal_9800, mcs1_mcs_mat1_2_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({new_AGEMA_signal_8315, new_AGEMA_signal_8314, mcs1_mcs_mat1_2_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1973], Fresh[1972], Fresh[1971]}), .c ({new_AGEMA_signal_9083, new_AGEMA_signal_9082, mcs1_mcs_mat1_2_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_8319, new_AGEMA_signal_8318, mcs1_mcs_mat1_2_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_9085, new_AGEMA_signal_9084, mcs1_mcs_mat1_2_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_9803, new_AGEMA_signal_9802, mcs1_mcs_mat1_2_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_8321, new_AGEMA_signal_8320, mcs1_mcs_mat1_2_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_9805, new_AGEMA_signal_9804, mcs1_mcs_mat1_2_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_10767, new_AGEMA_signal_10766, mcs1_mcs_mat1_2_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_10769, new_AGEMA_signal_10768, mcs1_mcs_mat1_2_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_9807, new_AGEMA_signal_9806, mcs1_mcs_mat1_2_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_11729, new_AGEMA_signal_11728, mcs1_mcs_mat1_2_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_9809, new_AGEMA_signal_9808, mcs1_mcs_mat1_2_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_10769, new_AGEMA_signal_10768, mcs1_mcs_mat1_2_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({new_AGEMA_signal_9809, new_AGEMA_signal_9808, mcs1_mcs_mat1_2_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1979], Fresh[1978], Fresh[1977]}), .c ({new_AGEMA_signal_8321, new_AGEMA_signal_8320, mcs1_mcs_mat1_2_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({new_AGEMA_signal_9085, new_AGEMA_signal_9084, mcs1_mcs_mat1_2_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_13645, new_AGEMA_signal_13644, mcs1_mcs_mat1_2_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_14107, new_AGEMA_signal_14106, mcs1_mcs_mat1_2_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_14539, new_AGEMA_signal_14538, mcs1_mcs_mat1_2_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_14541, new_AGEMA_signal_14540, mcs1_mcs_mat1_2_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_13643, new_AGEMA_signal_13642, mcs1_mcs_mat1_2_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_15023, new_AGEMA_signal_15022, mcs1_mcs_mat1_2_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, mcs1_mcs_mat1_2_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_13643, new_AGEMA_signal_13642, mcs1_mcs_mat1_2_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({new_AGEMA_signal_14541, new_AGEMA_signal_14540, mcs1_mcs_mat1_2_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_15025, new_AGEMA_signal_15024, mcs1_mcs_mat1_2_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_10771, new_AGEMA_signal_10770, mcs1_mcs_mat1_2_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_14107, new_AGEMA_signal_14106, mcs1_mcs_mat1_2_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_14541, new_AGEMA_signal_14540, mcs1_mcs_mat1_2_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_11731, new_AGEMA_signal_11730, mcs1_mcs_mat1_2_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_13649, new_AGEMA_signal_13648, mcs1_mcs_mat1_2_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_14107, new_AGEMA_signal_14106, mcs1_mcs_mat1_2_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_13647, new_AGEMA_signal_13646, mcs1_mcs_mat1_2_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_14109, new_AGEMA_signal_14108, mcs1_mcs_mat1_2_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_14543, new_AGEMA_signal_14542, mcs1_mcs_mat1_2_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_13645, new_AGEMA_signal_13644, mcs1_mcs_mat1_2_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_11731, new_AGEMA_signal_11730, mcs1_mcs_mat1_2_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_14109, new_AGEMA_signal_14108, mcs1_mcs_mat1_2_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, mcs1_mcs_mat1_2_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_13645, new_AGEMA_signal_13644, mcs1_mcs_mat1_2_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1985], Fresh[1984], Fresh[1983]}), .c ({new_AGEMA_signal_13649, new_AGEMA_signal_13648, mcs1_mcs_mat1_2_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({new_AGEMA_signal_11731, new_AGEMA_signal_11730, mcs1_mcs_mat1_2_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1991], Fresh[1990], Fresh[1989]}), .c ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, mcs1_mcs_mat1_2_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_9089, new_AGEMA_signal_9088, mcs1_mcs_mat1_2_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_9813, new_AGEMA_signal_9812, mcs1_mcs_mat1_2_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_12591, new_AGEMA_signal_12590, mcs1_mcs_mat1_2_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_8323, new_AGEMA_signal_8322, mcs1_mcs_mat1_2_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_13163, new_AGEMA_signal_13162, mcs1_mcs_mat1_2_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_11733, new_AGEMA_signal_11732, mcs1_mcs_mat1_2_mcs_out[47]}), .b ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_12591, new_AGEMA_signal_12590, mcs1_mcs_mat1_2_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_10775, new_AGEMA_signal_10774, mcs1_mcs_mat1_2_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .c ({new_AGEMA_signal_11733, new_AGEMA_signal_11732, mcs1_mcs_mat1_2_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_7777, new_AGEMA_signal_7776, mcs1_mcs_mat1_2_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_9815, new_AGEMA_signal_9814, mcs1_mcs_mat1_2_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_10775, new_AGEMA_signal_10774, mcs1_mcs_mat1_2_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({new_AGEMA_signal_9815, new_AGEMA_signal_9814, mcs1_mcs_mat1_2_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1997], Fresh[1996], Fresh[1995]}), .c ({new_AGEMA_signal_8323, new_AGEMA_signal_8322, mcs1_mcs_mat1_2_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({new_AGEMA_signal_9089, new_AGEMA_signal_9088, mcs1_mcs_mat1_2_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_10777, new_AGEMA_signal_10776, mcs1_mcs_mat1_2_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_9091, new_AGEMA_signal_9090, mcs1_mcs_mat1_2_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_11735, new_AGEMA_signal_11734, mcs1_mcs_mat1_2_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_9817, new_AGEMA_signal_9816, mcs1_mcs_mat1_2_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8325, new_AGEMA_signal_8324, mcs1_mcs_mat1_2_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_10777, new_AGEMA_signal_10776, mcs1_mcs_mat1_2_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_10779, new_AGEMA_signal_10778, mcs1_mcs_mat1_2_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_9821, new_AGEMA_signal_9820, mcs1_mcs_mat1_2_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_11737, new_AGEMA_signal_11736, mcs1_mcs_mat1_2_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_10781, new_AGEMA_signal_10780, mcs1_mcs_mat1_2_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_7779, new_AGEMA_signal_7778, mcs1_mcs_mat1_2_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_11739, new_AGEMA_signal_11738, mcs1_mcs_mat1_2_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_9817, new_AGEMA_signal_9816, mcs1_mcs_mat1_2_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9093, new_AGEMA_signal_9092, mcs1_mcs_mat1_2_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_10781, new_AGEMA_signal_10780, mcs1_mcs_mat1_2_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_9819, new_AGEMA_signal_9818, mcs1_mcs_mat1_2_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_9093, new_AGEMA_signal_9092, mcs1_mcs_mat1_2_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_10783, new_AGEMA_signal_10782, mcs1_mcs_mat1_2_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2003], Fresh[2002], Fresh[2001]}), .c ({new_AGEMA_signal_9821, new_AGEMA_signal_9820, mcs1_mcs_mat1_2_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({new_AGEMA_signal_8325, new_AGEMA_signal_8324, mcs1_mcs_mat1_2_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2009], Fresh[2008], Fresh[2007]}), .c ({new_AGEMA_signal_9093, new_AGEMA_signal_9092, mcs1_mcs_mat1_2_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_14545, new_AGEMA_signal_14544, mcs1_mcs_mat1_2_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_10785, new_AGEMA_signal_10784, mcs1_mcs_mat1_2_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_15027, new_AGEMA_signal_15026, mcs1_mcs_mat1_2_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, mcs1_mcs_mat1_2_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_13165, new_AGEMA_signal_13164, mcs1_mcs_mat1_2_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_13651, new_AGEMA_signal_13650, mcs1_mcs_mat1_2_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({new_AGEMA_signal_14545, new_AGEMA_signal_14544, mcs1_mcs_mat1_2_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_15029, new_AGEMA_signal_15028, mcs1_mcs_mat1_2_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_13653, new_AGEMA_signal_13652, mcs1_mcs_mat1_2_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_14111, new_AGEMA_signal_14110, mcs1_mcs_mat1_2_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_14545, new_AGEMA_signal_14544, mcs1_mcs_mat1_2_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_13655, new_AGEMA_signal_13654, mcs1_mcs_mat1_2_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_13169, new_AGEMA_signal_13168, mcs1_mcs_mat1_2_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_14111, new_AGEMA_signal_14110, mcs1_mcs_mat1_2_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_13655, new_AGEMA_signal_13654, mcs1_mcs_mat1_2_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, mcs1_mcs_mat1_2_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_14113, new_AGEMA_signal_14112, mcs1_mcs_mat1_2_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_12593, new_AGEMA_signal_12592, mcs1_mcs_mat1_2_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, mcs1_mcs_mat1_2_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({new_AGEMA_signal_11741, new_AGEMA_signal_11740, mcs1_mcs_mat1_2_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_12593, new_AGEMA_signal_12592, mcs1_mcs_mat1_2_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({new_AGEMA_signal_13655, new_AGEMA_signal_13654, mcs1_mcs_mat1_2_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2015], Fresh[2014], Fresh[2013]}), .c ({new_AGEMA_signal_11741, new_AGEMA_signal_11740, mcs1_mcs_mat1_2_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({new_AGEMA_signal_13169, new_AGEMA_signal_13168, mcs1_mcs_mat1_2_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_9823, new_AGEMA_signal_9822, mcs1_mcs_mat1_2_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_9095, new_AGEMA_signal_9094, mcs1_mcs_mat1_2_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_10787, new_AGEMA_signal_10786, mcs1_mcs_mat1_2_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_8327, new_AGEMA_signal_8326, mcs1_mcs_mat1_2_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_8779, new_AGEMA_signal_8778, mcs1_mcs_mat1_2_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_12595, new_AGEMA_signal_12594, mcs1_mcs_mat1_2_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_9825, new_AGEMA_signal_9824, mcs1_mcs_mat1_2_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_13171, new_AGEMA_signal_13170, mcs1_mcs_mat1_2_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2021], Fresh[2020], Fresh[2019]}), .c ({new_AGEMA_signal_9825, new_AGEMA_signal_9824, mcs1_mcs_mat1_2_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({new_AGEMA_signal_8327, new_AGEMA_signal_8326, mcs1_mcs_mat1_2_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2027], Fresh[2026], Fresh[2025]}), .c ({new_AGEMA_signal_9095, new_AGEMA_signal_9094, mcs1_mcs_mat1_2_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_11745, new_AGEMA_signal_11744, mcs1_mcs_mat1_2_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_10791, new_AGEMA_signal_10790, mcs1_mcs_mat1_2_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, mcs1_mcs_mat1_2_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_8331, new_AGEMA_signal_8330, mcs1_mcs_mat1_2_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_10793, new_AGEMA_signal_10792, mcs1_mcs_mat1_2_mcs_out[29]}), .c ({new_AGEMA_signal_11745, new_AGEMA_signal_11744, mcs1_mcs_mat1_2_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_8329, new_AGEMA_signal_8328, mcs1_mcs_mat1_2_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_10791, new_AGEMA_signal_10790, mcs1_mcs_mat1_2_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_11747, new_AGEMA_signal_11746, mcs1_mcs_mat1_2_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, mcs1_mcs_mat1_2_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .c ({new_AGEMA_signal_10791, new_AGEMA_signal_10790, mcs1_mcs_mat1_2_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_11749, new_AGEMA_signal_11748, mcs1_mcs_mat1_2_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_9827, new_AGEMA_signal_9826, mcs1_mcs_mat1_2_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_12599, new_AGEMA_signal_12598, mcs1_mcs_mat1_2_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_10795, new_AGEMA_signal_10794, mcs1_mcs_mat1_2_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_9829, new_AGEMA_signal_9828, mcs1_mcs_mat1_2_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_11749, new_AGEMA_signal_11748, mcs1_mcs_mat1_2_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_9097, new_AGEMA_signal_9096, mcs1_mcs_mat1_2_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_9829, new_AGEMA_signal_9828, mcs1_mcs_mat1_2_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, mcs1_mcs_mat1_2_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8331, new_AGEMA_signal_8330, mcs1_mcs_mat1_2_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_10795, new_AGEMA_signal_10794, mcs1_mcs_mat1_2_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, mcs1_mcs_mat1_2_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2033], Fresh[2032], Fresh[2031]}), .c ({new_AGEMA_signal_8331, new_AGEMA_signal_8330, mcs1_mcs_mat1_2_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({new_AGEMA_signal_9097, new_AGEMA_signal_9096, mcs1_mcs_mat1_2_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_9833, new_AGEMA_signal_9832, mcs1_mcs_mat1_2_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_10797, new_AGEMA_signal_10796, mcs1_mcs_mat1_2_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_9099, new_AGEMA_signal_9098, mcs1_mcs_mat1_2_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8333, new_AGEMA_signal_8332, mcs1_mcs_mat1_2_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_9833, new_AGEMA_signal_9832, mcs1_mcs_mat1_2_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_10799, new_AGEMA_signal_10798, mcs1_mcs_mat1_2_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_11751, new_AGEMA_signal_11750, mcs1_mcs_mat1_2_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_9837, new_AGEMA_signal_9836, mcs1_mcs_mat1_2_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8333, new_AGEMA_signal_8332, mcs1_mcs_mat1_2_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_10799, new_AGEMA_signal_10798, mcs1_mcs_mat1_2_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_11753, new_AGEMA_signal_11752, mcs1_mcs_mat1_2_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .c ({new_AGEMA_signal_12601, new_AGEMA_signal_12600, mcs1_mcs_mat1_2_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_9837, new_AGEMA_signal_9836, mcs1_mcs_mat1_2_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_10801, new_AGEMA_signal_10800, mcs1_mcs_mat1_2_mcs_out[24]}), .c ({new_AGEMA_signal_11753, new_AGEMA_signal_11752, mcs1_mcs_mat1_2_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_9835, new_AGEMA_signal_9834, mcs1_mcs_mat1_2_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .c ({new_AGEMA_signal_10801, new_AGEMA_signal_10800, mcs1_mcs_mat1_2_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_9099, new_AGEMA_signal_9098, mcs1_mcs_mat1_2_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7785, new_AGEMA_signal_7784, mcs1_mcs_mat1_2_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_9835, new_AGEMA_signal_9834, mcs1_mcs_mat1_2_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2039], Fresh[2038], Fresh[2037]}), .c ({new_AGEMA_signal_9837, new_AGEMA_signal_9836, mcs1_mcs_mat1_2_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({new_AGEMA_signal_8333, new_AGEMA_signal_8332, mcs1_mcs_mat1_2_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2045], Fresh[2044], Fresh[2043]}), .c ({new_AGEMA_signal_9099, new_AGEMA_signal_9098, mcs1_mcs_mat1_2_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_13657, new_AGEMA_signal_13656, mcs1_mcs_mat1_2_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .c ({new_AGEMA_signal_14115, new_AGEMA_signal_14114, mcs1_mcs_mat1_2_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, mcs1_mcs_mat1_2_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_11755, new_AGEMA_signal_11754, mcs1_mcs_mat1_2_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_13657, new_AGEMA_signal_13656, mcs1_mcs_mat1_2_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_14117, new_AGEMA_signal_14116, mcs1_mcs_mat1_2_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .c ({new_AGEMA_signal_14547, new_AGEMA_signal_14546, mcs1_mcs_mat1_2_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_13661, new_AGEMA_signal_13660, mcs1_mcs_mat1_2_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_11755, new_AGEMA_signal_11754, mcs1_mcs_mat1_2_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_14117, new_AGEMA_signal_14116, mcs1_mcs_mat1_2_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_14549, new_AGEMA_signal_14548, mcs1_mcs_mat1_2_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_15031, new_AGEMA_signal_15030, mcs1_mcs_mat1_2_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_13661, new_AGEMA_signal_13660, mcs1_mcs_mat1_2_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_14119, new_AGEMA_signal_14118, mcs1_mcs_mat1_2_mcs_out[20]}), .c ({new_AGEMA_signal_14549, new_AGEMA_signal_14548, mcs1_mcs_mat1_2_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_13659, new_AGEMA_signal_13658, mcs1_mcs_mat1_2_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_14119, new_AGEMA_signal_14118, mcs1_mcs_mat1_2_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, mcs1_mcs_mat1_2_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_10803, new_AGEMA_signal_10802, mcs1_mcs_mat1_2_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_13659, new_AGEMA_signal_13658, mcs1_mcs_mat1_2_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({new_AGEMA_signal_13661, new_AGEMA_signal_13660, mcs1_mcs_mat1_2_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2051], Fresh[2050], Fresh[2049]}), .c ({new_AGEMA_signal_11755, new_AGEMA_signal_11754, mcs1_mcs_mat1_2_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, mcs1_mcs_mat1_2_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_9839, new_AGEMA_signal_9838, mcs1_mcs_mat1_2_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_9845, new_AGEMA_signal_9844, mcs1_mcs_mat1_2_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_10805, new_AGEMA_signal_10804, mcs1_mcs_mat1_2_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_10807, new_AGEMA_signal_10806, mcs1_mcs_mat1_2_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_7787, new_AGEMA_signal_7786, mcs1_mcs_mat1_2_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_11757, new_AGEMA_signal_11756, mcs1_mcs_mat1_2_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_11759, new_AGEMA_signal_11758, mcs1_mcs_mat1_2_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_8335, new_AGEMA_signal_8334, mcs1_mcs_mat1_2_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_12603, new_AGEMA_signal_12602, mcs1_mcs_mat1_2_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7528, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_10807, new_AGEMA_signal_10806, mcs1_mcs_mat1_2_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_11759, new_AGEMA_signal_11758, mcs1_mcs_mat1_2_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_9841, new_AGEMA_signal_9840, mcs1_mcs_mat1_2_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .c ({new_AGEMA_signal_10807, new_AGEMA_signal_10806, mcs1_mcs_mat1_2_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_9101, new_AGEMA_signal_9100, mcs1_mcs_mat1_2_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_9103, new_AGEMA_signal_9102, mcs1_mcs_mat1_2_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_9841, new_AGEMA_signal_9840, mcs1_mcs_mat1_2_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_9843, new_AGEMA_signal_9842, mcs1_mcs_mat1_2_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_8335, new_AGEMA_signal_8334, mcs1_mcs_mat1_2_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_10809, new_AGEMA_signal_10808, mcs1_mcs_mat1_2_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2057], Fresh[2056], Fresh[2055]}), .c ({new_AGEMA_signal_9845, new_AGEMA_signal_9844, mcs1_mcs_mat1_2_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({new_AGEMA_signal_8335, new_AGEMA_signal_8334, mcs1_mcs_mat1_2_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2063], Fresh[2062], Fresh[2061]}), .c ({new_AGEMA_signal_9103, new_AGEMA_signal_9102, mcs1_mcs_mat1_2_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_11765, new_AGEMA_signal_11764, mcs1_mcs_mat1_2_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_8781, new_AGEMA_signal_8780, mcs1_mcs_mat1_2_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_12605, new_AGEMA_signal_12604, mcs1_mcs_mat1_2_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_10815, new_AGEMA_signal_10814, mcs1_mcs_mat1_2_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_10811, new_AGEMA_signal_10810, mcs1_mcs_mat1_2_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_11761, new_AGEMA_signal_11760, mcs1_mcs_mat1_2_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_9849, new_AGEMA_signal_9848, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_8337, new_AGEMA_signal_8336, mcs1_mcs_mat1_2_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_10811, new_AGEMA_signal_10810, mcs1_mcs_mat1_2_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_8781, new_AGEMA_signal_8780, mcs1_mcs_mat1_2_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_10813, new_AGEMA_signal_10812, mcs1_mcs_mat1_2_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_11763, new_AGEMA_signal_11762, mcs1_mcs_mat1_2_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_9847, new_AGEMA_signal_9846, mcs1_mcs_mat1_2_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_9849, new_AGEMA_signal_9848, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_10813, new_AGEMA_signal_10812, mcs1_mcs_mat1_2_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_7789, new_AGEMA_signal_7788, mcs1_mcs_mat1_2_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_8337, new_AGEMA_signal_8336, mcs1_mcs_mat1_2_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8781, new_AGEMA_signal_8780, mcs1_mcs_mat1_2_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_12607, new_AGEMA_signal_12606, mcs1_mcs_mat1_2_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_13175, new_AGEMA_signal_13174, mcs1_mcs_mat1_2_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_11765, new_AGEMA_signal_11764, mcs1_mcs_mat1_2_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_9849, new_AGEMA_signal_9848, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_12607, new_AGEMA_signal_12606, mcs1_mcs_mat1_2_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_10815, new_AGEMA_signal_10814, mcs1_mcs_mat1_2_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_11765, new_AGEMA_signal_11764, mcs1_mcs_mat1_2_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_9847, new_AGEMA_signal_9846, mcs1_mcs_mat1_2_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_10815, new_AGEMA_signal_10814, mcs1_mcs_mat1_2_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_7493, new_AGEMA_signal_7492, shiftr_out[116]}), .b ({new_AGEMA_signal_9105, new_AGEMA_signal_9104, mcs1_mcs_mat1_2_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_9847, new_AGEMA_signal_9846, mcs1_mcs_mat1_2_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({new_AGEMA_signal_9849, new_AGEMA_signal_9848, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2069], Fresh[2068], Fresh[2067]}), .c ({new_AGEMA_signal_8337, new_AGEMA_signal_8336, mcs1_mcs_mat1_2_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({new_AGEMA_signal_9105, new_AGEMA_signal_9104, mcs1_mcs_mat1_2_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_8783, new_AGEMA_signal_8782, mcs1_mcs_mat1_2_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .c ({new_AGEMA_signal_9107, new_AGEMA_signal_9106, mcs1_mcs_mat1_2_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_10819, new_AGEMA_signal_10818, mcs1_mcs_mat1_2_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_11767, new_AGEMA_signal_11766, mcs1_mcs_mat1_2_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_9851, new_AGEMA_signal_9850, mcs1_mcs_mat1_2_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_10817, new_AGEMA_signal_10816, mcs1_mcs_mat1_2_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_9109, new_AGEMA_signal_9108, mcs1_mcs_mat1_2_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_8783, new_AGEMA_signal_8782, mcs1_mcs_mat1_2_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_9851, new_AGEMA_signal_9850, mcs1_mcs_mat1_2_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_7791, new_AGEMA_signal_7790, mcs1_mcs_mat1_2_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8339, new_AGEMA_signal_8338, mcs1_mcs_mat1_2_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_8783, new_AGEMA_signal_8782, mcs1_mcs_mat1_2_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_11769, new_AGEMA_signal_11768, mcs1_mcs_mat1_2_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, shiftr_out[84]}), .c ({new_AGEMA_signal_12609, new_AGEMA_signal_12608, mcs1_mcs_mat1_2_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_7791, new_AGEMA_signal_7790, mcs1_mcs_mat1_2_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_10819, new_AGEMA_signal_10818, mcs1_mcs_mat1_2_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_11769, new_AGEMA_signal_11768, mcs1_mcs_mat1_2_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_9853, new_AGEMA_signal_9852, mcs1_mcs_mat1_2_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_9109, new_AGEMA_signal_9108, mcs1_mcs_mat1_2_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_10819, new_AGEMA_signal_10818, mcs1_mcs_mat1_2_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2075], Fresh[2074], Fresh[2073]}), .c ({new_AGEMA_signal_9853, new_AGEMA_signal_9852, mcs1_mcs_mat1_2_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({new_AGEMA_signal_8339, new_AGEMA_signal_8338, mcs1_mcs_mat1_2_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, shiftr_out[87]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2081], Fresh[2080], Fresh[2079]}), .c ({new_AGEMA_signal_9109, new_AGEMA_signal_9108, mcs1_mcs_mat1_2_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_15587, new_AGEMA_signal_15586, mcs1_mcs_mat1_2_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, mcs1_mcs_mat1_2_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_16055, new_AGEMA_signal_16054, mcs1_mcs_mat1_2_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_15033, new_AGEMA_signal_15032, mcs1_mcs_mat1_2_mcs_out[7]}), .b ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .c ({new_AGEMA_signal_15587, new_AGEMA_signal_15586, mcs1_mcs_mat1_2_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_14551, new_AGEMA_signal_14550, mcs1_mcs_mat1_2_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .c ({new_AGEMA_signal_15033, new_AGEMA_signal_15032, mcs1_mcs_mat1_2_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_14121, new_AGEMA_signal_14120, mcs1_mcs_mat1_2_mcs_out[6]}), .b ({new_AGEMA_signal_11773, new_AGEMA_signal_11772, mcs1_mcs_mat1_2_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_14551, new_AGEMA_signal_14550, mcs1_mcs_mat1_2_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_11771, new_AGEMA_signal_11770, mcs1_mcs_mat1_2_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_13663, new_AGEMA_signal_13662, mcs1_mcs_mat1_2_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_14121, new_AGEMA_signal_14120, mcs1_mcs_mat1_2_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, shiftr_out[53]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({new_AGEMA_signal_13663, new_AGEMA_signal_13662, mcs1_mcs_mat1_2_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[54]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2087], Fresh[2086], Fresh[2085]}), .c ({new_AGEMA_signal_11773, new_AGEMA_signal_11772, mcs1_mcs_mat1_2_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12383, new_AGEMA_signal_12382, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, mcs1_mcs_mat1_2_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_9111, new_AGEMA_signal_9110, mcs1_mcs_mat1_2_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_9855, new_AGEMA_signal_9854, mcs1_mcs_mat1_2_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_10825, new_AGEMA_signal_10824, mcs1_mcs_mat1_2_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .b ({new_AGEMA_signal_9113, new_AGEMA_signal_9112, mcs1_mcs_mat1_2_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_9855, new_AGEMA_signal_9854, mcs1_mcs_mat1_2_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_10827, new_AGEMA_signal_10826, mcs1_mcs_mat1_2_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_8341, new_AGEMA_signal_8340, mcs1_mcs_mat1_2_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_11775, new_AGEMA_signal_11774, mcs1_mcs_mat1_2_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_10829, new_AGEMA_signal_10828, mcs1_mcs_mat1_2_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_9859, new_AGEMA_signal_9858, mcs1_mcs_mat1_2_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_11777, new_AGEMA_signal_11776, mcs1_mcs_mat1_2_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_9861, new_AGEMA_signal_9860, mcs1_mcs_mat1_2_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_7793, new_AGEMA_signal_7792, mcs1_mcs_mat1_2_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_10829, new_AGEMA_signal_10828, mcs1_mcs_mat1_2_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, shiftr_out[21]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2093], Fresh[2092], Fresh[2091]}), .c ({new_AGEMA_signal_9861, new_AGEMA_signal_9860, mcs1_mcs_mat1_2_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, shiftr_out[22]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({new_AGEMA_signal_8341, new_AGEMA_signal_8340, mcs1_mcs_mat1_2_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2099], Fresh[2098], Fresh[2097]}), .c ({new_AGEMA_signal_9113, new_AGEMA_signal_9112, mcs1_mcs_mat1_2_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U96 ( .a ({new_AGEMA_signal_13181, new_AGEMA_signal_13180, mcs1_mcs_mat1_3_n128}), .b ({new_AGEMA_signal_15035, new_AGEMA_signal_15034, mcs1_mcs_mat1_3_n127}), .c ({temp_next_s2[81], temp_next_s1[81], temp_next_s0[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U95 ( .a ({new_AGEMA_signal_14597, new_AGEMA_signal_14596, mcs1_mcs_mat1_3_mcs_out[41]}), .b ({new_AGEMA_signal_9933, new_AGEMA_signal_9932, mcs1_mcs_mat1_3_mcs_out[45]}), .c ({new_AGEMA_signal_15035, new_AGEMA_signal_15034, mcs1_mcs_mat1_3_n127}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U94 ( .a ({new_AGEMA_signal_8787, new_AGEMA_signal_8786, mcs1_mcs_mat1_3_mcs_out[33]}), .b ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, mcs1_mcs_mat1_3_mcs_out[37]}), .c ({new_AGEMA_signal_13181, new_AGEMA_signal_13180, mcs1_mcs_mat1_3_n128}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U93 ( .a ({new_AGEMA_signal_13665, new_AGEMA_signal_13664, mcs1_mcs_mat1_3_n126}), .b ({new_AGEMA_signal_14553, new_AGEMA_signal_14552, mcs1_mcs_mat1_3_n125}), .c ({temp_next_s2[80], temp_next_s1[80], temp_next_s0[80]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U92 ( .a ({new_AGEMA_signal_14163, new_AGEMA_signal_14162, mcs1_mcs_mat1_3_mcs_out[40]}), .b ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, mcs1_mcs_mat1_3_mcs_out[44]}), .c ({new_AGEMA_signal_14553, new_AGEMA_signal_14552, mcs1_mcs_mat1_3_n125}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U91 ( .a ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, mcs1_mcs_mat1_3_mcs_out[32]}), .b ({new_AGEMA_signal_10899, new_AGEMA_signal_10898, mcs1_mcs_mat1_3_mcs_out[36]}), .c ({new_AGEMA_signal_13665, new_AGEMA_signal_13664, mcs1_mcs_mat1_3_n126}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U90 ( .a ({new_AGEMA_signal_11779, new_AGEMA_signal_11778, mcs1_mcs_mat1_3_n124}), .b ({new_AGEMA_signal_14555, new_AGEMA_signal_14554, mcs1_mcs_mat1_3_n123}), .c ({temp_next_s2[51], temp_next_s1[51], temp_next_s0[51]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U89 ( .a ({new_AGEMA_signal_14165, new_AGEMA_signal_14164, mcs1_mcs_mat1_3_mcs_out[27]}), .b ({new_AGEMA_signal_12667, new_AGEMA_signal_12666, mcs1_mcs_mat1_3_mcs_out[31]}), .c ({new_AGEMA_signal_14555, new_AGEMA_signal_14554, mcs1_mcs_mat1_3_n123}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U88 ( .a ({new_AGEMA_signal_10919, new_AGEMA_signal_10918, mcs1_mcs_mat1_3_mcs_out[19]}), .b ({new_AGEMA_signal_10913, new_AGEMA_signal_10912, mcs1_mcs_mat1_3_mcs_out[23]}), .c ({new_AGEMA_signal_11779, new_AGEMA_signal_11778, mcs1_mcs_mat1_3_n124}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U87 ( .a ({new_AGEMA_signal_12611, new_AGEMA_signal_12610, mcs1_mcs_mat1_3_n122}), .b ({new_AGEMA_signal_15041, new_AGEMA_signal_15040, mcs1_mcs_mat1_3_n121}), .c ({temp_next_s2[50], temp_next_s1[50], temp_next_s0[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U86 ( .a ({new_AGEMA_signal_14599, new_AGEMA_signal_14598, mcs1_mcs_mat1_3_mcs_out[26]}), .b ({new_AGEMA_signal_11869, new_AGEMA_signal_11868, mcs1_mcs_mat1_3_mcs_out[30]}), .c ({new_AGEMA_signal_15041, new_AGEMA_signal_15040, mcs1_mcs_mat1_3_n121}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U85 ( .a ({new_AGEMA_signal_11879, new_AGEMA_signal_11878, mcs1_mcs_mat1_3_mcs_out[18]}), .b ({new_AGEMA_signal_11875, new_AGEMA_signal_11874, mcs1_mcs_mat1_3_mcs_out[22]}), .c ({new_AGEMA_signal_12611, new_AGEMA_signal_12610, mcs1_mcs_mat1_3_n122}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U84 ( .a ({new_AGEMA_signal_13183, new_AGEMA_signal_13182, mcs1_mcs_mat1_3_n120}), .b ({new_AGEMA_signal_15593, new_AGEMA_signal_15592, mcs1_mcs_mat1_3_n119}), .c ({temp_next_s2[49], temp_next_s1[49], temp_next_s0[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U83 ( .a ({new_AGEMA_signal_15079, new_AGEMA_signal_15078, mcs1_mcs_mat1_3_mcs_out[25]}), .b ({new_AGEMA_signal_10907, new_AGEMA_signal_10906, mcs1_mcs_mat1_3_mcs_out[29]}), .c ({new_AGEMA_signal_15593, new_AGEMA_signal_15592, mcs1_mcs_mat1_3_n119}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U82 ( .a ({new_AGEMA_signal_12673, new_AGEMA_signal_12672, mcs1_mcs_mat1_3_mcs_out[17]}), .b ({new_AGEMA_signal_12671, new_AGEMA_signal_12670, mcs1_mcs_mat1_3_mcs_out[21]}), .c ({new_AGEMA_signal_13183, new_AGEMA_signal_13182, mcs1_mcs_mat1_3_n120}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U81 ( .a ({new_AGEMA_signal_11781, new_AGEMA_signal_11780, mcs1_mcs_mat1_3_n118}), .b ({new_AGEMA_signal_14557, new_AGEMA_signal_14556, mcs1_mcs_mat1_3_n117}), .c ({temp_next_s2[48], temp_next_s1[48], temp_next_s0[48]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U80 ( .a ({new_AGEMA_signal_14169, new_AGEMA_signal_14168, mcs1_mcs_mat1_3_mcs_out[24]}), .b ({new_AGEMA_signal_12669, new_AGEMA_signal_12668, mcs1_mcs_mat1_3_mcs_out[28]}), .c ({new_AGEMA_signal_14557, new_AGEMA_signal_14556, mcs1_mcs_mat1_3_n117}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U79 ( .a ({new_AGEMA_signal_10923, new_AGEMA_signal_10922, mcs1_mcs_mat1_3_mcs_out[16]}), .b ({new_AGEMA_signal_10917, new_AGEMA_signal_10916, mcs1_mcs_mat1_3_mcs_out[20]}), .c ({new_AGEMA_signal_11781, new_AGEMA_signal_11780, mcs1_mcs_mat1_3_n118}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U78 ( .a ({new_AGEMA_signal_13667, new_AGEMA_signal_13666, mcs1_mcs_mat1_3_n116}), .b ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, mcs1_mcs_mat1_3_n115}), .c ({temp_next_s2[19], temp_next_s1[19], temp_next_s0[19]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U77 ( .a ({new_AGEMA_signal_10935, new_AGEMA_signal_10934, mcs1_mcs_mat1_3_mcs_out[3]}), .b ({new_AGEMA_signal_12681, new_AGEMA_signal_12680, mcs1_mcs_mat1_3_mcs_out[7]}), .c ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, mcs1_mcs_mat1_3_n115}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U76 ( .a ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, mcs1_mcs_mat1_3_mcs_out[11]}), .b ({new_AGEMA_signal_12675, new_AGEMA_signal_12674, mcs1_mcs_mat1_3_mcs_out[15]}), .c ({new_AGEMA_signal_13667, new_AGEMA_signal_13666, mcs1_mcs_mat1_3_n116}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U75 ( .a ({new_AGEMA_signal_13187, new_AGEMA_signal_13186, mcs1_mcs_mat1_3_n114}), .b ({new_AGEMA_signal_15595, new_AGEMA_signal_15594, mcs1_mcs_mat1_3_n113}), .c ({new_AGEMA_signal_16059, new_AGEMA_signal_16058, mcs_out[243]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U74 ( .a ({new_AGEMA_signal_15069, new_AGEMA_signal_15068, mcs1_mcs_mat1_3_mcs_out[123]}), .b ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_15595, new_AGEMA_signal_15594, mcs1_mcs_mat1_3_n113}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U73 ( .a ({new_AGEMA_signal_11803, new_AGEMA_signal_11802, mcs1_mcs_mat1_3_mcs_out[115]}), .b ({new_AGEMA_signal_12623, new_AGEMA_signal_12622, mcs1_mcs_mat1_3_mcs_out[119]}), .c ({new_AGEMA_signal_13187, new_AGEMA_signal_13186, mcs1_mcs_mat1_3_n114}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U72 ( .a ({new_AGEMA_signal_13189, new_AGEMA_signal_13188, mcs1_mcs_mat1_3_n112}), .b ({new_AGEMA_signal_14125, new_AGEMA_signal_14124, mcs1_mcs_mat1_3_n111}), .c ({new_AGEMA_signal_14559, new_AGEMA_signal_14558, mcs_out[242]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U71 ( .a ({new_AGEMA_signal_13681, new_AGEMA_signal_13680, mcs1_mcs_mat1_3_mcs_out[122]}), .b ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_14125, new_AGEMA_signal_14124, mcs1_mcs_mat1_3_n111}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U70 ( .a ({new_AGEMA_signal_10837, new_AGEMA_signal_10836, mcs1_mcs_mat1_3_mcs_out[114]}), .b ({new_AGEMA_signal_12625, new_AGEMA_signal_12624, mcs1_mcs_mat1_3_mcs_out[118]}), .c ({new_AGEMA_signal_13189, new_AGEMA_signal_13188, mcs1_mcs_mat1_3_n112}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U69 ( .a ({new_AGEMA_signal_15045, new_AGEMA_signal_15044, mcs1_mcs_mat1_3_n110}), .b ({new_AGEMA_signal_11783, new_AGEMA_signal_11782, mcs1_mcs_mat1_3_n109}), .c ({temp_next_s2[18], temp_next_s1[18], temp_next_s0[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U68 ( .a ({new_AGEMA_signal_10937, new_AGEMA_signal_10936, mcs1_mcs_mat1_3_mcs_out[2]}), .b ({new_AGEMA_signal_10933, new_AGEMA_signal_10932, mcs1_mcs_mat1_3_mcs_out[6]}), .c ({new_AGEMA_signal_11783, new_AGEMA_signal_11782, mcs1_mcs_mat1_3_n109}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U67 ( .a ({new_AGEMA_signal_14603, new_AGEMA_signal_14602, mcs1_mcs_mat1_3_mcs_out[10]}), .b ({new_AGEMA_signal_11883, new_AGEMA_signal_11882, mcs1_mcs_mat1_3_mcs_out[14]}), .c ({new_AGEMA_signal_15045, new_AGEMA_signal_15044, mcs1_mcs_mat1_3_n110}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U66 ( .a ({new_AGEMA_signal_12613, new_AGEMA_signal_12612, mcs1_mcs_mat1_3_n108}), .b ({new_AGEMA_signal_15599, new_AGEMA_signal_15598, mcs1_mcs_mat1_3_n107}), .c ({new_AGEMA_signal_16061, new_AGEMA_signal_16060, mcs_out[241]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U65 ( .a ({new_AGEMA_signal_15071, new_AGEMA_signal_15070, mcs1_mcs_mat1_3_mcs_out[121]}), .b ({new_AGEMA_signal_9115, new_AGEMA_signal_9114, mcs1_mcs_mat1_3_mcs_out[125]}), .c ({new_AGEMA_signal_15599, new_AGEMA_signal_15598, mcs1_mcs_mat1_3_n107}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U64 ( .a ({new_AGEMA_signal_9869, new_AGEMA_signal_9868, mcs1_mcs_mat1_3_mcs_out[113]}), .b ({new_AGEMA_signal_11801, new_AGEMA_signal_11800, mcs1_mcs_mat1_3_mcs_out[117]}), .c ({new_AGEMA_signal_12613, new_AGEMA_signal_12612, mcs1_mcs_mat1_3_n108}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U63 ( .a ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, mcs1_mcs_mat1_3_n106}), .b ({new_AGEMA_signal_15047, new_AGEMA_signal_15046, mcs1_mcs_mat1_3_n105}), .c ({new_AGEMA_signal_15601, new_AGEMA_signal_15600, mcs_out[240]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U62 ( .a ({new_AGEMA_signal_14577, new_AGEMA_signal_14576, mcs1_mcs_mat1_3_mcs_out[120]}), .b ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_15047, new_AGEMA_signal_15046, mcs1_mcs_mat1_3_n105}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U61 ( .a ({new_AGEMA_signal_12627, new_AGEMA_signal_12626, mcs1_mcs_mat1_3_mcs_out[112]}), .b ({new_AGEMA_signal_10835, new_AGEMA_signal_10834, mcs1_mcs_mat1_3_mcs_out[116]}), .c ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, mcs1_mcs_mat1_3_n106}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U60 ( .a ({new_AGEMA_signal_15049, new_AGEMA_signal_15048, mcs1_mcs_mat1_3_n104}), .b ({new_AGEMA_signal_13193, new_AGEMA_signal_13192, mcs1_mcs_mat1_3_n103}), .c ({new_AGEMA_signal_15603, new_AGEMA_signal_15602, mcs_out[211]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U59 ( .a ({new_AGEMA_signal_12629, new_AGEMA_signal_12628, mcs1_mcs_mat1_3_mcs_out[111]}), .b ({new_AGEMA_signal_12637, new_AGEMA_signal_12636, mcs1_mcs_mat1_3_mcs_out[99]}), .c ({new_AGEMA_signal_13193, new_AGEMA_signal_13192, mcs1_mcs_mat1_3_n103}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U58 ( .a ({new_AGEMA_signal_11813, new_AGEMA_signal_11812, mcs1_mcs_mat1_3_mcs_out[103]}), .b ({new_AGEMA_signal_14579, new_AGEMA_signal_14578, mcs1_mcs_mat1_3_mcs_out[107]}), .c ({new_AGEMA_signal_15049, new_AGEMA_signal_15048, mcs1_mcs_mat1_3_n104}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U57 ( .a ({new_AGEMA_signal_15051, new_AGEMA_signal_15050, mcs1_mcs_mat1_3_n102}), .b ({new_AGEMA_signal_13195, new_AGEMA_signal_13194, mcs1_mcs_mat1_3_n101}), .c ({new_AGEMA_signal_15605, new_AGEMA_signal_15604, mcs_out[210]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U56 ( .a ({new_AGEMA_signal_12631, new_AGEMA_signal_12630, mcs1_mcs_mat1_3_mcs_out[110]}), .b ({new_AGEMA_signal_10855, new_AGEMA_signal_10854, mcs1_mcs_mat1_3_mcs_out[98]}), .c ({new_AGEMA_signal_13195, new_AGEMA_signal_13194, mcs1_mcs_mat1_3_n101}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U55 ( .a ({new_AGEMA_signal_9879, new_AGEMA_signal_9878, mcs1_mcs_mat1_3_mcs_out[102]}), .b ({new_AGEMA_signal_14581, new_AGEMA_signal_14580, mcs1_mcs_mat1_3_mcs_out[106]}), .c ({new_AGEMA_signal_15051, new_AGEMA_signal_15050, mcs1_mcs_mat1_3_n102}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U54 ( .a ({new_AGEMA_signal_15053, new_AGEMA_signal_15052, mcs1_mcs_mat1_3_n100}), .b ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, mcs1_mcs_mat1_3_n99}), .c ({new_AGEMA_signal_15607, new_AGEMA_signal_15606, mcs_out[209]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U53 ( .a ({new_AGEMA_signal_12633, new_AGEMA_signal_12632, mcs1_mcs_mat1_3_mcs_out[109]}), .b ({new_AGEMA_signal_9133, new_AGEMA_signal_9132, mcs1_mcs_mat1_3_mcs_out[97]}), .c ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, mcs1_mcs_mat1_3_n99}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U52 ( .a ({new_AGEMA_signal_10851, new_AGEMA_signal_10850, mcs1_mcs_mat1_3_mcs_out[101]}), .b ({new_AGEMA_signal_14583, new_AGEMA_signal_14582, mcs1_mcs_mat1_3_mcs_out[105]}), .c ({new_AGEMA_signal_15053, new_AGEMA_signal_15052, mcs1_mcs_mat1_3_n100}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U51 ( .a ({new_AGEMA_signal_15609, new_AGEMA_signal_15608, mcs1_mcs_mat1_3_n98}), .b ({new_AGEMA_signal_14127, new_AGEMA_signal_14126, mcs1_mcs_mat1_3_n97}), .c ({new_AGEMA_signal_16063, new_AGEMA_signal_16062, mcs_out[208]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U50 ( .a ({new_AGEMA_signal_12635, new_AGEMA_signal_12634, mcs1_mcs_mat1_3_mcs_out[108]}), .b ({new_AGEMA_signal_13689, new_AGEMA_signal_13688, mcs1_mcs_mat1_3_mcs_out[96]}), .c ({new_AGEMA_signal_14127, new_AGEMA_signal_14126, mcs1_mcs_mat1_3_n97}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U49 ( .a ({new_AGEMA_signal_11815, new_AGEMA_signal_11814, mcs1_mcs_mat1_3_mcs_out[100]}), .b ({new_AGEMA_signal_15073, new_AGEMA_signal_15072, mcs1_mcs_mat1_3_mcs_out[104]}), .c ({new_AGEMA_signal_15609, new_AGEMA_signal_15608, mcs1_mcs_mat1_3_n98}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U48 ( .a ({new_AGEMA_signal_11785, new_AGEMA_signal_11784, mcs1_mcs_mat1_3_n96}), .b ({new_AGEMA_signal_13669, new_AGEMA_signal_13668, mcs1_mcs_mat1_3_n95}), .c ({new_AGEMA_signal_14129, new_AGEMA_signal_14128, mcs_out[179]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U47 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_11819, new_AGEMA_signal_11818, mcs1_mcs_mat1_3_mcs_out[95]}), .c ({new_AGEMA_signal_13669, new_AGEMA_signal_13668, mcs1_mcs_mat1_3_n95}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U46 ( .a ({new_AGEMA_signal_10861, new_AGEMA_signal_10860, mcs1_mcs_mat1_3_mcs_out[83]}), .b ({new_AGEMA_signal_9895, new_AGEMA_signal_9894, mcs1_mcs_mat1_3_mcs_out[87]}), .c ({new_AGEMA_signal_11785, new_AGEMA_signal_11784, mcs1_mcs_mat1_3_n96}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U45 ( .a ({new_AGEMA_signal_11787, new_AGEMA_signal_11786, mcs1_mcs_mat1_3_n94}), .b ({new_AGEMA_signal_13671, new_AGEMA_signal_13670, mcs1_mcs_mat1_3_n93}), .c ({new_AGEMA_signal_14131, new_AGEMA_signal_14130, mcs_out[178]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U43 ( .a ({new_AGEMA_signal_10863, new_AGEMA_signal_10862, mcs1_mcs_mat1_3_mcs_out[82]}), .b ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_11787, new_AGEMA_signal_11786, mcs1_mcs_mat1_3_n94}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U42 ( .a ({new_AGEMA_signal_11789, new_AGEMA_signal_11788, mcs1_mcs_mat1_3_n92}), .b ({new_AGEMA_signal_13673, new_AGEMA_signal_13672, mcs1_mcs_mat1_3_n91}), .c ({new_AGEMA_signal_14133, new_AGEMA_signal_14132, mcs_out[177]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U41 ( .a ({new_AGEMA_signal_13225, new_AGEMA_signal_13224, mcs1_mcs_mat1_3_mcs_out[89]}), .b ({new_AGEMA_signal_9891, new_AGEMA_signal_9890, mcs1_mcs_mat1_3_mcs_out[93]}), .c ({new_AGEMA_signal_13673, new_AGEMA_signal_13672, mcs1_mcs_mat1_3_n91}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U40 ( .a ({new_AGEMA_signal_10865, new_AGEMA_signal_10864, mcs1_mcs_mat1_3_mcs_out[81]}), .b ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_11789, new_AGEMA_signal_11788, mcs1_mcs_mat1_3_n92}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U39 ( .a ({new_AGEMA_signal_12615, new_AGEMA_signal_12614, mcs1_mcs_mat1_3_n90}), .b ({new_AGEMA_signal_13199, new_AGEMA_signal_13198, mcs1_mcs_mat1_3_n89}), .c ({new_AGEMA_signal_13675, new_AGEMA_signal_13674, mcs_out[176]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U38 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_12639, new_AGEMA_signal_12638, mcs1_mcs_mat1_3_mcs_out[92]}), .c ({new_AGEMA_signal_13199, new_AGEMA_signal_13198, mcs1_mcs_mat1_3_n89}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U37 ( .a ({new_AGEMA_signal_11823, new_AGEMA_signal_11822, mcs1_mcs_mat1_3_mcs_out[80]}), .b ({new_AGEMA_signal_10859, new_AGEMA_signal_10858, mcs1_mcs_mat1_3_mcs_out[84]}), .c ({new_AGEMA_signal_12615, new_AGEMA_signal_12614, mcs1_mcs_mat1_3_n90}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U36 ( .a ({new_AGEMA_signal_12617, new_AGEMA_signal_12616, mcs1_mcs_mat1_3_n88}), .b ({new_AGEMA_signal_14561, new_AGEMA_signal_14560, mcs1_mcs_mat1_3_n87}), .c ({temp_next_s2[17], temp_next_s1[17], temp_next_s0[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U35 ( .a ({new_AGEMA_signal_9179, new_AGEMA_signal_9178, mcs1_mcs_mat1_3_mcs_out[5]}), .b ({new_AGEMA_signal_14171, new_AGEMA_signal_14170, mcs1_mcs_mat1_3_mcs_out[9]}), .c ({new_AGEMA_signal_14561, new_AGEMA_signal_14560, mcs1_mcs_mat1_3_n87}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U34 ( .a ({new_AGEMA_signal_11885, new_AGEMA_signal_11884, mcs1_mcs_mat1_3_mcs_out[13]}), .b ({new_AGEMA_signal_11893, new_AGEMA_signal_11892, mcs1_mcs_mat1_3_mcs_out[1]}), .c ({new_AGEMA_signal_12617, new_AGEMA_signal_12616, mcs1_mcs_mat1_3_n88}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U33 ( .a ({new_AGEMA_signal_13201, new_AGEMA_signal_13200, mcs1_mcs_mat1_3_n86}), .b ({new_AGEMA_signal_14135, new_AGEMA_signal_14134, mcs1_mcs_mat1_3_n85}), .c ({new_AGEMA_signal_14563, new_AGEMA_signal_14562, mcs_out[147]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U32 ( .a ({new_AGEMA_signal_13691, new_AGEMA_signal_13690, mcs1_mcs_mat1_3_mcs_out[75]}), .b ({new_AGEMA_signal_11825, new_AGEMA_signal_11824, mcs1_mcs_mat1_3_mcs_out[79]}), .c ({new_AGEMA_signal_14135, new_AGEMA_signal_14134, mcs1_mcs_mat1_3_n85}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U31 ( .a ({new_AGEMA_signal_12649, new_AGEMA_signal_12648, mcs1_mcs_mat1_3_mcs_out[67]}), .b ({new_AGEMA_signal_11833, new_AGEMA_signal_11832, mcs1_mcs_mat1_3_mcs_out[71]}), .c ({new_AGEMA_signal_13201, new_AGEMA_signal_13200, mcs1_mcs_mat1_3_n86}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U30 ( .a ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, mcs1_mcs_mat1_3_n84}), .b ({new_AGEMA_signal_15611, new_AGEMA_signal_15610, mcs1_mcs_mat1_3_n83}), .c ({new_AGEMA_signal_16065, new_AGEMA_signal_16064, mcs_out[146]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U29 ( .a ({new_AGEMA_signal_15075, new_AGEMA_signal_15074, mcs1_mcs_mat1_3_mcs_out[74]}), .b ({new_AGEMA_signal_8361, new_AGEMA_signal_8360, mcs1_mcs_mat1_3_mcs_out[78]}), .c ({new_AGEMA_signal_15611, new_AGEMA_signal_15610, mcs1_mcs_mat1_3_n83}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U28 ( .a ({new_AGEMA_signal_11839, new_AGEMA_signal_11838, mcs1_mcs_mat1_3_mcs_out[66]}), .b ({new_AGEMA_signal_12645, new_AGEMA_signal_12644, mcs1_mcs_mat1_3_mcs_out[70]}), .c ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, mcs1_mcs_mat1_3_n84}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U27 ( .a ({new_AGEMA_signal_13205, new_AGEMA_signal_13204, mcs1_mcs_mat1_3_n82}), .b ({new_AGEMA_signal_14565, new_AGEMA_signal_14564, mcs1_mcs_mat1_3_n81}), .c ({new_AGEMA_signal_15057, new_AGEMA_signal_15056, mcs_out[145]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U26 ( .a ({new_AGEMA_signal_14147, new_AGEMA_signal_14146, mcs1_mcs_mat1_3_mcs_out[73]}), .b ({new_AGEMA_signal_9905, new_AGEMA_signal_9904, mcs1_mcs_mat1_3_mcs_out[77]}), .c ({new_AGEMA_signal_14565, new_AGEMA_signal_14564, mcs1_mcs_mat1_3_n81}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U25 ( .a ({new_AGEMA_signal_9915, new_AGEMA_signal_9914, mcs1_mcs_mat1_3_mcs_out[65]}), .b ({new_AGEMA_signal_12647, new_AGEMA_signal_12646, mcs1_mcs_mat1_3_mcs_out[69]}), .c ({new_AGEMA_signal_13205, new_AGEMA_signal_13204, mcs1_mcs_mat1_3_n82}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U24 ( .a ({new_AGEMA_signal_13677, new_AGEMA_signal_13676, mcs1_mcs_mat1_3_n80}), .b ({new_AGEMA_signal_15613, new_AGEMA_signal_15612, mcs1_mcs_mat1_3_n79}), .c ({new_AGEMA_signal_16067, new_AGEMA_signal_16066, mcs_out[144]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U23 ( .a ({new_AGEMA_signal_15077, new_AGEMA_signal_15076, mcs1_mcs_mat1_3_mcs_out[72]}), .b ({new_AGEMA_signal_12641, new_AGEMA_signal_12640, mcs1_mcs_mat1_3_mcs_out[76]}), .c ({new_AGEMA_signal_15613, new_AGEMA_signal_15612, mcs1_mcs_mat1_3_n79}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U22 ( .a ({new_AGEMA_signal_13229, new_AGEMA_signal_13228, mcs1_mcs_mat1_3_mcs_out[64]}), .b ({new_AGEMA_signal_11837, new_AGEMA_signal_11836, mcs1_mcs_mat1_3_mcs_out[68]}), .c ({new_AGEMA_signal_13677, new_AGEMA_signal_13676, mcs1_mcs_mat1_3_n80}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U21 ( .a ({new_AGEMA_signal_12619, new_AGEMA_signal_12618, mcs1_mcs_mat1_3_n78}), .b ({new_AGEMA_signal_14567, new_AGEMA_signal_14566, mcs1_mcs_mat1_3_n77}), .c ({temp_next_s2[115], temp_next_s1[115], temp_next_s0[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U20 ( .a ({new_AGEMA_signal_14151, new_AGEMA_signal_14150, mcs1_mcs_mat1_3_mcs_out[59]}), .b ({new_AGEMA_signal_11843, new_AGEMA_signal_11842, mcs1_mcs_mat1_3_mcs_out[63]}), .c ({new_AGEMA_signal_14567, new_AGEMA_signal_14566, mcs1_mcs_mat1_3_n77}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U19 ( .a ({new_AGEMA_signal_9931, new_AGEMA_signal_9930, mcs1_mcs_mat1_3_mcs_out[51]}), .b ({new_AGEMA_signal_11853, new_AGEMA_signal_11852, mcs1_mcs_mat1_3_mcs_out[55]}), .c ({new_AGEMA_signal_12619, new_AGEMA_signal_12618, mcs1_mcs_mat1_3_n78}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U18 ( .a ({new_AGEMA_signal_13207, new_AGEMA_signal_13206, mcs1_mcs_mat1_3_n76}), .b ({new_AGEMA_signal_14137, new_AGEMA_signal_14136, mcs1_mcs_mat1_3_n75}), .c ({temp_next_s2[114], temp_next_s1[114], temp_next_s0[114]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U17 ( .a ({new_AGEMA_signal_13697, new_AGEMA_signal_13696, mcs1_mcs_mat1_3_mcs_out[58]}), .b ({new_AGEMA_signal_10879, new_AGEMA_signal_10878, mcs1_mcs_mat1_3_mcs_out[62]}), .c ({new_AGEMA_signal_14137, new_AGEMA_signal_14136, mcs1_mcs_mat1_3_n75}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U16 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_12655, new_AGEMA_signal_12654, mcs1_mcs_mat1_3_mcs_out[54]}), .c ({new_AGEMA_signal_13207, new_AGEMA_signal_13206, mcs1_mcs_mat1_3_n76}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U15 ( .a ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, mcs1_mcs_mat1_3_n74}), .b ({new_AGEMA_signal_14571, new_AGEMA_signal_14570, mcs1_mcs_mat1_3_n73}), .c ({temp_next_s2[113], temp_next_s1[113], temp_next_s0[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U14 ( .a ({new_AGEMA_signal_14153, new_AGEMA_signal_14152, mcs1_mcs_mat1_3_mcs_out[57]}), .b ({new_AGEMA_signal_10881, new_AGEMA_signal_10880, mcs1_mcs_mat1_3_mcs_out[61]}), .c ({new_AGEMA_signal_14571, new_AGEMA_signal_14570, mcs1_mcs_mat1_3_n73}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U13 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_12657, new_AGEMA_signal_12656, mcs1_mcs_mat1_3_mcs_out[53]}), .c ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, mcs1_mcs_mat1_3_n74}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U12 ( .a ({new_AGEMA_signal_12621, new_AGEMA_signal_12620, mcs1_mcs_mat1_3_n72}), .b ({new_AGEMA_signal_15063, new_AGEMA_signal_15062, mcs1_mcs_mat1_3_n71}), .c ({temp_next_s2[112], temp_next_s1[112], temp_next_s0[112]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U11 ( .a ({new_AGEMA_signal_14591, new_AGEMA_signal_14590, mcs1_mcs_mat1_3_mcs_out[56]}), .b ({new_AGEMA_signal_12653, new_AGEMA_signal_12652, mcs1_mcs_mat1_3_mcs_out[60]}), .c ({new_AGEMA_signal_15063, new_AGEMA_signal_15062, mcs1_mcs_mat1_3_n71}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U10 ( .a ({new_AGEMA_signal_10891, new_AGEMA_signal_10890, mcs1_mcs_mat1_3_mcs_out[48]}), .b ({new_AGEMA_signal_11857, new_AGEMA_signal_11856, mcs1_mcs_mat1_3_mcs_out[52]}), .c ({new_AGEMA_signal_12621, new_AGEMA_signal_12620, mcs1_mcs_mat1_3_n72}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U9 ( .a ({new_AGEMA_signal_13211, new_AGEMA_signal_13210, mcs1_mcs_mat1_3_n70}), .b ({new_AGEMA_signal_15065, new_AGEMA_signal_15064, mcs1_mcs_mat1_3_n69}), .c ({temp_next_s2[83], temp_next_s1[83], temp_next_s0[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U8 ( .a ({new_AGEMA_signal_14593, new_AGEMA_signal_14592, mcs1_mcs_mat1_3_mcs_out[43]}), .b ({new_AGEMA_signal_11859, new_AGEMA_signal_11858, mcs1_mcs_mat1_3_mcs_out[47]}), .c ({new_AGEMA_signal_15065, new_AGEMA_signal_15064, mcs1_mcs_mat1_3_n69}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U7 ( .a ({new_AGEMA_signal_11865, new_AGEMA_signal_11864, mcs1_mcs_mat1_3_mcs_out[35]}), .b ({new_AGEMA_signal_12661, new_AGEMA_signal_12660, mcs1_mcs_mat1_3_mcs_out[39]}), .c ({new_AGEMA_signal_13211, new_AGEMA_signal_13210, mcs1_mcs_mat1_3_n70}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U6 ( .a ({new_AGEMA_signal_11791, new_AGEMA_signal_11790, mcs1_mcs_mat1_3_n68}), .b ({new_AGEMA_signal_15067, new_AGEMA_signal_15066, mcs1_mcs_mat1_3_n67}), .c ({temp_next_s2[82], temp_next_s1[82], temp_next_s0[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U5 ( .a ({new_AGEMA_signal_14595, new_AGEMA_signal_14594, mcs1_mcs_mat1_3_mcs_out[42]}), .b ({new_AGEMA_signal_9157, new_AGEMA_signal_9156, mcs1_mcs_mat1_3_mcs_out[46]}), .c ({new_AGEMA_signal_15067, new_AGEMA_signal_15066, mcs1_mcs_mat1_3_n67}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U4 ( .a ({new_AGEMA_signal_10901, new_AGEMA_signal_10900, mcs1_mcs_mat1_3_mcs_out[34]}), .b ({new_AGEMA_signal_9937, new_AGEMA_signal_9936, mcs1_mcs_mat1_3_mcs_out[38]}), .c ({new_AGEMA_signal_11791, new_AGEMA_signal_11790, mcs1_mcs_mat1_3_n68}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U3 ( .a ({new_AGEMA_signal_13679, new_AGEMA_signal_13678, mcs1_mcs_mat1_3_n66}), .b ({new_AGEMA_signal_15621, new_AGEMA_signal_15620, mcs1_mcs_mat1_3_n65}), .c ({temp_next_s2[16], temp_next_s1[16], temp_next_s0[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U2 ( .a ({new_AGEMA_signal_13721, new_AGEMA_signal_13720, mcs1_mcs_mat1_3_mcs_out[4]}), .b ({new_AGEMA_signal_15081, new_AGEMA_signal_15080, mcs1_mcs_mat1_3_mcs_out[8]}), .c ({new_AGEMA_signal_15621, new_AGEMA_signal_15620, mcs1_mcs_mat1_3_n65}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_U1 ( .a ({new_AGEMA_signal_11895, new_AGEMA_signal_11894, mcs1_mcs_mat1_3_mcs_out[0]}), .b ({new_AGEMA_signal_13243, new_AGEMA_signal_13242, mcs1_mcs_mat1_3_mcs_out[12]}), .c ({new_AGEMA_signal_13679, new_AGEMA_signal_13678, mcs1_mcs_mat1_3_n66}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_14573, new_AGEMA_signal_14572, mcs1_mcs_mat1_3_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_15069, new_AGEMA_signal_15068, mcs1_mcs_mat1_3_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_14139, new_AGEMA_signal_14138, mcs1_mcs_mat1_3_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_10831, new_AGEMA_signal_10830, mcs1_mcs_mat1_3_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_14573, new_AGEMA_signal_14572, mcs1_mcs_mat1_3_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, mcs1_mcs_mat1_3_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_13213, new_AGEMA_signal_13212, mcs1_mcs_mat1_3_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_13681, new_AGEMA_signal_13680, mcs1_mcs_mat1_3_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_11795, new_AGEMA_signal_11794, mcs1_mcs_mat1_3_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .c ({new_AGEMA_signal_13213, new_AGEMA_signal_13212, mcs1_mcs_mat1_3_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_14575, new_AGEMA_signal_14574, mcs1_mcs_mat1_3_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .c ({new_AGEMA_signal_15071, new_AGEMA_signal_15070, mcs1_mcs_mat1_3_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_14139, new_AGEMA_signal_14138, mcs1_mcs_mat1_3_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_14575, new_AGEMA_signal_14574, mcs1_mcs_mat1_3_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_13683, new_AGEMA_signal_13682, mcs1_mcs_mat1_3_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, mcs1_mcs_mat1_3_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_14139, new_AGEMA_signal_14138, mcs1_mcs_mat1_3_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_14141, new_AGEMA_signal_14140, mcs1_mcs_mat1_3_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_14577, new_AGEMA_signal_14576, mcs1_mcs_mat1_3_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_13683, new_AGEMA_signal_13682, mcs1_mcs_mat1_3_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_11795, new_AGEMA_signal_11794, mcs1_mcs_mat1_3_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_14141, new_AGEMA_signal_14140, mcs1_mcs_mat1_3_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({new_AGEMA_signal_13683, new_AGEMA_signal_13682, mcs1_mcs_mat1_3_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2105], Fresh[2104], Fresh[2103]}), .c ({new_AGEMA_signal_11795, new_AGEMA_signal_11794, mcs1_mcs_mat1_3_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, mcs1_mcs_mat1_3_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_11797, new_AGEMA_signal_11796, mcs1_mcs_mat1_3_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .c ({new_AGEMA_signal_12623, new_AGEMA_signal_12622, mcs1_mcs_mat1_3_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_10833, new_AGEMA_signal_10832, mcs1_mcs_mat1_3_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9121, new_AGEMA_signal_9120, mcs1_mcs_mat1_3_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_11797, new_AGEMA_signal_11796, mcs1_mcs_mat1_3_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_11799, new_AGEMA_signal_11798, mcs1_mcs_mat1_3_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_9865, new_AGEMA_signal_9864, mcs1_mcs_mat1_3_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_12625, new_AGEMA_signal_12624, mcs1_mcs_mat1_3_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_10833, new_AGEMA_signal_10832, mcs1_mcs_mat1_3_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .c ({new_AGEMA_signal_11799, new_AGEMA_signal_11798, mcs1_mcs_mat1_3_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_10833, new_AGEMA_signal_10832, mcs1_mcs_mat1_3_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9863, new_AGEMA_signal_9862, mcs1_mcs_mat1_3_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_11801, new_AGEMA_signal_11800, mcs1_mcs_mat1_3_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_9867, new_AGEMA_signal_9866, mcs1_mcs_mat1_3_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_8343, new_AGEMA_signal_8342, mcs1_mcs_mat1_3_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_10833, new_AGEMA_signal_10832, mcs1_mcs_mat1_3_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_9119, new_AGEMA_signal_9118, mcs1_mcs_mat1_3_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_9865, new_AGEMA_signal_9864, mcs1_mcs_mat1_3_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_10835, new_AGEMA_signal_10834, mcs1_mcs_mat1_3_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_7795, new_AGEMA_signal_7794, mcs1_mcs_mat1_3_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_9121, new_AGEMA_signal_9120, mcs1_mcs_mat1_3_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_9865, new_AGEMA_signal_9864, mcs1_mcs_mat1_3_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_8343, new_AGEMA_signal_8342, mcs1_mcs_mat1_3_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_9119, new_AGEMA_signal_9118, mcs1_mcs_mat1_3_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2111], Fresh[2110], Fresh[2109]}), .c ({new_AGEMA_signal_9867, new_AGEMA_signal_9866, mcs1_mcs_mat1_3_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({new_AGEMA_signal_8343, new_AGEMA_signal_8342, mcs1_mcs_mat1_3_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2117], Fresh[2116], Fresh[2115]}), .c ({new_AGEMA_signal_9121, new_AGEMA_signal_9120, mcs1_mcs_mat1_3_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_10839, new_AGEMA_signal_10838, mcs1_mcs_mat1_3_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_8345, new_AGEMA_signal_8344, mcs1_mcs_mat1_3_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_11803, new_AGEMA_signal_11802, mcs1_mcs_mat1_3_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_9123, new_AGEMA_signal_9122, mcs1_mcs_mat1_3_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_9125, new_AGEMA_signal_9124, mcs1_mcs_mat1_3_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_9869, new_AGEMA_signal_9868, mcs1_mcs_mat1_3_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_10841, new_AGEMA_signal_10840, mcs1_mcs_mat1_3_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_11805, new_AGEMA_signal_11804, mcs1_mcs_mat1_3_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_12627, new_AGEMA_signal_12626, mcs1_mcs_mat1_3_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_10839, new_AGEMA_signal_10838, mcs1_mcs_mat1_3_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_11805, new_AGEMA_signal_11804, mcs1_mcs_mat1_3_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_7797, new_AGEMA_signal_7796, mcs1_mcs_mat1_3_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9873, new_AGEMA_signal_9872, mcs1_mcs_mat1_3_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_10839, new_AGEMA_signal_10838, mcs1_mcs_mat1_3_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_8347, new_AGEMA_signal_8346, mcs1_mcs_mat1_3_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_9871, new_AGEMA_signal_9870, mcs1_mcs_mat1_3_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_10841, new_AGEMA_signal_10840, mcs1_mcs_mat1_3_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({new_AGEMA_signal_9873, new_AGEMA_signal_9872, mcs1_mcs_mat1_3_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2123], Fresh[2122], Fresh[2121]}), .c ({new_AGEMA_signal_8347, new_AGEMA_signal_8346, mcs1_mcs_mat1_3_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({new_AGEMA_signal_9125, new_AGEMA_signal_9124, mcs1_mcs_mat1_3_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({new_AGEMA_signal_11807, new_AGEMA_signal_11806, mcs1_mcs_mat1_3_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12629, new_AGEMA_signal_12628, mcs1_mcs_mat1_3_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({new_AGEMA_signal_11809, new_AGEMA_signal_11808, mcs1_mcs_mat1_3_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12631, new_AGEMA_signal_12630, mcs1_mcs_mat1_3_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_9127, new_AGEMA_signal_9126, mcs1_mcs_mat1_3_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_11807, new_AGEMA_signal_11806, mcs1_mcs_mat1_3_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12633, new_AGEMA_signal_12632, mcs1_mcs_mat1_3_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_8349, new_AGEMA_signal_8348, mcs1_mcs_mat1_3_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_10843, new_AGEMA_signal_10842, mcs1_mcs_mat1_3_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_11807, new_AGEMA_signal_11806, mcs1_mcs_mat1_3_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_9875, new_AGEMA_signal_9874, mcs1_mcs_mat1_3_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_11809, new_AGEMA_signal_11808, mcs1_mcs_mat1_3_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12635, new_AGEMA_signal_12634, mcs1_mcs_mat1_3_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_10845, new_AGEMA_signal_10844, mcs1_mcs_mat1_3_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_11809, new_AGEMA_signal_11808, mcs1_mcs_mat1_3_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_9127, new_AGEMA_signal_9126, mcs1_mcs_mat1_3_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_9877, new_AGEMA_signal_9876, mcs1_mcs_mat1_3_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_10845, new_AGEMA_signal_10844, mcs1_mcs_mat1_3_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2129], Fresh[2128], Fresh[2127]}), .c ({new_AGEMA_signal_9877, new_AGEMA_signal_9876, mcs1_mcs_mat1_3_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({new_AGEMA_signal_8349, new_AGEMA_signal_8348, mcs1_mcs_mat1_3_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2135], Fresh[2134], Fresh[2133]}), .c ({new_AGEMA_signal_9127, new_AGEMA_signal_9126, mcs1_mcs_mat1_3_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_14145, new_AGEMA_signal_14144, mcs1_mcs_mat1_3_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_14143, new_AGEMA_signal_14142, mcs1_mcs_mat1_3_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_14579, new_AGEMA_signal_14578, mcs1_mcs_mat1_3_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_14143, new_AGEMA_signal_14142, mcs1_mcs_mat1_3_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_13217, new_AGEMA_signal_13216, mcs1_mcs_mat1_3_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_14581, new_AGEMA_signal_14580, mcs1_mcs_mat1_3_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_11811, new_AGEMA_signal_11810, mcs1_mcs_mat1_3_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .c ({new_AGEMA_signal_13217, new_AGEMA_signal_13216, mcs1_mcs_mat1_3_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_14143, new_AGEMA_signal_14142, mcs1_mcs_mat1_3_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_14583, new_AGEMA_signal_14582, mcs1_mcs_mat1_3_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_13687, new_AGEMA_signal_13686, mcs1_mcs_mat1_3_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_10847, new_AGEMA_signal_10846, mcs1_mcs_mat1_3_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_14143, new_AGEMA_signal_14142, mcs1_mcs_mat1_3_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_14585, new_AGEMA_signal_14584, mcs1_mcs_mat1_3_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_15073, new_AGEMA_signal_15072, mcs1_mcs_mat1_3_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_14145, new_AGEMA_signal_14144, mcs1_mcs_mat1_3_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_13687, new_AGEMA_signal_13686, mcs1_mcs_mat1_3_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_14585, new_AGEMA_signal_14584, mcs1_mcs_mat1_3_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_13685, new_AGEMA_signal_13684, mcs1_mcs_mat1_3_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .c ({new_AGEMA_signal_14145, new_AGEMA_signal_14144, mcs1_mcs_mat1_3_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_11811, new_AGEMA_signal_11810, mcs1_mcs_mat1_3_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_13219, new_AGEMA_signal_13218, mcs1_mcs_mat1_3_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_13685, new_AGEMA_signal_13684, mcs1_mcs_mat1_3_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({new_AGEMA_signal_13687, new_AGEMA_signal_13686, mcs1_mcs_mat1_3_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2141], Fresh[2140], Fresh[2139]}), .c ({new_AGEMA_signal_11811, new_AGEMA_signal_11810, mcs1_mcs_mat1_3_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({new_AGEMA_signal_13219, new_AGEMA_signal_13218, mcs1_mcs_mat1_3_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_9129, new_AGEMA_signal_9128, mcs1_mcs_mat1_3_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_10849, new_AGEMA_signal_10848, mcs1_mcs_mat1_3_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_11813, new_AGEMA_signal_11812, mcs1_mcs_mat1_3_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_9885, new_AGEMA_signal_9884, mcs1_mcs_mat1_3_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_10849, new_AGEMA_signal_10848, mcs1_mcs_mat1_3_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_9881, new_AGEMA_signal_9880, mcs1_mcs_mat1_3_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_9131, new_AGEMA_signal_9130, mcs1_mcs_mat1_3_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_10851, new_AGEMA_signal_10850, mcs1_mcs_mat1_3_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_9883, new_AGEMA_signal_9882, mcs1_mcs_mat1_3_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_10853, new_AGEMA_signal_10852, mcs1_mcs_mat1_3_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_11815, new_AGEMA_signal_11814, mcs1_mcs_mat1_3_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_7801, new_AGEMA_signal_7800, mcs1_mcs_mat1_3_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_9885, new_AGEMA_signal_9884, mcs1_mcs_mat1_3_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_10853, new_AGEMA_signal_10852, mcs1_mcs_mat1_3_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_8351, new_AGEMA_signal_8350, mcs1_mcs_mat1_3_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .c ({new_AGEMA_signal_9883, new_AGEMA_signal_9882, mcs1_mcs_mat1_3_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2147], Fresh[2146], Fresh[2145]}), .c ({new_AGEMA_signal_9885, new_AGEMA_signal_9884, mcs1_mcs_mat1_3_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({new_AGEMA_signal_8351, new_AGEMA_signal_8350, mcs1_mcs_mat1_3_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2153], Fresh[2152], Fresh[2151]}), .c ({new_AGEMA_signal_9131, new_AGEMA_signal_9130, mcs1_mcs_mat1_3_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, mcs1_mcs_mat1_3_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_9135, new_AGEMA_signal_9134, mcs1_mcs_mat1_3_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_13689, new_AGEMA_signal_13688, mcs1_mcs_mat1_3_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_12637, new_AGEMA_signal_12636, mcs1_mcs_mat1_3_mcs_out[99]}), .b ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .c ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, mcs1_mcs_mat1_3_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_11817, new_AGEMA_signal_11816, mcs1_mcs_mat1_3_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .c ({new_AGEMA_signal_12637, new_AGEMA_signal_12636, mcs1_mcs_mat1_3_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_10855, new_AGEMA_signal_10854, mcs1_mcs_mat1_3_mcs_out[98]}), .b ({new_AGEMA_signal_8355, new_AGEMA_signal_8354, mcs1_mcs_mat1_3_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_11817, new_AGEMA_signal_11816, mcs1_mcs_mat1_3_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_8353, new_AGEMA_signal_8352, mcs1_mcs_mat1_3_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_9887, new_AGEMA_signal_9886, mcs1_mcs_mat1_3_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_10855, new_AGEMA_signal_10854, mcs1_mcs_mat1_3_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({new_AGEMA_signal_9887, new_AGEMA_signal_9886, mcs1_mcs_mat1_3_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2159], Fresh[2158], Fresh[2157]}), .c ({new_AGEMA_signal_8355, new_AGEMA_signal_8354, mcs1_mcs_mat1_3_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({new_AGEMA_signal_9135, new_AGEMA_signal_9134, mcs1_mcs_mat1_3_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_10857, new_AGEMA_signal_10856, mcs1_mcs_mat1_3_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_11819, new_AGEMA_signal_11818, mcs1_mcs_mat1_3_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_9139, new_AGEMA_signal_9138, mcs1_mcs_mat1_3_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_9141, new_AGEMA_signal_9140, mcs1_mcs_mat1_3_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_9891, new_AGEMA_signal_9890, mcs1_mcs_mat1_3_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_11821, new_AGEMA_signal_11820, mcs1_mcs_mat1_3_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_8357, new_AGEMA_signal_8356, mcs1_mcs_mat1_3_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_12639, new_AGEMA_signal_12638, mcs1_mcs_mat1_3_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_10857, new_AGEMA_signal_10856, mcs1_mcs_mat1_3_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_11821, new_AGEMA_signal_11820, mcs1_mcs_mat1_3_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_7805, new_AGEMA_signal_7804, mcs1_mcs_mat1_3_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_9893, new_AGEMA_signal_9892, mcs1_mcs_mat1_3_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_10857, new_AGEMA_signal_10856, mcs1_mcs_mat1_3_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2165], Fresh[2164], Fresh[2163]}), .c ({new_AGEMA_signal_9893, new_AGEMA_signal_9892, mcs1_mcs_mat1_3_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({new_AGEMA_signal_8357, new_AGEMA_signal_8356, mcs1_mcs_mat1_3_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2171], Fresh[2170], Fresh[2169]}), .c ({new_AGEMA_signal_9141, new_AGEMA_signal_9140, mcs1_mcs_mat1_3_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_9901, new_AGEMA_signal_9900, mcs1_mcs_mat1_3_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_9903, new_AGEMA_signal_9902, mcs1_mcs_mat1_3_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_10861, new_AGEMA_signal_10860, mcs1_mcs_mat1_3_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_9897, new_AGEMA_signal_9896, mcs1_mcs_mat1_3_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_7807, new_AGEMA_signal_7806, mcs1_mcs_mat1_3_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_10863, new_AGEMA_signal_10862, mcs1_mcs_mat1_3_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_9143, new_AGEMA_signal_9142, mcs1_mcs_mat1_3_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_9897, new_AGEMA_signal_9896, mcs1_mcs_mat1_3_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_9899, new_AGEMA_signal_9898, mcs1_mcs_mat1_3_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_10865, new_AGEMA_signal_10864, mcs1_mcs_mat1_3_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_8359, new_AGEMA_signal_8358, mcs1_mcs_mat1_3_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_9143, new_AGEMA_signal_9142, mcs1_mcs_mat1_3_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_9899, new_AGEMA_signal_9898, mcs1_mcs_mat1_3_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_10867, new_AGEMA_signal_10866, mcs1_mcs_mat1_3_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .c ({new_AGEMA_signal_11823, new_AGEMA_signal_11822, mcs1_mcs_mat1_3_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_9901, new_AGEMA_signal_9900, mcs1_mcs_mat1_3_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_8359, new_AGEMA_signal_8358, mcs1_mcs_mat1_3_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_10867, new_AGEMA_signal_10866, mcs1_mcs_mat1_3_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({new_AGEMA_signal_9903, new_AGEMA_signal_9902, mcs1_mcs_mat1_3_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2177], Fresh[2176], Fresh[2175]}), .c ({new_AGEMA_signal_8359, new_AGEMA_signal_8358, mcs1_mcs_mat1_3_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({new_AGEMA_signal_9143, new_AGEMA_signal_9142, mcs1_mcs_mat1_3_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_10869, new_AGEMA_signal_10868, mcs1_mcs_mat1_3_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_11825, new_AGEMA_signal_11824, mcs1_mcs_mat1_3_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_9145, new_AGEMA_signal_9144, mcs1_mcs_mat1_3_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_9905, new_AGEMA_signal_9904, mcs1_mcs_mat1_3_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_11827, new_AGEMA_signal_11826, mcs1_mcs_mat1_3_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_8363, new_AGEMA_signal_8362, mcs1_mcs_mat1_3_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_12641, new_AGEMA_signal_12640, mcs1_mcs_mat1_3_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_10869, new_AGEMA_signal_10868, mcs1_mcs_mat1_3_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .c ({new_AGEMA_signal_11827, new_AGEMA_signal_11826, mcs1_mcs_mat1_3_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_7809, new_AGEMA_signal_7808, mcs1_mcs_mat1_3_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_9907, new_AGEMA_signal_9906, mcs1_mcs_mat1_3_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_10869, new_AGEMA_signal_10868, mcs1_mcs_mat1_3_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2183], Fresh[2182], Fresh[2181]}), .c ({new_AGEMA_signal_9907, new_AGEMA_signal_9906, mcs1_mcs_mat1_3_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({new_AGEMA_signal_8363, new_AGEMA_signal_8362, mcs1_mcs_mat1_3_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2189], Fresh[2188], Fresh[2187]}), .c ({new_AGEMA_signal_9145, new_AGEMA_signal_9144, mcs1_mcs_mat1_3_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_14587, new_AGEMA_signal_14586, mcs1_mcs_mat1_3_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_15075, new_AGEMA_signal_15074, mcs1_mcs_mat1_3_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_14149, new_AGEMA_signal_14148, mcs1_mcs_mat1_3_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_13693, new_AGEMA_signal_13692, mcs1_mcs_mat1_3_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_14587, new_AGEMA_signal_14586, mcs1_mcs_mat1_3_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_12643, new_AGEMA_signal_12642, mcs1_mcs_mat1_3_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_13691, new_AGEMA_signal_13690, mcs1_mcs_mat1_3_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_13693, new_AGEMA_signal_13692, mcs1_mcs_mat1_3_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_12643, new_AGEMA_signal_12642, mcs1_mcs_mat1_3_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_14147, new_AGEMA_signal_14146, mcs1_mcs_mat1_3_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_11829, new_AGEMA_signal_11828, mcs1_mcs_mat1_3_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_11831, new_AGEMA_signal_11830, mcs1_mcs_mat1_3_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_12643, new_AGEMA_signal_12642, mcs1_mcs_mat1_3_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, mcs1_mcs_mat1_3_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .c ({new_AGEMA_signal_13693, new_AGEMA_signal_13692, mcs1_mcs_mat1_3_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_14589, new_AGEMA_signal_14588, mcs1_mcs_mat1_3_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_11829, new_AGEMA_signal_11828, mcs1_mcs_mat1_3_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_15077, new_AGEMA_signal_15076, mcs1_mcs_mat1_3_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_14149, new_AGEMA_signal_14148, mcs1_mcs_mat1_3_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, mcs1_mcs_mat1_3_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_14589, new_AGEMA_signal_14588, mcs1_mcs_mat1_3_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .b ({new_AGEMA_signal_13695, new_AGEMA_signal_13694, mcs1_mcs_mat1_3_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_14149, new_AGEMA_signal_14148, mcs1_mcs_mat1_3_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({new_AGEMA_signal_13695, new_AGEMA_signal_13694, mcs1_mcs_mat1_3_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2195], Fresh[2194], Fresh[2193]}), .c ({new_AGEMA_signal_11831, new_AGEMA_signal_11830, mcs1_mcs_mat1_3_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, mcs1_mcs_mat1_3_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_10873, new_AGEMA_signal_10872, mcs1_mcs_mat1_3_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_9147, new_AGEMA_signal_9146, mcs1_mcs_mat1_3_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_11833, new_AGEMA_signal_11832, mcs1_mcs_mat1_3_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_9911, new_AGEMA_signal_9910, mcs1_mcs_mat1_3_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_11835, new_AGEMA_signal_11834, mcs1_mcs_mat1_3_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12645, new_AGEMA_signal_12644, mcs1_mcs_mat1_3_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_10873, new_AGEMA_signal_10872, mcs1_mcs_mat1_3_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_11835, new_AGEMA_signal_11834, mcs1_mcs_mat1_3_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12647, new_AGEMA_signal_12646, mcs1_mcs_mat1_3_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_9147, new_AGEMA_signal_9146, mcs1_mcs_mat1_3_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_10875, new_AGEMA_signal_10874, mcs1_mcs_mat1_3_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_11835, new_AGEMA_signal_11834, mcs1_mcs_mat1_3_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, mcs1_mcs_mat1_3_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_9147, new_AGEMA_signal_9146, mcs1_mcs_mat1_3_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_9909, new_AGEMA_signal_9908, mcs1_mcs_mat1_3_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .c ({new_AGEMA_signal_10873, new_AGEMA_signal_10872, mcs1_mcs_mat1_3_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_9149, new_AGEMA_signal_9148, mcs1_mcs_mat1_3_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7811, new_AGEMA_signal_7810, mcs1_mcs_mat1_3_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_9909, new_AGEMA_signal_9908, mcs1_mcs_mat1_3_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_10875, new_AGEMA_signal_10874, mcs1_mcs_mat1_3_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_9911, new_AGEMA_signal_9910, mcs1_mcs_mat1_3_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_11837, new_AGEMA_signal_11836, mcs1_mcs_mat1_3_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_9149, new_AGEMA_signal_9148, mcs1_mcs_mat1_3_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_9911, new_AGEMA_signal_9910, mcs1_mcs_mat1_3_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({new_AGEMA_signal_9913, new_AGEMA_signal_9912, mcs1_mcs_mat1_3_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_10875, new_AGEMA_signal_10874, mcs1_mcs_mat1_3_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2201], Fresh[2200], Fresh[2199]}), .c ({new_AGEMA_signal_9913, new_AGEMA_signal_9912, mcs1_mcs_mat1_3_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, mcs1_mcs_mat1_3_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2207], Fresh[2206], Fresh[2205]}), .c ({new_AGEMA_signal_9149, new_AGEMA_signal_9148, mcs1_mcs_mat1_3_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_11841, new_AGEMA_signal_11840, mcs1_mcs_mat1_3_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_12649, new_AGEMA_signal_12648, mcs1_mcs_mat1_3_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({new_AGEMA_signal_10877, new_AGEMA_signal_10876, mcs1_mcs_mat1_3_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_11839, new_AGEMA_signal_11838, mcs1_mcs_mat1_3_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_12651, new_AGEMA_signal_12650, mcs1_mcs_mat1_3_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_9151, new_AGEMA_signal_9150, mcs1_mcs_mat1_3_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_13229, new_AGEMA_signal_13228, mcs1_mcs_mat1_3_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_11841, new_AGEMA_signal_11840, mcs1_mcs_mat1_3_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .c ({new_AGEMA_signal_12651, new_AGEMA_signal_12650, mcs1_mcs_mat1_3_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_8367, new_AGEMA_signal_8366, mcs1_mcs_mat1_3_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_10877, new_AGEMA_signal_10876, mcs1_mcs_mat1_3_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_11841, new_AGEMA_signal_11840, mcs1_mcs_mat1_3_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_7813, new_AGEMA_signal_7812, mcs1_mcs_mat1_3_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_9917, new_AGEMA_signal_9916, mcs1_mcs_mat1_3_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_10877, new_AGEMA_signal_10876, mcs1_mcs_mat1_3_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({new_AGEMA_signal_9917, new_AGEMA_signal_9916, mcs1_mcs_mat1_3_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2213], Fresh[2212], Fresh[2211]}), .c ({new_AGEMA_signal_8367, new_AGEMA_signal_8366, mcs1_mcs_mat1_3_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({new_AGEMA_signal_9151, new_AGEMA_signal_9150, mcs1_mcs_mat1_3_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_10883, new_AGEMA_signal_10882, mcs1_mcs_mat1_3_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_9153, new_AGEMA_signal_9152, mcs1_mcs_mat1_3_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_11843, new_AGEMA_signal_11842, mcs1_mcs_mat1_3_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_8369, new_AGEMA_signal_8368, mcs1_mcs_mat1_3_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_9919, new_AGEMA_signal_9918, mcs1_mcs_mat1_3_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_10879, new_AGEMA_signal_10878, mcs1_mcs_mat1_3_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({new_AGEMA_signal_9921, new_AGEMA_signal_9920, mcs1_mcs_mat1_3_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_10881, new_AGEMA_signal_10880, mcs1_mcs_mat1_3_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2219], Fresh[2218], Fresh[2217]}), .c ({new_AGEMA_signal_9921, new_AGEMA_signal_9920, mcs1_mcs_mat1_3_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({new_AGEMA_signal_8369, new_AGEMA_signal_8368, mcs1_mcs_mat1_3_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2225], Fresh[2224], Fresh[2223]}), .c ({new_AGEMA_signal_9153, new_AGEMA_signal_9152, mcs1_mcs_mat1_3_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_11849, new_AGEMA_signal_11848, mcs1_mcs_mat1_3_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_13231, new_AGEMA_signal_13230, mcs1_mcs_mat1_3_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_13697, new_AGEMA_signal_13696, mcs1_mcs_mat1_3_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_11851, new_AGEMA_signal_11850, mcs1_mcs_mat1_3_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_13699, new_AGEMA_signal_13698, mcs1_mcs_mat1_3_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_14153, new_AGEMA_signal_14152, mcs1_mcs_mat1_3_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_14155, new_AGEMA_signal_14154, mcs1_mcs_mat1_3_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_13701, new_AGEMA_signal_13700, mcs1_mcs_mat1_3_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_14591, new_AGEMA_signal_14590, mcs1_mcs_mat1_3_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_13703, new_AGEMA_signal_13702, mcs1_mcs_mat1_3_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_14155, new_AGEMA_signal_14154, mcs1_mcs_mat1_3_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({new_AGEMA_signal_13703, new_AGEMA_signal_13702, mcs1_mcs_mat1_3_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2231], Fresh[2230], Fresh[2229]}), .c ({new_AGEMA_signal_11851, new_AGEMA_signal_11850, mcs1_mcs_mat1_3_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({new_AGEMA_signal_13231, new_AGEMA_signal_13230, mcs1_mcs_mat1_3_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_9925, new_AGEMA_signal_9924, mcs1_mcs_mat1_3_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_10887, new_AGEMA_signal_10886, mcs1_mcs_mat1_3_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_11853, new_AGEMA_signal_11852, mcs1_mcs_mat1_3_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_11855, new_AGEMA_signal_11854, mcs1_mcs_mat1_3_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_9923, new_AGEMA_signal_9922, mcs1_mcs_mat1_3_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_12655, new_AGEMA_signal_12654, mcs1_mcs_mat1_3_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_9155, new_AGEMA_signal_9154, mcs1_mcs_mat1_3_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_9923, new_AGEMA_signal_9922, mcs1_mcs_mat1_3_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({new_AGEMA_signal_11855, new_AGEMA_signal_11854, mcs1_mcs_mat1_3_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_12657, new_AGEMA_signal_12656, mcs1_mcs_mat1_3_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_7817, new_AGEMA_signal_7816, mcs1_mcs_mat1_3_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_10887, new_AGEMA_signal_10886, mcs1_mcs_mat1_3_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_11855, new_AGEMA_signal_11854, mcs1_mcs_mat1_3_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, mcs1_mcs_mat1_3_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_9929, new_AGEMA_signal_9928, mcs1_mcs_mat1_3_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_10887, new_AGEMA_signal_10886, mcs1_mcs_mat1_3_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_9927, new_AGEMA_signal_9926, mcs1_mcs_mat1_3_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_10889, new_AGEMA_signal_10888, mcs1_mcs_mat1_3_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_11857, new_AGEMA_signal_11856, mcs1_mcs_mat1_3_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_9925, new_AGEMA_signal_9924, mcs1_mcs_mat1_3_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, mcs1_mcs_mat1_3_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_10889, new_AGEMA_signal_10888, mcs1_mcs_mat1_3_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_9155, new_AGEMA_signal_9154, mcs1_mcs_mat1_3_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_9925, new_AGEMA_signal_9924, mcs1_mcs_mat1_3_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2237], Fresh[2236], Fresh[2235]}), .c ({new_AGEMA_signal_9929, new_AGEMA_signal_9928, mcs1_mcs_mat1_3_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, mcs1_mcs_mat1_3_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2243], Fresh[2242], Fresh[2241]}), .c ({new_AGEMA_signal_9155, new_AGEMA_signal_9154, mcs1_mcs_mat1_3_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_9159, new_AGEMA_signal_9158, mcs1_mcs_mat1_3_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_9933, new_AGEMA_signal_9932, mcs1_mcs_mat1_3_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_12659, new_AGEMA_signal_12658, mcs1_mcs_mat1_3_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_8373, new_AGEMA_signal_8372, mcs1_mcs_mat1_3_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, mcs1_mcs_mat1_3_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_11859, new_AGEMA_signal_11858, mcs1_mcs_mat1_3_mcs_out[47]}), .b ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_12659, new_AGEMA_signal_12658, mcs1_mcs_mat1_3_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_10893, new_AGEMA_signal_10892, mcs1_mcs_mat1_3_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .c ({new_AGEMA_signal_11859, new_AGEMA_signal_11858, mcs1_mcs_mat1_3_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_7819, new_AGEMA_signal_7818, mcs1_mcs_mat1_3_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_9935, new_AGEMA_signal_9934, mcs1_mcs_mat1_3_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_10893, new_AGEMA_signal_10892, mcs1_mcs_mat1_3_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({new_AGEMA_signal_9935, new_AGEMA_signal_9934, mcs1_mcs_mat1_3_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2249], Fresh[2248], Fresh[2247]}), .c ({new_AGEMA_signal_8373, new_AGEMA_signal_8372, mcs1_mcs_mat1_3_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({new_AGEMA_signal_9159, new_AGEMA_signal_9158, mcs1_mcs_mat1_3_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_14157, new_AGEMA_signal_14156, mcs1_mcs_mat1_3_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_13235, new_AGEMA_signal_13234, mcs1_mcs_mat1_3_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_14593, new_AGEMA_signal_14592, mcs1_mcs_mat1_3_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_13705, new_AGEMA_signal_13704, mcs1_mcs_mat1_3_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_11861, new_AGEMA_signal_11860, mcs1_mcs_mat1_3_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_14157, new_AGEMA_signal_14156, mcs1_mcs_mat1_3_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_14159, new_AGEMA_signal_14158, mcs1_mcs_mat1_3_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_13709, new_AGEMA_signal_13708, mcs1_mcs_mat1_3_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_14595, new_AGEMA_signal_14594, mcs1_mcs_mat1_3_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_14161, new_AGEMA_signal_14160, mcs1_mcs_mat1_3_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_10895, new_AGEMA_signal_10894, mcs1_mcs_mat1_3_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_14597, new_AGEMA_signal_14596, mcs1_mcs_mat1_3_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_13705, new_AGEMA_signal_13704, mcs1_mcs_mat1_3_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_13237, new_AGEMA_signal_13236, mcs1_mcs_mat1_3_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_14161, new_AGEMA_signal_14160, mcs1_mcs_mat1_3_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_13707, new_AGEMA_signal_13706, mcs1_mcs_mat1_3_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_13237, new_AGEMA_signal_13236, mcs1_mcs_mat1_3_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_14163, new_AGEMA_signal_14162, mcs1_mcs_mat1_3_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2255], Fresh[2254], Fresh[2253]}), .c ({new_AGEMA_signal_13709, new_AGEMA_signal_13708, mcs1_mcs_mat1_3_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({new_AGEMA_signal_11861, new_AGEMA_signal_11860, mcs1_mcs_mat1_3_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2261], Fresh[2260], Fresh[2259]}), .c ({new_AGEMA_signal_13237, new_AGEMA_signal_13236, mcs1_mcs_mat1_3_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_11863, new_AGEMA_signal_11862, mcs1_mcs_mat1_3_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_7821, new_AGEMA_signal_7820, mcs1_mcs_mat1_3_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_12661, new_AGEMA_signal_12660, mcs1_mcs_mat1_3_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_9163, new_AGEMA_signal_9162, mcs1_mcs_mat1_3_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_9161, new_AGEMA_signal_9160, mcs1_mcs_mat1_3_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_9937, new_AGEMA_signal_9936, mcs1_mcs_mat1_3_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({new_AGEMA_signal_11863, new_AGEMA_signal_11862, mcs1_mcs_mat1_3_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, mcs1_mcs_mat1_3_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_9939, new_AGEMA_signal_9938, mcs1_mcs_mat1_3_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_10897, new_AGEMA_signal_10896, mcs1_mcs_mat1_3_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_11863, new_AGEMA_signal_11862, mcs1_mcs_mat1_3_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_9941, new_AGEMA_signal_9940, mcs1_mcs_mat1_3_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9165, new_AGEMA_signal_9164, mcs1_mcs_mat1_3_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_10897, new_AGEMA_signal_10896, mcs1_mcs_mat1_3_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_9941, new_AGEMA_signal_9940, mcs1_mcs_mat1_3_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9163, new_AGEMA_signal_9162, mcs1_mcs_mat1_3_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_10899, new_AGEMA_signal_10898, mcs1_mcs_mat1_3_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_8785, new_AGEMA_signal_8784, mcs1_mcs_mat1_3_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_9163, new_AGEMA_signal_9162, mcs1_mcs_mat1_3_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({new_AGEMA_signal_8375, new_AGEMA_signal_8374, mcs1_mcs_mat1_3_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_8785, new_AGEMA_signal_8784, mcs1_mcs_mat1_3_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({new_AGEMA_signal_9941, new_AGEMA_signal_9940, mcs1_mcs_mat1_3_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2267], Fresh[2266], Fresh[2265]}), .c ({new_AGEMA_signal_8375, new_AGEMA_signal_8374, mcs1_mcs_mat1_3_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({new_AGEMA_signal_9165, new_AGEMA_signal_9164, mcs1_mcs_mat1_3_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_9943, new_AGEMA_signal_9942, mcs1_mcs_mat1_3_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_9167, new_AGEMA_signal_9166, mcs1_mcs_mat1_3_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_10901, new_AGEMA_signal_10900, mcs1_mcs_mat1_3_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, mcs1_mcs_mat1_3_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_8787, new_AGEMA_signal_8786, mcs1_mcs_mat1_3_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_12665, new_AGEMA_signal_12664, mcs1_mcs_mat1_3_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_9945, new_AGEMA_signal_9944, mcs1_mcs_mat1_3_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, mcs1_mcs_mat1_3_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2273], Fresh[2272], Fresh[2271]}), .c ({new_AGEMA_signal_9945, new_AGEMA_signal_9944, mcs1_mcs_mat1_3_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, mcs1_mcs_mat1_3_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2279], Fresh[2278], Fresh[2277]}), .c ({new_AGEMA_signal_9167, new_AGEMA_signal_9166, mcs1_mcs_mat1_3_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_11867, new_AGEMA_signal_11866, mcs1_mcs_mat1_3_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_10905, new_AGEMA_signal_10904, mcs1_mcs_mat1_3_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_12667, new_AGEMA_signal_12666, mcs1_mcs_mat1_3_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_8381, new_AGEMA_signal_8380, mcs1_mcs_mat1_3_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_10907, new_AGEMA_signal_10906, mcs1_mcs_mat1_3_mcs_out[29]}), .c ({new_AGEMA_signal_11867, new_AGEMA_signal_11866, mcs1_mcs_mat1_3_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_8379, new_AGEMA_signal_8378, mcs1_mcs_mat1_3_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_10905, new_AGEMA_signal_10904, mcs1_mcs_mat1_3_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_11869, new_AGEMA_signal_11868, mcs1_mcs_mat1_3_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_9951, new_AGEMA_signal_9950, mcs1_mcs_mat1_3_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .c ({new_AGEMA_signal_10905, new_AGEMA_signal_10904, mcs1_mcs_mat1_3_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_11871, new_AGEMA_signal_11870, mcs1_mcs_mat1_3_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_9947, new_AGEMA_signal_9946, mcs1_mcs_mat1_3_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_12669, new_AGEMA_signal_12668, mcs1_mcs_mat1_3_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_10909, new_AGEMA_signal_10908, mcs1_mcs_mat1_3_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_9949, new_AGEMA_signal_9948, mcs1_mcs_mat1_3_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_11871, new_AGEMA_signal_11870, mcs1_mcs_mat1_3_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_9169, new_AGEMA_signal_9168, mcs1_mcs_mat1_3_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_9949, new_AGEMA_signal_9948, mcs1_mcs_mat1_3_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_9951, new_AGEMA_signal_9950, mcs1_mcs_mat1_3_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8381, new_AGEMA_signal_8380, mcs1_mcs_mat1_3_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_10909, new_AGEMA_signal_10908, mcs1_mcs_mat1_3_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({new_AGEMA_signal_9951, new_AGEMA_signal_9950, mcs1_mcs_mat1_3_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2285], Fresh[2284], Fresh[2283]}), .c ({new_AGEMA_signal_8381, new_AGEMA_signal_8380, mcs1_mcs_mat1_3_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({new_AGEMA_signal_9169, new_AGEMA_signal_9168, mcs1_mcs_mat1_3_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_13711, new_AGEMA_signal_13710, mcs1_mcs_mat1_3_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_14165, new_AGEMA_signal_14164, mcs1_mcs_mat1_3_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_13241, new_AGEMA_signal_13240, mcs1_mcs_mat1_3_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_11873, new_AGEMA_signal_11872, mcs1_mcs_mat1_3_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_13711, new_AGEMA_signal_13710, mcs1_mcs_mat1_3_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_14167, new_AGEMA_signal_14166, mcs1_mcs_mat1_3_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_14599, new_AGEMA_signal_14598, mcs1_mcs_mat1_3_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_13715, new_AGEMA_signal_13714, mcs1_mcs_mat1_3_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_11873, new_AGEMA_signal_11872, mcs1_mcs_mat1_3_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_14167, new_AGEMA_signal_14166, mcs1_mcs_mat1_3_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_14601, new_AGEMA_signal_14600, mcs1_mcs_mat1_3_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .c ({new_AGEMA_signal_15079, new_AGEMA_signal_15078, mcs1_mcs_mat1_3_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_13715, new_AGEMA_signal_13714, mcs1_mcs_mat1_3_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_14169, new_AGEMA_signal_14168, mcs1_mcs_mat1_3_mcs_out[24]}), .c ({new_AGEMA_signal_14601, new_AGEMA_signal_14600, mcs1_mcs_mat1_3_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_13713, new_AGEMA_signal_13712, mcs1_mcs_mat1_3_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .c ({new_AGEMA_signal_14169, new_AGEMA_signal_14168, mcs1_mcs_mat1_3_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_13241, new_AGEMA_signal_13240, mcs1_mcs_mat1_3_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_10911, new_AGEMA_signal_10910, mcs1_mcs_mat1_3_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_13713, new_AGEMA_signal_13712, mcs1_mcs_mat1_3_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2291], Fresh[2290], Fresh[2289]}), .c ({new_AGEMA_signal_13715, new_AGEMA_signal_13714, mcs1_mcs_mat1_3_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({new_AGEMA_signal_11873, new_AGEMA_signal_11872, mcs1_mcs_mat1_3_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2297], Fresh[2296], Fresh[2295]}), .c ({new_AGEMA_signal_13241, new_AGEMA_signal_13240, mcs1_mcs_mat1_3_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_9953, new_AGEMA_signal_9952, mcs1_mcs_mat1_3_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .c ({new_AGEMA_signal_10913, new_AGEMA_signal_10912, mcs1_mcs_mat1_3_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_9171, new_AGEMA_signal_9170, mcs1_mcs_mat1_3_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, mcs1_mcs_mat1_3_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_9953, new_AGEMA_signal_9952, mcs1_mcs_mat1_3_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_10915, new_AGEMA_signal_10914, mcs1_mcs_mat1_3_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .c ({new_AGEMA_signal_11875, new_AGEMA_signal_11874, mcs1_mcs_mat1_3_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_9957, new_AGEMA_signal_9956, mcs1_mcs_mat1_3_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, mcs1_mcs_mat1_3_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_10915, new_AGEMA_signal_10914, mcs1_mcs_mat1_3_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_11877, new_AGEMA_signal_11876, mcs1_mcs_mat1_3_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_12671, new_AGEMA_signal_12670, mcs1_mcs_mat1_3_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_9957, new_AGEMA_signal_9956, mcs1_mcs_mat1_3_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_10917, new_AGEMA_signal_10916, mcs1_mcs_mat1_3_mcs_out[20]}), .c ({new_AGEMA_signal_11877, new_AGEMA_signal_11876, mcs1_mcs_mat1_3_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_9955, new_AGEMA_signal_9954, mcs1_mcs_mat1_3_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_10917, new_AGEMA_signal_10916, mcs1_mcs_mat1_3_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_9171, new_AGEMA_signal_9170, mcs1_mcs_mat1_3_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7827, new_AGEMA_signal_7826, mcs1_mcs_mat1_3_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_9955, new_AGEMA_signal_9954, mcs1_mcs_mat1_3_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({new_AGEMA_signal_9957, new_AGEMA_signal_9956, mcs1_mcs_mat1_3_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2303], Fresh[2302], Fresh[2301]}), .c ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, mcs1_mcs_mat1_3_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({new_AGEMA_signal_9171, new_AGEMA_signal_9170, mcs1_mcs_mat1_3_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_9959, new_AGEMA_signal_9958, mcs1_mcs_mat1_3_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_9965, new_AGEMA_signal_9964, mcs1_mcs_mat1_3_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_10919, new_AGEMA_signal_10918, mcs1_mcs_mat1_3_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_10921, new_AGEMA_signal_10920, mcs1_mcs_mat1_3_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_7829, new_AGEMA_signal_7828, mcs1_mcs_mat1_3_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_11879, new_AGEMA_signal_11878, mcs1_mcs_mat1_3_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_11881, new_AGEMA_signal_11880, mcs1_mcs_mat1_3_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_8385, new_AGEMA_signal_8384, mcs1_mcs_mat1_3_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_12673, new_AGEMA_signal_12672, mcs1_mcs_mat1_3_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_10921, new_AGEMA_signal_10920, mcs1_mcs_mat1_3_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_11881, new_AGEMA_signal_11880, mcs1_mcs_mat1_3_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_9961, new_AGEMA_signal_9960, mcs1_mcs_mat1_3_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .c ({new_AGEMA_signal_10921, new_AGEMA_signal_10920, mcs1_mcs_mat1_3_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_9173, new_AGEMA_signal_9172, mcs1_mcs_mat1_3_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_9175, new_AGEMA_signal_9174, mcs1_mcs_mat1_3_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_9961, new_AGEMA_signal_9960, mcs1_mcs_mat1_3_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_9963, new_AGEMA_signal_9962, mcs1_mcs_mat1_3_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_8385, new_AGEMA_signal_8384, mcs1_mcs_mat1_3_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_10923, new_AGEMA_signal_10922, mcs1_mcs_mat1_3_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2309], Fresh[2308], Fresh[2307]}), .c ({new_AGEMA_signal_9965, new_AGEMA_signal_9964, mcs1_mcs_mat1_3_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({new_AGEMA_signal_8385, new_AGEMA_signal_8384, mcs1_mcs_mat1_3_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2315], Fresh[2314], Fresh[2313]}), .c ({new_AGEMA_signal_9175, new_AGEMA_signal_9174, mcs1_mcs_mat1_3_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_11887, new_AGEMA_signal_11886, mcs1_mcs_mat1_3_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_8789, new_AGEMA_signal_8788, mcs1_mcs_mat1_3_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_12675, new_AGEMA_signal_12674, mcs1_mcs_mat1_3_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_10929, new_AGEMA_signal_10928, mcs1_mcs_mat1_3_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_10925, new_AGEMA_signal_10924, mcs1_mcs_mat1_3_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_11883, new_AGEMA_signal_11882, mcs1_mcs_mat1_3_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_9969, new_AGEMA_signal_9968, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_8387, new_AGEMA_signal_8386, mcs1_mcs_mat1_3_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_10925, new_AGEMA_signal_10924, mcs1_mcs_mat1_3_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_8789, new_AGEMA_signal_8788, mcs1_mcs_mat1_3_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_10927, new_AGEMA_signal_10926, mcs1_mcs_mat1_3_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_11885, new_AGEMA_signal_11884, mcs1_mcs_mat1_3_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_9967, new_AGEMA_signal_9966, mcs1_mcs_mat1_3_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_9969, new_AGEMA_signal_9968, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_10927, new_AGEMA_signal_10926, mcs1_mcs_mat1_3_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_7831, new_AGEMA_signal_7830, mcs1_mcs_mat1_3_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_8387, new_AGEMA_signal_8386, mcs1_mcs_mat1_3_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8789, new_AGEMA_signal_8788, mcs1_mcs_mat1_3_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_12677, new_AGEMA_signal_12676, mcs1_mcs_mat1_3_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_13243, new_AGEMA_signal_13242, mcs1_mcs_mat1_3_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_11887, new_AGEMA_signal_11886, mcs1_mcs_mat1_3_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_9969, new_AGEMA_signal_9968, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_12677, new_AGEMA_signal_12676, mcs1_mcs_mat1_3_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_10929, new_AGEMA_signal_10928, mcs1_mcs_mat1_3_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_11887, new_AGEMA_signal_11886, mcs1_mcs_mat1_3_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_9967, new_AGEMA_signal_9966, mcs1_mcs_mat1_3_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_10929, new_AGEMA_signal_10928, mcs1_mcs_mat1_3_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, shiftr_out[112]}), .b ({new_AGEMA_signal_9177, new_AGEMA_signal_9176, mcs1_mcs_mat1_3_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_9967, new_AGEMA_signal_9966, mcs1_mcs_mat1_3_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({new_AGEMA_signal_9969, new_AGEMA_signal_9968, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2321], Fresh[2320], Fresh[2319]}), .c ({new_AGEMA_signal_8387, new_AGEMA_signal_8386, mcs1_mcs_mat1_3_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({new_AGEMA_signal_9177, new_AGEMA_signal_9176, mcs1_mcs_mat1_3_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_12679, new_AGEMA_signal_12678, mcs1_mcs_mat1_3_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .c ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, mcs1_mcs_mat1_3_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_14173, new_AGEMA_signal_14172, mcs1_mcs_mat1_3_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_14603, new_AGEMA_signal_14602, mcs1_mcs_mat1_3_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_13717, new_AGEMA_signal_13716, mcs1_mcs_mat1_3_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_14171, new_AGEMA_signal_14170, mcs1_mcs_mat1_3_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_13247, new_AGEMA_signal_13246, mcs1_mcs_mat1_3_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_12679, new_AGEMA_signal_12678, mcs1_mcs_mat1_3_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_13717, new_AGEMA_signal_13716, mcs1_mcs_mat1_3_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_10931, new_AGEMA_signal_10930, mcs1_mcs_mat1_3_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_11889, new_AGEMA_signal_11888, mcs1_mcs_mat1_3_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_12679, new_AGEMA_signal_12678, mcs1_mcs_mat1_3_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_14605, new_AGEMA_signal_14604, mcs1_mcs_mat1_3_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_9503, new_AGEMA_signal_9502, shiftr_out[80]}), .c ({new_AGEMA_signal_15081, new_AGEMA_signal_15080, mcs1_mcs_mat1_3_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_10931, new_AGEMA_signal_10930, mcs1_mcs_mat1_3_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_14173, new_AGEMA_signal_14172, mcs1_mcs_mat1_3_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_14605, new_AGEMA_signal_14604, mcs1_mcs_mat1_3_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_13719, new_AGEMA_signal_13718, mcs1_mcs_mat1_3_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_13247, new_AGEMA_signal_13246, mcs1_mcs_mat1_3_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_14173, new_AGEMA_signal_14172, mcs1_mcs_mat1_3_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2327], Fresh[2326], Fresh[2325]}), .c ({new_AGEMA_signal_13719, new_AGEMA_signal_13718, mcs1_mcs_mat1_3_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10463, new_AGEMA_signal_10462, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({new_AGEMA_signal_11889, new_AGEMA_signal_11888, mcs1_mcs_mat1_3_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, shiftr_out[83]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2333], Fresh[2332], Fresh[2331]}), .c ({new_AGEMA_signal_13247, new_AGEMA_signal_13246, mcs1_mcs_mat1_3_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_13249, new_AGEMA_signal_13248, mcs1_mcs_mat1_3_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_9181, new_AGEMA_signal_9180, mcs1_mcs_mat1_3_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_13721, new_AGEMA_signal_13720, mcs1_mcs_mat1_3_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_12681, new_AGEMA_signal_12680, mcs1_mcs_mat1_3_mcs_out[7]}), .b ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .c ({new_AGEMA_signal_13249, new_AGEMA_signal_13248, mcs1_mcs_mat1_3_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_11891, new_AGEMA_signal_11890, mcs1_mcs_mat1_3_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .c ({new_AGEMA_signal_12681, new_AGEMA_signal_12680, mcs1_mcs_mat1_3_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_10933, new_AGEMA_signal_10932, mcs1_mcs_mat1_3_mcs_out[6]}), .b ({new_AGEMA_signal_8391, new_AGEMA_signal_8390, mcs1_mcs_mat1_3_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_11891, new_AGEMA_signal_11890, mcs1_mcs_mat1_3_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, mcs1_mcs_mat1_3_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_9971, new_AGEMA_signal_9970, mcs1_mcs_mat1_3_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_10933, new_AGEMA_signal_10932, mcs1_mcs_mat1_3_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, shiftr_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({new_AGEMA_signal_9971, new_AGEMA_signal_9970, mcs1_mcs_mat1_3_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, shiftr_out[50]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2339], Fresh[2338], Fresh[2337]}), .c ({new_AGEMA_signal_8391, new_AGEMA_signal_8390, mcs1_mcs_mat1_3_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({new_AGEMA_signal_9181, new_AGEMA_signal_9180, mcs1_mcs_mat1_3_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_9183, new_AGEMA_signal_9182, mcs1_mcs_mat1_3_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_9973, new_AGEMA_signal_9972, mcs1_mcs_mat1_3_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_10937, new_AGEMA_signal_10936, mcs1_mcs_mat1_3_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .b ({new_AGEMA_signal_9185, new_AGEMA_signal_9184, mcs1_mcs_mat1_3_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_9973, new_AGEMA_signal_9972, mcs1_mcs_mat1_3_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_10939, new_AGEMA_signal_10938, mcs1_mcs_mat1_3_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_8393, new_AGEMA_signal_8392, mcs1_mcs_mat1_3_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_11893, new_AGEMA_signal_11892, mcs1_mcs_mat1_3_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_10941, new_AGEMA_signal_10940, mcs1_mcs_mat1_3_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_9977, new_AGEMA_signal_9976, mcs1_mcs_mat1_3_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_11895, new_AGEMA_signal_11894, mcs1_mcs_mat1_3_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_9979, new_AGEMA_signal_9978, mcs1_mcs_mat1_3_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_7835, new_AGEMA_signal_7834, mcs1_mcs_mat1_3_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_10941, new_AGEMA_signal_10940, mcs1_mcs_mat1_3_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, shiftr_out[17]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2345], Fresh[2344], Fresh[2343]}), .c ({new_AGEMA_signal_9979, new_AGEMA_signal_9978, mcs1_mcs_mat1_3_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, shiftr_out[18]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({new_AGEMA_signal_8393, new_AGEMA_signal_8392, mcs1_mcs_mat1_3_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2351], Fresh[2350], Fresh[2349]}), .c ({new_AGEMA_signal_9185, new_AGEMA_signal_9184, mcs1_mcs_mat1_3_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U96 ( .a ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, mcs1_mcs_mat1_4_n128}), .b ({new_AGEMA_signal_14175, new_AGEMA_signal_14174, mcs1_mcs_mat1_4_n127}), .c ({temp_next_s2[77], temp_next_s1[77], temp_next_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U95 ( .a ({new_AGEMA_signal_11983, new_AGEMA_signal_11982, mcs1_mcs_mat1_4_mcs_out[41]}), .b ({new_AGEMA_signal_13759, new_AGEMA_signal_13758, mcs1_mcs_mat1_4_mcs_out[45]}), .c ({new_AGEMA_signal_14175, new_AGEMA_signal_14174, mcs1_mcs_mat1_4_n127}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U94 ( .a ({new_AGEMA_signal_8795, new_AGEMA_signal_8794, mcs1_mcs_mat1_4_mcs_out[33]}), .b ({new_AGEMA_signal_12731, new_AGEMA_signal_12730, mcs1_mcs_mat1_4_mcs_out[37]}), .c ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, mcs1_mcs_mat1_4_n128}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U93 ( .a ({new_AGEMA_signal_13723, new_AGEMA_signal_13722, mcs1_mcs_mat1_4_n126}), .b ({new_AGEMA_signal_16071, new_AGEMA_signal_16070, mcs1_mcs_mat1_4_n125}), .c ({temp_next_s2[76], temp_next_s1[76], temp_next_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U92 ( .a ({new_AGEMA_signal_11017, new_AGEMA_signal_11016, mcs1_mcs_mat1_4_mcs_out[40]}), .b ({new_AGEMA_signal_15657, new_AGEMA_signal_15656, mcs1_mcs_mat1_4_mcs_out[44]}), .c ({new_AGEMA_signal_16071, new_AGEMA_signal_16070, mcs1_mcs_mat1_4_n125}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U91 ( .a ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, mcs1_mcs_mat1_4_mcs_out[32]}), .b ({new_AGEMA_signal_11021, new_AGEMA_signal_11020, mcs1_mcs_mat1_4_mcs_out[36]}), .c ({new_AGEMA_signal_13723, new_AGEMA_signal_13722, mcs1_mcs_mat1_4_n126}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U90 ( .a ({new_AGEMA_signal_11897, new_AGEMA_signal_11896, mcs1_mcs_mat1_4_n124}), .b ({new_AGEMA_signal_15623, new_AGEMA_signal_15622, mcs1_mcs_mat1_4_n123}), .c ({temp_next_s2[47], temp_next_s1[47], temp_next_s0[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U89 ( .a ({new_AGEMA_signal_11029, new_AGEMA_signal_11028, mcs1_mcs_mat1_4_mcs_out[27]}), .b ({new_AGEMA_signal_15119, new_AGEMA_signal_15118, mcs1_mcs_mat1_4_mcs_out[31]}), .c ({new_AGEMA_signal_15623, new_AGEMA_signal_15622, mcs1_mcs_mat1_4_n123}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U88 ( .a ({new_AGEMA_signal_11041, new_AGEMA_signal_11040, mcs1_mcs_mat1_4_mcs_out[19]}), .b ({new_AGEMA_signal_11035, new_AGEMA_signal_11034, mcs1_mcs_mat1_4_mcs_out[23]}), .c ({new_AGEMA_signal_11897, new_AGEMA_signal_11896, mcs1_mcs_mat1_4_n124}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U87 ( .a ({new_AGEMA_signal_12683, new_AGEMA_signal_12682, mcs1_mcs_mat1_4_n122}), .b ({new_AGEMA_signal_15083, new_AGEMA_signal_15082, mcs1_mcs_mat1_4_n121}), .c ({temp_next_s2[46], temp_next_s1[46], temp_next_s0[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U86 ( .a ({new_AGEMA_signal_11993, new_AGEMA_signal_11992, mcs1_mcs_mat1_4_mcs_out[26]}), .b ({new_AGEMA_signal_14641, new_AGEMA_signal_14640, mcs1_mcs_mat1_4_mcs_out[30]}), .c ({new_AGEMA_signal_15083, new_AGEMA_signal_15082, mcs1_mcs_mat1_4_n121}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U85 ( .a ({new_AGEMA_signal_12001, new_AGEMA_signal_12000, mcs1_mcs_mat1_4_mcs_out[18]}), .b ({new_AGEMA_signal_11997, new_AGEMA_signal_11996, mcs1_mcs_mat1_4_mcs_out[22]}), .c ({new_AGEMA_signal_12683, new_AGEMA_signal_12682, mcs1_mcs_mat1_4_n122}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U84 ( .a ({new_AGEMA_signal_13253, new_AGEMA_signal_13252, mcs1_mcs_mat1_4_n120}), .b ({new_AGEMA_signal_14609, new_AGEMA_signal_14608, mcs1_mcs_mat1_4_n119}), .c ({temp_next_s2[45], temp_next_s1[45], temp_next_s0[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U83 ( .a ({new_AGEMA_signal_12735, new_AGEMA_signal_12734, mcs1_mcs_mat1_4_mcs_out[25]}), .b ({new_AGEMA_signal_14209, new_AGEMA_signal_14208, mcs1_mcs_mat1_4_mcs_out[29]}), .c ({new_AGEMA_signal_14609, new_AGEMA_signal_14608, mcs1_mcs_mat1_4_n119}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U82 ( .a ({new_AGEMA_signal_12739, new_AGEMA_signal_12738, mcs1_mcs_mat1_4_mcs_out[17]}), .b ({new_AGEMA_signal_12737, new_AGEMA_signal_12736, mcs1_mcs_mat1_4_mcs_out[21]}), .c ({new_AGEMA_signal_13253, new_AGEMA_signal_13252, mcs1_mcs_mat1_4_n120}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U81 ( .a ({new_AGEMA_signal_11899, new_AGEMA_signal_11898, mcs1_mcs_mat1_4_n118}), .b ({new_AGEMA_signal_15627, new_AGEMA_signal_15626, mcs1_mcs_mat1_4_n117}), .c ({temp_next_s2[44], temp_next_s1[44], temp_next_s0[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U80 ( .a ({new_AGEMA_signal_11033, new_AGEMA_signal_11032, mcs1_mcs_mat1_4_mcs_out[24]}), .b ({new_AGEMA_signal_15121, new_AGEMA_signal_15120, mcs1_mcs_mat1_4_mcs_out[28]}), .c ({new_AGEMA_signal_15627, new_AGEMA_signal_15626, mcs1_mcs_mat1_4_n117}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U79 ( .a ({new_AGEMA_signal_11045, new_AGEMA_signal_11044, mcs1_mcs_mat1_4_mcs_out[16]}), .b ({new_AGEMA_signal_11039, new_AGEMA_signal_11038, mcs1_mcs_mat1_4_mcs_out[20]}), .c ({new_AGEMA_signal_11899, new_AGEMA_signal_11898, mcs1_mcs_mat1_4_n118}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U78 ( .a ({new_AGEMA_signal_15629, new_AGEMA_signal_15628, mcs1_mcs_mat1_4_n116}), .b ({new_AGEMA_signal_13255, new_AGEMA_signal_13254, mcs1_mcs_mat1_4_n115}), .c ({temp_next_s2[15], temp_next_s1[15], temp_next_s0[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U77 ( .a ({new_AGEMA_signal_11055, new_AGEMA_signal_11054, mcs1_mcs_mat1_4_mcs_out[3]}), .b ({new_AGEMA_signal_12745, new_AGEMA_signal_12744, mcs1_mcs_mat1_4_mcs_out[7]}), .c ({new_AGEMA_signal_13255, new_AGEMA_signal_13254, mcs1_mcs_mat1_4_n115}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U76 ( .a ({new_AGEMA_signal_9251, new_AGEMA_signal_9250, mcs1_mcs_mat1_4_mcs_out[11]}), .b ({new_AGEMA_signal_15123, new_AGEMA_signal_15122, mcs1_mcs_mat1_4_mcs_out[15]}), .c ({new_AGEMA_signal_15629, new_AGEMA_signal_15628, mcs1_mcs_mat1_4_n116}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U75 ( .a ({new_AGEMA_signal_13259, new_AGEMA_signal_13258, mcs1_mcs_mat1_4_n114}), .b ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, mcs1_mcs_mat1_4_n113}), .c ({new_AGEMA_signal_13725, new_AGEMA_signal_13724, mcs_out[239]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U74 ( .a ({new_AGEMA_signal_12699, new_AGEMA_signal_12698, mcs1_mcs_mat1_4_mcs_out[123]}), .b ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, mcs1_mcs_mat1_4_n113}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U73 ( .a ({new_AGEMA_signal_11925, new_AGEMA_signal_11924, mcs1_mcs_mat1_4_mcs_out[115]}), .b ({new_AGEMA_signal_12703, new_AGEMA_signal_12702, mcs1_mcs_mat1_4_mcs_out[119]}), .c ({new_AGEMA_signal_13259, new_AGEMA_signal_13258, mcs1_mcs_mat1_4_n114}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U72 ( .a ({new_AGEMA_signal_13261, new_AGEMA_signal_13260, mcs1_mcs_mat1_4_n112}), .b ({new_AGEMA_signal_13727, new_AGEMA_signal_13726, mcs1_mcs_mat1_4_n111}), .c ({new_AGEMA_signal_14177, new_AGEMA_signal_14176, mcs_out[238]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U71 ( .a ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, mcs1_mcs_mat1_4_mcs_out[122]}), .b ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_13727, new_AGEMA_signal_13726, mcs1_mcs_mat1_4_n111}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U70 ( .a ({new_AGEMA_signal_10951, new_AGEMA_signal_10950, mcs1_mcs_mat1_4_mcs_out[114]}), .b ({new_AGEMA_signal_12705, new_AGEMA_signal_12704, mcs1_mcs_mat1_4_mcs_out[118]}), .c ({new_AGEMA_signal_13261, new_AGEMA_signal_13260, mcs1_mcs_mat1_4_n112}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U69 ( .a ({new_AGEMA_signal_15087, new_AGEMA_signal_15086, mcs1_mcs_mat1_4_n110}), .b ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, mcs1_mcs_mat1_4_n109}), .c ({temp_next_s2[14], temp_next_s1[14], temp_next_s0[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U68 ( .a ({new_AGEMA_signal_11057, new_AGEMA_signal_11056, mcs1_mcs_mat1_4_mcs_out[2]}), .b ({new_AGEMA_signal_11053, new_AGEMA_signal_11052, mcs1_mcs_mat1_4_mcs_out[6]}), .c ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, mcs1_mcs_mat1_4_n109}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U67 ( .a ({new_AGEMA_signal_12007, new_AGEMA_signal_12006, mcs1_mcs_mat1_4_mcs_out[10]}), .b ({new_AGEMA_signal_14645, new_AGEMA_signal_14644, mcs1_mcs_mat1_4_mcs_out[14]}), .c ({new_AGEMA_signal_15087, new_AGEMA_signal_15086, mcs1_mcs_mat1_4_n110}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U66 ( .a ({new_AGEMA_signal_12685, new_AGEMA_signal_12684, mcs1_mcs_mat1_4_n108}), .b ({new_AGEMA_signal_13729, new_AGEMA_signal_13728, mcs1_mcs_mat1_4_n107}), .c ({new_AGEMA_signal_14179, new_AGEMA_signal_14178, mcs_out[237]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U65 ( .a ({new_AGEMA_signal_12701, new_AGEMA_signal_12700, mcs1_mcs_mat1_4_mcs_out[121]}), .b ({new_AGEMA_signal_13283, new_AGEMA_signal_13282, mcs1_mcs_mat1_4_mcs_out[125]}), .c ({new_AGEMA_signal_13729, new_AGEMA_signal_13728, mcs1_mcs_mat1_4_n107}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U64 ( .a ({new_AGEMA_signal_9991, new_AGEMA_signal_9990, mcs1_mcs_mat1_4_mcs_out[113]}), .b ({new_AGEMA_signal_11923, new_AGEMA_signal_11922, mcs1_mcs_mat1_4_mcs_out[117]}), .c ({new_AGEMA_signal_12685, new_AGEMA_signal_12684, mcs1_mcs_mat1_4_n108}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U63 ( .a ({new_AGEMA_signal_13265, new_AGEMA_signal_13264, mcs1_mcs_mat1_4_n106}), .b ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, mcs1_mcs_mat1_4_n105}), .c ({new_AGEMA_signal_13731, new_AGEMA_signal_13730, mcs_out[236]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U62 ( .a ({new_AGEMA_signal_11917, new_AGEMA_signal_11916, mcs1_mcs_mat1_4_mcs_out[120]}), .b ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, mcs1_mcs_mat1_4_n105}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U61 ( .a ({new_AGEMA_signal_12707, new_AGEMA_signal_12706, mcs1_mcs_mat1_4_mcs_out[112]}), .b ({new_AGEMA_signal_10949, new_AGEMA_signal_10948, mcs1_mcs_mat1_4_mcs_out[116]}), .c ({new_AGEMA_signal_13265, new_AGEMA_signal_13264, mcs1_mcs_mat1_4_n106}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U60 ( .a ({new_AGEMA_signal_12687, new_AGEMA_signal_12686, mcs1_mcs_mat1_4_n104}), .b ({new_AGEMA_signal_15633, new_AGEMA_signal_15632, mcs1_mcs_mat1_4_n103}), .c ({new_AGEMA_signal_16079, new_AGEMA_signal_16078, mcs_out[207]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U59 ( .a ({new_AGEMA_signal_15103, new_AGEMA_signal_15102, mcs1_mcs_mat1_4_mcs_out[111]}), .b ({new_AGEMA_signal_12711, new_AGEMA_signal_12710, mcs1_mcs_mat1_4_mcs_out[99]}), .c ({new_AGEMA_signal_15633, new_AGEMA_signal_15632, mcs1_mcs_mat1_4_n103}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U58 ( .a ({new_AGEMA_signal_11939, new_AGEMA_signal_11938, mcs1_mcs_mat1_4_mcs_out[103]}), .b ({new_AGEMA_signal_11931, new_AGEMA_signal_11930, mcs1_mcs_mat1_4_mcs_out[107]}), .c ({new_AGEMA_signal_12687, new_AGEMA_signal_12686, mcs1_mcs_mat1_4_n104}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U57 ( .a ({new_AGEMA_signal_12689, new_AGEMA_signal_12688, mcs1_mcs_mat1_4_n102}), .b ({new_AGEMA_signal_15635, new_AGEMA_signal_15634, mcs1_mcs_mat1_4_n101}), .c ({new_AGEMA_signal_16081, new_AGEMA_signal_16080, mcs_out[206]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U56 ( .a ({new_AGEMA_signal_15105, new_AGEMA_signal_15104, mcs1_mcs_mat1_4_mcs_out[110]}), .b ({new_AGEMA_signal_10969, new_AGEMA_signal_10968, mcs1_mcs_mat1_4_mcs_out[98]}), .c ({new_AGEMA_signal_15635, new_AGEMA_signal_15634, mcs1_mcs_mat1_4_n101}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U55 ( .a ({new_AGEMA_signal_10001, new_AGEMA_signal_10000, mcs1_mcs_mat1_4_mcs_out[102]}), .b ({new_AGEMA_signal_11933, new_AGEMA_signal_11932, mcs1_mcs_mat1_4_mcs_out[106]}), .c ({new_AGEMA_signal_12689, new_AGEMA_signal_12688, mcs1_mcs_mat1_4_n102}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U54 ( .a ({new_AGEMA_signal_12691, new_AGEMA_signal_12690, mcs1_mcs_mat1_4_n100}), .b ({new_AGEMA_signal_15637, new_AGEMA_signal_15636, mcs1_mcs_mat1_4_n99}), .c ({new_AGEMA_signal_16083, new_AGEMA_signal_16082, mcs_out[205]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U53 ( .a ({new_AGEMA_signal_15107, new_AGEMA_signal_15106, mcs1_mcs_mat1_4_mcs_out[109]}), .b ({new_AGEMA_signal_9209, new_AGEMA_signal_9208, mcs1_mcs_mat1_4_mcs_out[97]}), .c ({new_AGEMA_signal_15637, new_AGEMA_signal_15636, mcs1_mcs_mat1_4_n99}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U52 ( .a ({new_AGEMA_signal_10965, new_AGEMA_signal_10964, mcs1_mcs_mat1_4_mcs_out[101]}), .b ({new_AGEMA_signal_11935, new_AGEMA_signal_11934, mcs1_mcs_mat1_4_mcs_out[105]}), .c ({new_AGEMA_signal_12691, new_AGEMA_signal_12690, mcs1_mcs_mat1_4_n100}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U51 ( .a ({new_AGEMA_signal_13267, new_AGEMA_signal_13266, mcs1_mcs_mat1_4_n98}), .b ({new_AGEMA_signal_15639, new_AGEMA_signal_15638, mcs1_mcs_mat1_4_n97}), .c ({new_AGEMA_signal_16085, new_AGEMA_signal_16084, mcs_out[204]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U50 ( .a ({new_AGEMA_signal_15109, new_AGEMA_signal_15108, mcs1_mcs_mat1_4_mcs_out[108]}), .b ({new_AGEMA_signal_13743, new_AGEMA_signal_13742, mcs1_mcs_mat1_4_mcs_out[96]}), .c ({new_AGEMA_signal_15639, new_AGEMA_signal_15638, mcs1_mcs_mat1_4_n97}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U49 ( .a ({new_AGEMA_signal_11941, new_AGEMA_signal_11940, mcs1_mcs_mat1_4_mcs_out[100]}), .b ({new_AGEMA_signal_12709, new_AGEMA_signal_12708, mcs1_mcs_mat1_4_mcs_out[104]}), .c ({new_AGEMA_signal_13267, new_AGEMA_signal_13266, mcs1_mcs_mat1_4_n98}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U48 ( .a ({new_AGEMA_signal_11903, new_AGEMA_signal_11902, mcs1_mcs_mat1_4_n96}), .b ({new_AGEMA_signal_15089, new_AGEMA_signal_15088, mcs1_mcs_mat1_4_n95}), .c ({new_AGEMA_signal_15641, new_AGEMA_signal_15640, mcs_out[175]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U47 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_14625, new_AGEMA_signal_14624, mcs1_mcs_mat1_4_mcs_out[95]}), .c ({new_AGEMA_signal_15089, new_AGEMA_signal_15088, mcs1_mcs_mat1_4_n95}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U46 ( .a ({new_AGEMA_signal_10975, new_AGEMA_signal_10974, mcs1_mcs_mat1_4_mcs_out[83]}), .b ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, mcs1_mcs_mat1_4_mcs_out[87]}), .c ({new_AGEMA_signal_11903, new_AGEMA_signal_11902, mcs1_mcs_mat1_4_n96}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U45 ( .a ({new_AGEMA_signal_11905, new_AGEMA_signal_11904, mcs1_mcs_mat1_4_n94}), .b ({new_AGEMA_signal_14181, new_AGEMA_signal_14180, mcs1_mcs_mat1_4_n93}), .c ({new_AGEMA_signal_14611, new_AGEMA_signal_14610, mcs_out[174]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U43 ( .a ({new_AGEMA_signal_10977, new_AGEMA_signal_10976, mcs1_mcs_mat1_4_mcs_out[82]}), .b ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_11905, new_AGEMA_signal_11904, mcs1_mcs_mat1_4_n94}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U42 ( .a ({new_AGEMA_signal_11907, new_AGEMA_signal_11906, mcs1_mcs_mat1_4_n92}), .b ({new_AGEMA_signal_14183, new_AGEMA_signal_14182, mcs1_mcs_mat1_4_n91}), .c ({new_AGEMA_signal_14613, new_AGEMA_signal_14612, mcs_out[173]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U41 ( .a ({new_AGEMA_signal_9215, new_AGEMA_signal_9214, mcs1_mcs_mat1_4_mcs_out[89]}), .b ({new_AGEMA_signal_13747, new_AGEMA_signal_13746, mcs1_mcs_mat1_4_mcs_out[93]}), .c ({new_AGEMA_signal_14183, new_AGEMA_signal_14182, mcs1_mcs_mat1_4_n91}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U40 ( .a ({new_AGEMA_signal_10979, new_AGEMA_signal_10978, mcs1_mcs_mat1_4_mcs_out[81]}), .b ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_11907, new_AGEMA_signal_11906, mcs1_mcs_mat1_4_n92}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U39 ( .a ({new_AGEMA_signal_12693, new_AGEMA_signal_12692, mcs1_mcs_mat1_4_n90}), .b ({new_AGEMA_signal_15643, new_AGEMA_signal_15642, mcs1_mcs_mat1_4_n89}), .c ({new_AGEMA_signal_16087, new_AGEMA_signal_16086, mcs_out[172]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U38 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_15111, new_AGEMA_signal_15110, mcs1_mcs_mat1_4_mcs_out[92]}), .c ({new_AGEMA_signal_15643, new_AGEMA_signal_15642, mcs1_mcs_mat1_4_n89}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U37 ( .a ({new_AGEMA_signal_11947, new_AGEMA_signal_11946, mcs1_mcs_mat1_4_mcs_out[80]}), .b ({new_AGEMA_signal_10973, new_AGEMA_signal_10972, mcs1_mcs_mat1_4_mcs_out[84]}), .c ({new_AGEMA_signal_12693, new_AGEMA_signal_12692, mcs1_mcs_mat1_4_n90}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U36 ( .a ({new_AGEMA_signal_15091, new_AGEMA_signal_15090, mcs1_mcs_mat1_4_n88}), .b ({new_AGEMA_signal_11909, new_AGEMA_signal_11908, mcs1_mcs_mat1_4_n87}), .c ({temp_next_s2[13], temp_next_s1[13], temp_next_s0[13]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U35 ( .a ({new_AGEMA_signal_9255, new_AGEMA_signal_9254, mcs1_mcs_mat1_4_mcs_out[5]}), .b ({new_AGEMA_signal_11049, new_AGEMA_signal_11048, mcs1_mcs_mat1_4_mcs_out[9]}), .c ({new_AGEMA_signal_11909, new_AGEMA_signal_11908, mcs1_mcs_mat1_4_n87}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U34 ( .a ({new_AGEMA_signal_14647, new_AGEMA_signal_14646, mcs1_mcs_mat1_4_mcs_out[13]}), .b ({new_AGEMA_signal_12013, new_AGEMA_signal_12012, mcs1_mcs_mat1_4_mcs_out[1]}), .c ({new_AGEMA_signal_15091, new_AGEMA_signal_15090, mcs1_mcs_mat1_4_n88}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U33 ( .a ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, mcs1_mcs_mat1_4_n86}), .b ({new_AGEMA_signal_15093, new_AGEMA_signal_15092, mcs1_mcs_mat1_4_n85}), .c ({new_AGEMA_signal_15647, new_AGEMA_signal_15646, mcs_out[143]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U32 ( .a ({new_AGEMA_signal_10021, new_AGEMA_signal_10020, mcs1_mcs_mat1_4_mcs_out[75]}), .b ({new_AGEMA_signal_14629, new_AGEMA_signal_14628, mcs1_mcs_mat1_4_mcs_out[79]}), .c ({new_AGEMA_signal_15093, new_AGEMA_signal_15092, mcs1_mcs_mat1_4_n85}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U31 ( .a ({new_AGEMA_signal_12721, new_AGEMA_signal_12720, mcs1_mcs_mat1_4_mcs_out[67]}), .b ({new_AGEMA_signal_11957, new_AGEMA_signal_11956, mcs1_mcs_mat1_4_mcs_out[71]}), .c ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, mcs1_mcs_mat1_4_n86}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U30 ( .a ({new_AGEMA_signal_13273, new_AGEMA_signal_13272, mcs1_mcs_mat1_4_n84}), .b ({new_AGEMA_signal_13271, new_AGEMA_signal_13270, mcs1_mcs_mat1_4_n83}), .c ({new_AGEMA_signal_13733, new_AGEMA_signal_13732, mcs_out[142]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U29 ( .a ({new_AGEMA_signal_12713, new_AGEMA_signal_12712, mcs1_mcs_mat1_4_mcs_out[74]}), .b ({new_AGEMA_signal_11949, new_AGEMA_signal_11948, mcs1_mcs_mat1_4_mcs_out[78]}), .c ({new_AGEMA_signal_13271, new_AGEMA_signal_13270, mcs1_mcs_mat1_4_n83}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U28 ( .a ({new_AGEMA_signal_11963, new_AGEMA_signal_11962, mcs1_mcs_mat1_4_mcs_out[66]}), .b ({new_AGEMA_signal_12717, new_AGEMA_signal_12716, mcs1_mcs_mat1_4_mcs_out[70]}), .c ({new_AGEMA_signal_13273, new_AGEMA_signal_13272, mcs1_mcs_mat1_4_n84}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U27 ( .a ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, mcs1_mcs_mat1_4_n82}), .b ({new_AGEMA_signal_14185, new_AGEMA_signal_14184, mcs1_mcs_mat1_4_n81}), .c ({new_AGEMA_signal_14615, new_AGEMA_signal_14614, mcs_out[141]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U26 ( .a ({new_AGEMA_signal_10985, new_AGEMA_signal_10984, mcs1_mcs_mat1_4_mcs_out[73]}), .b ({new_AGEMA_signal_13751, new_AGEMA_signal_13750, mcs1_mcs_mat1_4_mcs_out[77]}), .c ({new_AGEMA_signal_14185, new_AGEMA_signal_14184, mcs1_mcs_mat1_4_n81}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U25 ( .a ({new_AGEMA_signal_10033, new_AGEMA_signal_10032, mcs1_mcs_mat1_4_mcs_out[65]}), .b ({new_AGEMA_signal_12719, new_AGEMA_signal_12718, mcs1_mcs_mat1_4_mcs_out[69]}), .c ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, mcs1_mcs_mat1_4_n82}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U24 ( .a ({new_AGEMA_signal_13735, new_AGEMA_signal_13734, mcs1_mcs_mat1_4_n80}), .b ({new_AGEMA_signal_15649, new_AGEMA_signal_15648, mcs1_mcs_mat1_4_n79}), .c ({new_AGEMA_signal_16089, new_AGEMA_signal_16088, mcs_out[140]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U23 ( .a ({new_AGEMA_signal_12715, new_AGEMA_signal_12714, mcs1_mcs_mat1_4_mcs_out[72]}), .b ({new_AGEMA_signal_15113, new_AGEMA_signal_15112, mcs1_mcs_mat1_4_mcs_out[76]}), .c ({new_AGEMA_signal_15649, new_AGEMA_signal_15648, mcs1_mcs_mat1_4_n79}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U22 ( .a ({new_AGEMA_signal_13297, new_AGEMA_signal_13296, mcs1_mcs_mat1_4_mcs_out[64]}), .b ({new_AGEMA_signal_11961, new_AGEMA_signal_11960, mcs1_mcs_mat1_4_mcs_out[68]}), .c ({new_AGEMA_signal_13735, new_AGEMA_signal_13734, mcs1_mcs_mat1_4_n80}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U21 ( .a ({new_AGEMA_signal_12695, new_AGEMA_signal_12694, mcs1_mcs_mat1_4_n78}), .b ({new_AGEMA_signal_15095, new_AGEMA_signal_15094, mcs1_mcs_mat1_4_n77}), .c ({temp_next_s2[111], temp_next_s1[111], temp_next_s0[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U20 ( .a ({new_AGEMA_signal_10997, new_AGEMA_signal_10996, mcs1_mcs_mat1_4_mcs_out[59]}), .b ({new_AGEMA_signal_14633, new_AGEMA_signal_14632, mcs1_mcs_mat1_4_mcs_out[63]}), .c ({new_AGEMA_signal_15095, new_AGEMA_signal_15094, mcs1_mcs_mat1_4_n77}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U19 ( .a ({new_AGEMA_signal_10053, new_AGEMA_signal_10052, mcs1_mcs_mat1_4_mcs_out[51]}), .b ({new_AGEMA_signal_11971, new_AGEMA_signal_11970, mcs1_mcs_mat1_4_mcs_out[55]}), .c ({new_AGEMA_signal_12695, new_AGEMA_signal_12694, mcs1_mcs_mat1_4_n78}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U18 ( .a ({new_AGEMA_signal_13277, new_AGEMA_signal_13276, mcs1_mcs_mat1_4_n76}), .b ({new_AGEMA_signal_14617, new_AGEMA_signal_14616, mcs1_mcs_mat1_4_n75}), .c ({temp_next_s2[110], temp_next_s1[110], temp_next_s0[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U17 ( .a ({new_AGEMA_signal_10037, new_AGEMA_signal_10036, mcs1_mcs_mat1_4_mcs_out[58]}), .b ({new_AGEMA_signal_14199, new_AGEMA_signal_14198, mcs1_mcs_mat1_4_mcs_out[62]}), .c ({new_AGEMA_signal_14617, new_AGEMA_signal_14616, mcs1_mcs_mat1_4_n75}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U16 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_12725, new_AGEMA_signal_12724, mcs1_mcs_mat1_4_mcs_out[54]}), .c ({new_AGEMA_signal_13277, new_AGEMA_signal_13276, mcs1_mcs_mat1_4_n76}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U15 ( .a ({new_AGEMA_signal_13279, new_AGEMA_signal_13278, mcs1_mcs_mat1_4_n74}), .b ({new_AGEMA_signal_14619, new_AGEMA_signal_14618, mcs1_mcs_mat1_4_n73}), .c ({temp_next_s2[109], temp_next_s1[109], temp_next_s0[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U14 ( .a ({new_AGEMA_signal_10999, new_AGEMA_signal_10998, mcs1_mcs_mat1_4_mcs_out[57]}), .b ({new_AGEMA_signal_14201, new_AGEMA_signal_14200, mcs1_mcs_mat1_4_mcs_out[61]}), .c ({new_AGEMA_signal_14619, new_AGEMA_signal_14618, mcs1_mcs_mat1_4_n73}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U13 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_12727, new_AGEMA_signal_12726, mcs1_mcs_mat1_4_mcs_out[53]}), .c ({new_AGEMA_signal_13279, new_AGEMA_signal_13278, mcs1_mcs_mat1_4_n74}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U12 ( .a ({new_AGEMA_signal_12697, new_AGEMA_signal_12696, mcs1_mcs_mat1_4_n72}), .b ({new_AGEMA_signal_15653, new_AGEMA_signal_15652, mcs1_mcs_mat1_4_n71}), .c ({temp_next_s2[108], temp_next_s1[108], temp_next_s0[108]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U11 ( .a ({new_AGEMA_signal_11969, new_AGEMA_signal_11968, mcs1_mcs_mat1_4_mcs_out[56]}), .b ({new_AGEMA_signal_15115, new_AGEMA_signal_15114, mcs1_mcs_mat1_4_mcs_out[60]}), .c ({new_AGEMA_signal_15653, new_AGEMA_signal_15652, mcs1_mcs_mat1_4_n71}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U10 ( .a ({new_AGEMA_signal_11007, new_AGEMA_signal_11006, mcs1_mcs_mat1_4_mcs_out[48]}), .b ({new_AGEMA_signal_11975, new_AGEMA_signal_11974, mcs1_mcs_mat1_4_mcs_out[52]}), .c ({new_AGEMA_signal_12697, new_AGEMA_signal_12696, mcs1_mcs_mat1_4_n72}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U9 ( .a ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, mcs1_mcs_mat1_4_n70}), .b ({new_AGEMA_signal_15101, new_AGEMA_signal_15100, mcs1_mcs_mat1_4_n69}), .c ({temp_next_s2[79], temp_next_s1[79], temp_next_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U8 ( .a ({new_AGEMA_signal_11979, new_AGEMA_signal_11978, mcs1_mcs_mat1_4_mcs_out[43]}), .b ({new_AGEMA_signal_14637, new_AGEMA_signal_14636, mcs1_mcs_mat1_4_mcs_out[47]}), .c ({new_AGEMA_signal_15101, new_AGEMA_signal_15100, mcs1_mcs_mat1_4_n69}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U7 ( .a ({new_AGEMA_signal_11987, new_AGEMA_signal_11986, mcs1_mcs_mat1_4_mcs_out[35]}), .b ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, mcs1_mcs_mat1_4_mcs_out[39]}), .c ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, mcs1_mcs_mat1_4_n70}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U6 ( .a ({new_AGEMA_signal_11911, new_AGEMA_signal_11910, mcs1_mcs_mat1_4_n68}), .b ({new_AGEMA_signal_13737, new_AGEMA_signal_13736, mcs1_mcs_mat1_4_n67}), .c ({temp_next_s2[78], temp_next_s1[78], temp_next_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U5 ( .a ({new_AGEMA_signal_11981, new_AGEMA_signal_11980, mcs1_mcs_mat1_4_mcs_out[42]}), .b ({new_AGEMA_signal_13301, new_AGEMA_signal_13300, mcs1_mcs_mat1_4_mcs_out[46]}), .c ({new_AGEMA_signal_13737, new_AGEMA_signal_13736, mcs1_mcs_mat1_4_n67}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U4 ( .a ({new_AGEMA_signal_11023, new_AGEMA_signal_11022, mcs1_mcs_mat1_4_mcs_out[34]}), .b ({new_AGEMA_signal_10061, new_AGEMA_signal_10060, mcs1_mcs_mat1_4_mcs_out[38]}), .c ({new_AGEMA_signal_11911, new_AGEMA_signal_11910, mcs1_mcs_mat1_4_n68}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U3 ( .a ({new_AGEMA_signal_16093, new_AGEMA_signal_16092, mcs1_mcs_mat1_4_n66}), .b ({new_AGEMA_signal_14189, new_AGEMA_signal_14188, mcs1_mcs_mat1_4_n65}), .c ({temp_next_s2[12], temp_next_s1[12], temp_next_s0[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U2 ( .a ({new_AGEMA_signal_13773, new_AGEMA_signal_13772, mcs1_mcs_mat1_4_mcs_out[4]}), .b ({new_AGEMA_signal_12743, new_AGEMA_signal_12742, mcs1_mcs_mat1_4_mcs_out[8]}), .c ({new_AGEMA_signal_14189, new_AGEMA_signal_14188, mcs1_mcs_mat1_4_n65}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_U1 ( .a ({new_AGEMA_signal_12015, new_AGEMA_signal_12014, mcs1_mcs_mat1_4_mcs_out[0]}), .b ({new_AGEMA_signal_15659, new_AGEMA_signal_15658, mcs1_mcs_mat1_4_mcs_out[12]}), .c ({new_AGEMA_signal_16093, new_AGEMA_signal_16092, mcs1_mcs_mat1_4_n66}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_11913, new_AGEMA_signal_11912, mcs1_mcs_mat1_4_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_12699, new_AGEMA_signal_12698, mcs1_mcs_mat1_4_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_10943, new_AGEMA_signal_10942, mcs1_mcs_mat1_4_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_7837, new_AGEMA_signal_7836, mcs1_mcs_mat1_4_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_11913, new_AGEMA_signal_11912, mcs1_mcs_mat1_4_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, mcs1_mcs_mat1_4_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_9187, new_AGEMA_signal_9186, mcs1_mcs_mat1_4_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, mcs1_mcs_mat1_4_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_4_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .c ({new_AGEMA_signal_9187, new_AGEMA_signal_9186, mcs1_mcs_mat1_4_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_11915, new_AGEMA_signal_11914, mcs1_mcs_mat1_4_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .c ({new_AGEMA_signal_12701, new_AGEMA_signal_12700, mcs1_mcs_mat1_4_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_10943, new_AGEMA_signal_10942, mcs1_mcs_mat1_4_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_11915, new_AGEMA_signal_11914, mcs1_mcs_mat1_4_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_9983, new_AGEMA_signal_9982, mcs1_mcs_mat1_4_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9189, new_AGEMA_signal_9188, mcs1_mcs_mat1_4_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_10943, new_AGEMA_signal_10942, mcs1_mcs_mat1_4_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_10945, new_AGEMA_signal_10944, mcs1_mcs_mat1_4_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_11917, new_AGEMA_signal_11916, mcs1_mcs_mat1_4_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_9983, new_AGEMA_signal_9982, mcs1_mcs_mat1_4_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_4_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_10945, new_AGEMA_signal_10944, mcs1_mcs_mat1_4_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({new_AGEMA_signal_9983, new_AGEMA_signal_9982, mcs1_mcs_mat1_4_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2357], Fresh[2356], Fresh[2355]}), .c ({new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_4_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({new_AGEMA_signal_9189, new_AGEMA_signal_9188, mcs1_mcs_mat1_4_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_11919, new_AGEMA_signal_11918, mcs1_mcs_mat1_4_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .c ({new_AGEMA_signal_12703, new_AGEMA_signal_12702, mcs1_mcs_mat1_4_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_10947, new_AGEMA_signal_10946, mcs1_mcs_mat1_4_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9195, new_AGEMA_signal_9194, mcs1_mcs_mat1_4_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_11919, new_AGEMA_signal_11918, mcs1_mcs_mat1_4_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_11921, new_AGEMA_signal_11920, mcs1_mcs_mat1_4_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_9987, new_AGEMA_signal_9986, mcs1_mcs_mat1_4_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_12705, new_AGEMA_signal_12704, mcs1_mcs_mat1_4_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_10947, new_AGEMA_signal_10946, mcs1_mcs_mat1_4_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .c ({new_AGEMA_signal_11921, new_AGEMA_signal_11920, mcs1_mcs_mat1_4_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_10947, new_AGEMA_signal_10946, mcs1_mcs_mat1_4_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9985, new_AGEMA_signal_9984, mcs1_mcs_mat1_4_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_11923, new_AGEMA_signal_11922, mcs1_mcs_mat1_4_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_9989, new_AGEMA_signal_9988, mcs1_mcs_mat1_4_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_8399, new_AGEMA_signal_8398, mcs1_mcs_mat1_4_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_10947, new_AGEMA_signal_10946, mcs1_mcs_mat1_4_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_9193, new_AGEMA_signal_9192, mcs1_mcs_mat1_4_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_9987, new_AGEMA_signal_9986, mcs1_mcs_mat1_4_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_10949, new_AGEMA_signal_10948, mcs1_mcs_mat1_4_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_7839, new_AGEMA_signal_7838, mcs1_mcs_mat1_4_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_9195, new_AGEMA_signal_9194, mcs1_mcs_mat1_4_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_9987, new_AGEMA_signal_9986, mcs1_mcs_mat1_4_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_8399, new_AGEMA_signal_8398, mcs1_mcs_mat1_4_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_9193, new_AGEMA_signal_9192, mcs1_mcs_mat1_4_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2363], Fresh[2362], Fresh[2361]}), .c ({new_AGEMA_signal_9989, new_AGEMA_signal_9988, mcs1_mcs_mat1_4_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({new_AGEMA_signal_8399, new_AGEMA_signal_8398, mcs1_mcs_mat1_4_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2369], Fresh[2368], Fresh[2367]}), .c ({new_AGEMA_signal_9195, new_AGEMA_signal_9194, mcs1_mcs_mat1_4_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_10953, new_AGEMA_signal_10952, mcs1_mcs_mat1_4_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, mcs1_mcs_mat1_4_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_11925, new_AGEMA_signal_11924, mcs1_mcs_mat1_4_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_9197, new_AGEMA_signal_9196, mcs1_mcs_mat1_4_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_9199, new_AGEMA_signal_9198, mcs1_mcs_mat1_4_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_9991, new_AGEMA_signal_9990, mcs1_mcs_mat1_4_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_10955, new_AGEMA_signal_10954, mcs1_mcs_mat1_4_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_11927, new_AGEMA_signal_11926, mcs1_mcs_mat1_4_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_12707, new_AGEMA_signal_12706, mcs1_mcs_mat1_4_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_10953, new_AGEMA_signal_10952, mcs1_mcs_mat1_4_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_11927, new_AGEMA_signal_11926, mcs1_mcs_mat1_4_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_7841, new_AGEMA_signal_7840, mcs1_mcs_mat1_4_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_9995, new_AGEMA_signal_9994, mcs1_mcs_mat1_4_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_10953, new_AGEMA_signal_10952, mcs1_mcs_mat1_4_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, mcs1_mcs_mat1_4_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_10955, new_AGEMA_signal_10954, mcs1_mcs_mat1_4_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({new_AGEMA_signal_9995, new_AGEMA_signal_9994, mcs1_mcs_mat1_4_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2375], Fresh[2374], Fresh[2373]}), .c ({new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({new_AGEMA_signal_9199, new_AGEMA_signal_9198, mcs1_mcs_mat1_4_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({new_AGEMA_signal_14621, new_AGEMA_signal_14620, mcs1_mcs_mat1_4_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_15103, new_AGEMA_signal_15102, mcs1_mcs_mat1_4_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({new_AGEMA_signal_14623, new_AGEMA_signal_14622, mcs1_mcs_mat1_4_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_15105, new_AGEMA_signal_15104, mcs1_mcs_mat1_4_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_13285, new_AGEMA_signal_13284, mcs1_mcs_mat1_4_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_14621, new_AGEMA_signal_14620, mcs1_mcs_mat1_4_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_15107, new_AGEMA_signal_15106, mcs1_mcs_mat1_4_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_11929, new_AGEMA_signal_11928, mcs1_mcs_mat1_4_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_14191, new_AGEMA_signal_14190, mcs1_mcs_mat1_4_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_14621, new_AGEMA_signal_14620, mcs1_mcs_mat1_4_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_13739, new_AGEMA_signal_13738, mcs1_mcs_mat1_4_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_14623, new_AGEMA_signal_14622, mcs1_mcs_mat1_4_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_15109, new_AGEMA_signal_15108, mcs1_mcs_mat1_4_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_14193, new_AGEMA_signal_14192, mcs1_mcs_mat1_4_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_14623, new_AGEMA_signal_14622, mcs1_mcs_mat1_4_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_13285, new_AGEMA_signal_13284, mcs1_mcs_mat1_4_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_13741, new_AGEMA_signal_13740, mcs1_mcs_mat1_4_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_14193, new_AGEMA_signal_14192, mcs1_mcs_mat1_4_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2381], Fresh[2380], Fresh[2379]}), .c ({new_AGEMA_signal_13741, new_AGEMA_signal_13740, mcs1_mcs_mat1_4_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({new_AGEMA_signal_11929, new_AGEMA_signal_11928, mcs1_mcs_mat1_4_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2387], Fresh[2386], Fresh[2385]}), .c ({new_AGEMA_signal_13285, new_AGEMA_signal_13284, mcs1_mcs_mat1_4_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_10961, new_AGEMA_signal_10960, mcs1_mcs_mat1_4_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_10959, new_AGEMA_signal_10958, mcs1_mcs_mat1_4_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_11931, new_AGEMA_signal_11930, mcs1_mcs_mat1_4_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_10959, new_AGEMA_signal_10958, mcs1_mcs_mat1_4_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_9201, new_AGEMA_signal_9200, mcs1_mcs_mat1_4_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_11933, new_AGEMA_signal_11932, mcs1_mcs_mat1_4_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_8405, new_AGEMA_signal_8404, mcs1_mcs_mat1_4_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .c ({new_AGEMA_signal_9201, new_AGEMA_signal_9200, mcs1_mcs_mat1_4_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_10959, new_AGEMA_signal_10958, mcs1_mcs_mat1_4_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_11935, new_AGEMA_signal_11934, mcs1_mcs_mat1_4_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_9999, new_AGEMA_signal_9998, mcs1_mcs_mat1_4_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_7843, new_AGEMA_signal_7842, mcs1_mcs_mat1_4_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_10959, new_AGEMA_signal_10958, mcs1_mcs_mat1_4_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_11937, new_AGEMA_signal_11936, mcs1_mcs_mat1_4_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_12709, new_AGEMA_signal_12708, mcs1_mcs_mat1_4_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_10961, new_AGEMA_signal_10960, mcs1_mcs_mat1_4_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_9999, new_AGEMA_signal_9998, mcs1_mcs_mat1_4_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_11937, new_AGEMA_signal_11936, mcs1_mcs_mat1_4_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_9997, new_AGEMA_signal_9996, mcs1_mcs_mat1_4_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .c ({new_AGEMA_signal_10961, new_AGEMA_signal_10960, mcs1_mcs_mat1_4_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_8405, new_AGEMA_signal_8404, mcs1_mcs_mat1_4_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_9203, new_AGEMA_signal_9202, mcs1_mcs_mat1_4_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_9997, new_AGEMA_signal_9996, mcs1_mcs_mat1_4_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({new_AGEMA_signal_9999, new_AGEMA_signal_9998, mcs1_mcs_mat1_4_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2393], Fresh[2392], Fresh[2391]}), .c ({new_AGEMA_signal_8405, new_AGEMA_signal_8404, mcs1_mcs_mat1_4_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({new_AGEMA_signal_9203, new_AGEMA_signal_9202, mcs1_mcs_mat1_4_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_9205, new_AGEMA_signal_9204, mcs1_mcs_mat1_4_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_10963, new_AGEMA_signal_10962, mcs1_mcs_mat1_4_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_11939, new_AGEMA_signal_11938, mcs1_mcs_mat1_4_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_10007, new_AGEMA_signal_10006, mcs1_mcs_mat1_4_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_10963, new_AGEMA_signal_10962, mcs1_mcs_mat1_4_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_10003, new_AGEMA_signal_10002, mcs1_mcs_mat1_4_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_9207, new_AGEMA_signal_9206, mcs1_mcs_mat1_4_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_10965, new_AGEMA_signal_10964, mcs1_mcs_mat1_4_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_10005, new_AGEMA_signal_10004, mcs1_mcs_mat1_4_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_10967, new_AGEMA_signal_10966, mcs1_mcs_mat1_4_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_11941, new_AGEMA_signal_11940, mcs1_mcs_mat1_4_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_7845, new_AGEMA_signal_7844, mcs1_mcs_mat1_4_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_10007, new_AGEMA_signal_10006, mcs1_mcs_mat1_4_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_10967, new_AGEMA_signal_10966, mcs1_mcs_mat1_4_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, mcs1_mcs_mat1_4_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .c ({new_AGEMA_signal_10005, new_AGEMA_signal_10004, mcs1_mcs_mat1_4_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2399], Fresh[2398], Fresh[2397]}), .c ({new_AGEMA_signal_10007, new_AGEMA_signal_10006, mcs1_mcs_mat1_4_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, mcs1_mcs_mat1_4_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2405], Fresh[2404], Fresh[2403]}), .c ({new_AGEMA_signal_9207, new_AGEMA_signal_9206, mcs1_mcs_mat1_4_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, mcs1_mcs_mat1_4_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_9211, new_AGEMA_signal_9210, mcs1_mcs_mat1_4_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_13743, new_AGEMA_signal_13742, mcs1_mcs_mat1_4_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_12711, new_AGEMA_signal_12710, mcs1_mcs_mat1_4_mcs_out[99]}), .b ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .c ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, mcs1_mcs_mat1_4_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_11943, new_AGEMA_signal_11942, mcs1_mcs_mat1_4_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .c ({new_AGEMA_signal_12711, new_AGEMA_signal_12710, mcs1_mcs_mat1_4_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_10969, new_AGEMA_signal_10968, mcs1_mcs_mat1_4_mcs_out[98]}), .b ({new_AGEMA_signal_8411, new_AGEMA_signal_8410, mcs1_mcs_mat1_4_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_11943, new_AGEMA_signal_11942, mcs1_mcs_mat1_4_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_4_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_10009, new_AGEMA_signal_10008, mcs1_mcs_mat1_4_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_10969, new_AGEMA_signal_10968, mcs1_mcs_mat1_4_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({new_AGEMA_signal_10009, new_AGEMA_signal_10008, mcs1_mcs_mat1_4_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2411], Fresh[2410], Fresh[2409]}), .c ({new_AGEMA_signal_8411, new_AGEMA_signal_8410, mcs1_mcs_mat1_4_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({new_AGEMA_signal_9211, new_AGEMA_signal_9210, mcs1_mcs_mat1_4_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_14195, new_AGEMA_signal_14194, mcs1_mcs_mat1_4_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_14625, new_AGEMA_signal_14624, mcs1_mcs_mat1_4_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_13291, new_AGEMA_signal_13290, mcs1_mcs_mat1_4_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, mcs1_mcs_mat1_4_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_13747, new_AGEMA_signal_13746, mcs1_mcs_mat1_4_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_14627, new_AGEMA_signal_14626, mcs1_mcs_mat1_4_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_11945, new_AGEMA_signal_11944, mcs1_mcs_mat1_4_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_15111, new_AGEMA_signal_15110, mcs1_mcs_mat1_4_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_14195, new_AGEMA_signal_14194, mcs1_mcs_mat1_4_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_14627, new_AGEMA_signal_14626, mcs1_mcs_mat1_4_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_10971, new_AGEMA_signal_10970, mcs1_mcs_mat1_4_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_13749, new_AGEMA_signal_13748, mcs1_mcs_mat1_4_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_14195, new_AGEMA_signal_14194, mcs1_mcs_mat1_4_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2417], Fresh[2416], Fresh[2415]}), .c ({new_AGEMA_signal_13749, new_AGEMA_signal_13748, mcs1_mcs_mat1_4_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({new_AGEMA_signal_11945, new_AGEMA_signal_11944, mcs1_mcs_mat1_4_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2423], Fresh[2422], Fresh[2421]}), .c ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, mcs1_mcs_mat1_4_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_10017, new_AGEMA_signal_10016, mcs1_mcs_mat1_4_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_10019, new_AGEMA_signal_10018, mcs1_mcs_mat1_4_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_10975, new_AGEMA_signal_10974, mcs1_mcs_mat1_4_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_10013, new_AGEMA_signal_10012, mcs1_mcs_mat1_4_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_7849, new_AGEMA_signal_7848, mcs1_mcs_mat1_4_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_10977, new_AGEMA_signal_10976, mcs1_mcs_mat1_4_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_9217, new_AGEMA_signal_9216, mcs1_mcs_mat1_4_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_10013, new_AGEMA_signal_10012, mcs1_mcs_mat1_4_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_10015, new_AGEMA_signal_10014, mcs1_mcs_mat1_4_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_10979, new_AGEMA_signal_10978, mcs1_mcs_mat1_4_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, mcs1_mcs_mat1_4_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_9217, new_AGEMA_signal_9216, mcs1_mcs_mat1_4_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_10015, new_AGEMA_signal_10014, mcs1_mcs_mat1_4_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_10981, new_AGEMA_signal_10980, mcs1_mcs_mat1_4_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .c ({new_AGEMA_signal_11947, new_AGEMA_signal_11946, mcs1_mcs_mat1_4_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_10017, new_AGEMA_signal_10016, mcs1_mcs_mat1_4_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, mcs1_mcs_mat1_4_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_10981, new_AGEMA_signal_10980, mcs1_mcs_mat1_4_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({new_AGEMA_signal_10019, new_AGEMA_signal_10018, mcs1_mcs_mat1_4_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2429], Fresh[2428], Fresh[2427]}), .c ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, mcs1_mcs_mat1_4_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({new_AGEMA_signal_9217, new_AGEMA_signal_9216, mcs1_mcs_mat1_4_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_14197, new_AGEMA_signal_14196, mcs1_mcs_mat1_4_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_14629, new_AGEMA_signal_14628, mcs1_mcs_mat1_4_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_13295, new_AGEMA_signal_13294, mcs1_mcs_mat1_4_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_13751, new_AGEMA_signal_13750, mcs1_mcs_mat1_4_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_14631, new_AGEMA_signal_14630, mcs1_mcs_mat1_4_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_11951, new_AGEMA_signal_11950, mcs1_mcs_mat1_4_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_15113, new_AGEMA_signal_15112, mcs1_mcs_mat1_4_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_14197, new_AGEMA_signal_14196, mcs1_mcs_mat1_4_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .c ({new_AGEMA_signal_14631, new_AGEMA_signal_14630, mcs1_mcs_mat1_4_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_10983, new_AGEMA_signal_10982, mcs1_mcs_mat1_4_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_13753, new_AGEMA_signal_13752, mcs1_mcs_mat1_4_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_14197, new_AGEMA_signal_14196, mcs1_mcs_mat1_4_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2435], Fresh[2434], Fresh[2433]}), .c ({new_AGEMA_signal_13753, new_AGEMA_signal_13752, mcs1_mcs_mat1_4_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({new_AGEMA_signal_11951, new_AGEMA_signal_11950, mcs1_mcs_mat1_4_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2441], Fresh[2440], Fresh[2439]}), .c ({new_AGEMA_signal_13295, new_AGEMA_signal_13294, mcs1_mcs_mat1_4_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_11953, new_AGEMA_signal_11952, mcs1_mcs_mat1_4_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_12713, new_AGEMA_signal_12712, mcs1_mcs_mat1_4_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_10987, new_AGEMA_signal_10986, mcs1_mcs_mat1_4_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_10023, new_AGEMA_signal_10022, mcs1_mcs_mat1_4_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_11953, new_AGEMA_signal_11952, mcs1_mcs_mat1_4_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_8791, new_AGEMA_signal_8790, mcs1_mcs_mat1_4_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_10021, new_AGEMA_signal_10020, mcs1_mcs_mat1_4_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_10023, new_AGEMA_signal_10022, mcs1_mcs_mat1_4_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_8791, new_AGEMA_signal_8790, mcs1_mcs_mat1_4_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_10985, new_AGEMA_signal_10984, mcs1_mcs_mat1_4_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_4_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_8417, new_AGEMA_signal_8416, mcs1_mcs_mat1_4_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_8791, new_AGEMA_signal_8790, mcs1_mcs_mat1_4_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_9219, new_AGEMA_signal_9218, mcs1_mcs_mat1_4_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .c ({new_AGEMA_signal_10023, new_AGEMA_signal_10022, mcs1_mcs_mat1_4_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, mcs1_mcs_mat1_4_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_4_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_12715, new_AGEMA_signal_12714, mcs1_mcs_mat1_4_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_10987, new_AGEMA_signal_10986, mcs1_mcs_mat1_4_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9219, new_AGEMA_signal_9218, mcs1_mcs_mat1_4_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, mcs1_mcs_mat1_4_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .b ({new_AGEMA_signal_10025, new_AGEMA_signal_10024, mcs1_mcs_mat1_4_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_10987, new_AGEMA_signal_10986, mcs1_mcs_mat1_4_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({new_AGEMA_signal_10025, new_AGEMA_signal_10024, mcs1_mcs_mat1_4_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2447], Fresh[2446], Fresh[2445]}), .c ({new_AGEMA_signal_8417, new_AGEMA_signal_8416, mcs1_mcs_mat1_4_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({new_AGEMA_signal_9219, new_AGEMA_signal_9218, mcs1_mcs_mat1_4_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_10989, new_AGEMA_signal_10988, mcs1_mcs_mat1_4_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_9221, new_AGEMA_signal_9220, mcs1_mcs_mat1_4_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_11957, new_AGEMA_signal_11956, mcs1_mcs_mat1_4_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_10029, new_AGEMA_signal_10028, mcs1_mcs_mat1_4_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_11959, new_AGEMA_signal_11958, mcs1_mcs_mat1_4_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12717, new_AGEMA_signal_12716, mcs1_mcs_mat1_4_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_10989, new_AGEMA_signal_10988, mcs1_mcs_mat1_4_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_11959, new_AGEMA_signal_11958, mcs1_mcs_mat1_4_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12719, new_AGEMA_signal_12718, mcs1_mcs_mat1_4_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_9221, new_AGEMA_signal_9220, mcs1_mcs_mat1_4_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_10991, new_AGEMA_signal_10990, mcs1_mcs_mat1_4_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_11959, new_AGEMA_signal_11958, mcs1_mcs_mat1_4_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, mcs1_mcs_mat1_4_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_9221, new_AGEMA_signal_9220, mcs1_mcs_mat1_4_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_10027, new_AGEMA_signal_10026, mcs1_mcs_mat1_4_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .c ({new_AGEMA_signal_10989, new_AGEMA_signal_10988, mcs1_mcs_mat1_4_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_9223, new_AGEMA_signal_9222, mcs1_mcs_mat1_4_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7853, new_AGEMA_signal_7852, mcs1_mcs_mat1_4_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_10027, new_AGEMA_signal_10026, mcs1_mcs_mat1_4_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_10991, new_AGEMA_signal_10990, mcs1_mcs_mat1_4_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_10029, new_AGEMA_signal_10028, mcs1_mcs_mat1_4_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_11961, new_AGEMA_signal_11960, mcs1_mcs_mat1_4_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_9223, new_AGEMA_signal_9222, mcs1_mcs_mat1_4_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_10029, new_AGEMA_signal_10028, mcs1_mcs_mat1_4_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({new_AGEMA_signal_10031, new_AGEMA_signal_10030, mcs1_mcs_mat1_4_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_10991, new_AGEMA_signal_10990, mcs1_mcs_mat1_4_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2453], Fresh[2452], Fresh[2451]}), .c ({new_AGEMA_signal_10031, new_AGEMA_signal_10030, mcs1_mcs_mat1_4_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, mcs1_mcs_mat1_4_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2459], Fresh[2458], Fresh[2457]}), .c ({new_AGEMA_signal_9223, new_AGEMA_signal_9222, mcs1_mcs_mat1_4_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_11965, new_AGEMA_signal_11964, mcs1_mcs_mat1_4_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_12721, new_AGEMA_signal_12720, mcs1_mcs_mat1_4_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({new_AGEMA_signal_10993, new_AGEMA_signal_10992, mcs1_mcs_mat1_4_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_11963, new_AGEMA_signal_11962, mcs1_mcs_mat1_4_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_12723, new_AGEMA_signal_12722, mcs1_mcs_mat1_4_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_9225, new_AGEMA_signal_9224, mcs1_mcs_mat1_4_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_13297, new_AGEMA_signal_13296, mcs1_mcs_mat1_4_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_11965, new_AGEMA_signal_11964, mcs1_mcs_mat1_4_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .c ({new_AGEMA_signal_12723, new_AGEMA_signal_12722, mcs1_mcs_mat1_4_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_10993, new_AGEMA_signal_10992, mcs1_mcs_mat1_4_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_11965, new_AGEMA_signal_11964, mcs1_mcs_mat1_4_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_7855, new_AGEMA_signal_7854, mcs1_mcs_mat1_4_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_10035, new_AGEMA_signal_10034, mcs1_mcs_mat1_4_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_10993, new_AGEMA_signal_10992, mcs1_mcs_mat1_4_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({new_AGEMA_signal_10035, new_AGEMA_signal_10034, mcs1_mcs_mat1_4_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2465], Fresh[2464], Fresh[2463]}), .c ({new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2468], Fresh[2467], Fresh[2466]}), .c ({new_AGEMA_signal_9225, new_AGEMA_signal_9224, mcs1_mcs_mat1_4_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_14203, new_AGEMA_signal_14202, mcs1_mcs_mat1_4_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, mcs1_mcs_mat1_4_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_14633, new_AGEMA_signal_14632, mcs1_mcs_mat1_4_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_11967, new_AGEMA_signal_11966, mcs1_mcs_mat1_4_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_13755, new_AGEMA_signal_13754, mcs1_mcs_mat1_4_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_14199, new_AGEMA_signal_14198, mcs1_mcs_mat1_4_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({new_AGEMA_signal_13757, new_AGEMA_signal_13756, mcs1_mcs_mat1_4_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_14201, new_AGEMA_signal_14200, mcs1_mcs_mat1_4_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2471], Fresh[2470], Fresh[2469]}), .c ({new_AGEMA_signal_13757, new_AGEMA_signal_13756, mcs1_mcs_mat1_4_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({new_AGEMA_signal_11967, new_AGEMA_signal_11966, mcs1_mcs_mat1_4_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2477], Fresh[2476], Fresh[2475]}), .c ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, mcs1_mcs_mat1_4_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, mcs1_mcs_mat1_4_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_9227, new_AGEMA_signal_9226, mcs1_mcs_mat1_4_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_10037, new_AGEMA_signal_10036, mcs1_mcs_mat1_4_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_4_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_10039, new_AGEMA_signal_10038, mcs1_mcs_mat1_4_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_10999, new_AGEMA_signal_10998, mcs1_mcs_mat1_4_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_11001, new_AGEMA_signal_11000, mcs1_mcs_mat1_4_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_10041, new_AGEMA_signal_10040, mcs1_mcs_mat1_4_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_11969, new_AGEMA_signal_11968, mcs1_mcs_mat1_4_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_10043, new_AGEMA_signal_10042, mcs1_mcs_mat1_4_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_11001, new_AGEMA_signal_11000, mcs1_mcs_mat1_4_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2480], Fresh[2479], Fresh[2478]}), .c ({new_AGEMA_signal_10043, new_AGEMA_signal_10042, mcs1_mcs_mat1_4_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2483], Fresh[2482], Fresh[2481]}), .c ({new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_4_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({new_AGEMA_signal_9227, new_AGEMA_signal_9226, mcs1_mcs_mat1_4_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, mcs1_mcs_mat1_4_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_11003, new_AGEMA_signal_11002, mcs1_mcs_mat1_4_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_11971, new_AGEMA_signal_11970, mcs1_mcs_mat1_4_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_11973, new_AGEMA_signal_11972, mcs1_mcs_mat1_4_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_10045, new_AGEMA_signal_10044, mcs1_mcs_mat1_4_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_12725, new_AGEMA_signal_12724, mcs1_mcs_mat1_4_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_9229, new_AGEMA_signal_9228, mcs1_mcs_mat1_4_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_10045, new_AGEMA_signal_10044, mcs1_mcs_mat1_4_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({new_AGEMA_signal_11973, new_AGEMA_signal_11972, mcs1_mcs_mat1_4_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_12727, new_AGEMA_signal_12726, mcs1_mcs_mat1_4_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_7859, new_AGEMA_signal_7858, mcs1_mcs_mat1_4_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_11003, new_AGEMA_signal_11002, mcs1_mcs_mat1_4_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_11973, new_AGEMA_signal_11972, mcs1_mcs_mat1_4_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_8429, new_AGEMA_signal_8428, mcs1_mcs_mat1_4_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_10051, new_AGEMA_signal_10050, mcs1_mcs_mat1_4_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_11003, new_AGEMA_signal_11002, mcs1_mcs_mat1_4_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_10049, new_AGEMA_signal_10048, mcs1_mcs_mat1_4_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_11005, new_AGEMA_signal_11004, mcs1_mcs_mat1_4_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_11975, new_AGEMA_signal_11974, mcs1_mcs_mat1_4_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, mcs1_mcs_mat1_4_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8429, new_AGEMA_signal_8428, mcs1_mcs_mat1_4_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_11005, new_AGEMA_signal_11004, mcs1_mcs_mat1_4_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_9229, new_AGEMA_signal_9228, mcs1_mcs_mat1_4_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, mcs1_mcs_mat1_4_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2489], Fresh[2488], Fresh[2487]}), .c ({new_AGEMA_signal_10051, new_AGEMA_signal_10050, mcs1_mcs_mat1_4_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({new_AGEMA_signal_8429, new_AGEMA_signal_8428, mcs1_mcs_mat1_4_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2495], Fresh[2494], Fresh[2493]}), .c ({new_AGEMA_signal_9229, new_AGEMA_signal_9228, mcs1_mcs_mat1_4_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_13303, new_AGEMA_signal_13302, mcs1_mcs_mat1_4_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_13759, new_AGEMA_signal_13758, mcs1_mcs_mat1_4_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_15117, new_AGEMA_signal_15116, mcs1_mcs_mat1_4_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_11977, new_AGEMA_signal_11976, mcs1_mcs_mat1_4_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_15657, new_AGEMA_signal_15656, mcs1_mcs_mat1_4_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_14637, new_AGEMA_signal_14636, mcs1_mcs_mat1_4_mcs_out[47]}), .b ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_15117, new_AGEMA_signal_15116, mcs1_mcs_mat1_4_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_14205, new_AGEMA_signal_14204, mcs1_mcs_mat1_4_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .c ({new_AGEMA_signal_14637, new_AGEMA_signal_14636, mcs1_mcs_mat1_4_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_11009, new_AGEMA_signal_11008, mcs1_mcs_mat1_4_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_13761, new_AGEMA_signal_13760, mcs1_mcs_mat1_4_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_14205, new_AGEMA_signal_14204, mcs1_mcs_mat1_4_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({new_AGEMA_signal_13761, new_AGEMA_signal_13760, mcs1_mcs_mat1_4_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2501], Fresh[2500], Fresh[2499]}), .c ({new_AGEMA_signal_11977, new_AGEMA_signal_11976, mcs1_mcs_mat1_4_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2504], Fresh[2503], Fresh[2502]}), .c ({new_AGEMA_signal_13303, new_AGEMA_signal_13302, mcs1_mcs_mat1_4_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_11011, new_AGEMA_signal_11010, mcs1_mcs_mat1_4_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_9231, new_AGEMA_signal_9230, mcs1_mcs_mat1_4_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_11979, new_AGEMA_signal_11978, mcs1_mcs_mat1_4_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_10055, new_AGEMA_signal_10054, mcs1_mcs_mat1_4_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, mcs1_mcs_mat1_4_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_11011, new_AGEMA_signal_11010, mcs1_mcs_mat1_4_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_11013, new_AGEMA_signal_11012, mcs1_mcs_mat1_4_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_10059, new_AGEMA_signal_10058, mcs1_mcs_mat1_4_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_11981, new_AGEMA_signal_11980, mcs1_mcs_mat1_4_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_11015, new_AGEMA_signal_11014, mcs1_mcs_mat1_4_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_7861, new_AGEMA_signal_7860, mcs1_mcs_mat1_4_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_11983, new_AGEMA_signal_11982, mcs1_mcs_mat1_4_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_10055, new_AGEMA_signal_10054, mcs1_mcs_mat1_4_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9233, new_AGEMA_signal_9232, mcs1_mcs_mat1_4_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_11015, new_AGEMA_signal_11014, mcs1_mcs_mat1_4_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_10057, new_AGEMA_signal_10056, mcs1_mcs_mat1_4_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_9233, new_AGEMA_signal_9232, mcs1_mcs_mat1_4_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_11017, new_AGEMA_signal_11016, mcs1_mcs_mat1_4_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2507], Fresh[2506], Fresh[2505]}), .c ({new_AGEMA_signal_10059, new_AGEMA_signal_10058, mcs1_mcs_mat1_4_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, mcs1_mcs_mat1_4_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2513], Fresh[2512], Fresh[2511]}), .c ({new_AGEMA_signal_9233, new_AGEMA_signal_9232, mcs1_mcs_mat1_4_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_11985, new_AGEMA_signal_11984, mcs1_mcs_mat1_4_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_7863, new_AGEMA_signal_7862, mcs1_mcs_mat1_4_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, mcs1_mcs_mat1_4_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_9237, new_AGEMA_signal_9236, mcs1_mcs_mat1_4_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_9235, new_AGEMA_signal_9234, mcs1_mcs_mat1_4_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_10061, new_AGEMA_signal_10060, mcs1_mcs_mat1_4_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({new_AGEMA_signal_11985, new_AGEMA_signal_11984, mcs1_mcs_mat1_4_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_12731, new_AGEMA_signal_12730, mcs1_mcs_mat1_4_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_10063, new_AGEMA_signal_10062, mcs1_mcs_mat1_4_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_11019, new_AGEMA_signal_11018, mcs1_mcs_mat1_4_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_11985, new_AGEMA_signal_11984, mcs1_mcs_mat1_4_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_10065, new_AGEMA_signal_10064, mcs1_mcs_mat1_4_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9239, new_AGEMA_signal_9238, mcs1_mcs_mat1_4_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_11019, new_AGEMA_signal_11018, mcs1_mcs_mat1_4_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_10065, new_AGEMA_signal_10064, mcs1_mcs_mat1_4_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9237, new_AGEMA_signal_9236, mcs1_mcs_mat1_4_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_11021, new_AGEMA_signal_11020, mcs1_mcs_mat1_4_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_8793, new_AGEMA_signal_8792, mcs1_mcs_mat1_4_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_9237, new_AGEMA_signal_9236, mcs1_mcs_mat1_4_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({new_AGEMA_signal_8433, new_AGEMA_signal_8432, mcs1_mcs_mat1_4_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_8793, new_AGEMA_signal_8792, mcs1_mcs_mat1_4_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2516], Fresh[2515], Fresh[2514]}), .c ({new_AGEMA_signal_10065, new_AGEMA_signal_10064, mcs1_mcs_mat1_4_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2519], Fresh[2518], Fresh[2517]}), .c ({new_AGEMA_signal_8433, new_AGEMA_signal_8432, mcs1_mcs_mat1_4_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({new_AGEMA_signal_9239, new_AGEMA_signal_9238, mcs1_mcs_mat1_4_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_10067, new_AGEMA_signal_10066, mcs1_mcs_mat1_4_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_9241, new_AGEMA_signal_9240, mcs1_mcs_mat1_4_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_11023, new_AGEMA_signal_11022, mcs1_mcs_mat1_4_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_8435, new_AGEMA_signal_8434, mcs1_mcs_mat1_4_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_8795, new_AGEMA_signal_8794, mcs1_mcs_mat1_4_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_12733, new_AGEMA_signal_12732, mcs1_mcs_mat1_4_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_10069, new_AGEMA_signal_10068, mcs1_mcs_mat1_4_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, mcs1_mcs_mat1_4_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2525], Fresh[2524], Fresh[2523]}), .c ({new_AGEMA_signal_10069, new_AGEMA_signal_10068, mcs1_mcs_mat1_4_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2528], Fresh[2527], Fresh[2526]}), .c ({new_AGEMA_signal_8435, new_AGEMA_signal_8434, mcs1_mcs_mat1_4_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2531], Fresh[2530], Fresh[2529]}), .c ({new_AGEMA_signal_9241, new_AGEMA_signal_9240, mcs1_mcs_mat1_4_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_14639, new_AGEMA_signal_14638, mcs1_mcs_mat1_4_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_14207, new_AGEMA_signal_14206, mcs1_mcs_mat1_4_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_15119, new_AGEMA_signal_15118, mcs1_mcs_mat1_4_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_11991, new_AGEMA_signal_11990, mcs1_mcs_mat1_4_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_14209, new_AGEMA_signal_14208, mcs1_mcs_mat1_4_mcs_out[29]}), .c ({new_AGEMA_signal_14639, new_AGEMA_signal_14638, mcs1_mcs_mat1_4_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_11989, new_AGEMA_signal_11988, mcs1_mcs_mat1_4_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_14207, new_AGEMA_signal_14206, mcs1_mcs_mat1_4_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_14641, new_AGEMA_signal_14640, mcs1_mcs_mat1_4_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_13767, new_AGEMA_signal_13766, mcs1_mcs_mat1_4_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .c ({new_AGEMA_signal_14207, new_AGEMA_signal_14206, mcs1_mcs_mat1_4_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_14643, new_AGEMA_signal_14642, mcs1_mcs_mat1_4_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_13763, new_AGEMA_signal_13762, mcs1_mcs_mat1_4_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_15121, new_AGEMA_signal_15120, mcs1_mcs_mat1_4_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_14211, new_AGEMA_signal_14210, mcs1_mcs_mat1_4_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_13765, new_AGEMA_signal_13764, mcs1_mcs_mat1_4_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_14643, new_AGEMA_signal_14642, mcs1_mcs_mat1_4_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_13307, new_AGEMA_signal_13306, mcs1_mcs_mat1_4_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_13765, new_AGEMA_signal_13764, mcs1_mcs_mat1_4_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_13767, new_AGEMA_signal_13766, mcs1_mcs_mat1_4_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_11991, new_AGEMA_signal_11990, mcs1_mcs_mat1_4_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_14211, new_AGEMA_signal_14210, mcs1_mcs_mat1_4_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({new_AGEMA_signal_13767, new_AGEMA_signal_13766, mcs1_mcs_mat1_4_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2537], Fresh[2536], Fresh[2535]}), .c ({new_AGEMA_signal_11991, new_AGEMA_signal_11990, mcs1_mcs_mat1_4_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2540], Fresh[2539], Fresh[2538]}), .c ({new_AGEMA_signal_13307, new_AGEMA_signal_13306, mcs1_mcs_mat1_4_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_10071, new_AGEMA_signal_10070, mcs1_mcs_mat1_4_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_11029, new_AGEMA_signal_11028, mcs1_mcs_mat1_4_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_9243, new_AGEMA_signal_9242, mcs1_mcs_mat1_4_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8437, new_AGEMA_signal_8436, mcs1_mcs_mat1_4_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_10071, new_AGEMA_signal_10070, mcs1_mcs_mat1_4_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_11031, new_AGEMA_signal_11030, mcs1_mcs_mat1_4_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_11993, new_AGEMA_signal_11992, mcs1_mcs_mat1_4_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_10075, new_AGEMA_signal_10074, mcs1_mcs_mat1_4_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8437, new_AGEMA_signal_8436, mcs1_mcs_mat1_4_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_11031, new_AGEMA_signal_11030, mcs1_mcs_mat1_4_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_11995, new_AGEMA_signal_11994, mcs1_mcs_mat1_4_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .c ({new_AGEMA_signal_12735, new_AGEMA_signal_12734, mcs1_mcs_mat1_4_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_10075, new_AGEMA_signal_10074, mcs1_mcs_mat1_4_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_11033, new_AGEMA_signal_11032, mcs1_mcs_mat1_4_mcs_out[24]}), .c ({new_AGEMA_signal_11995, new_AGEMA_signal_11994, mcs1_mcs_mat1_4_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_10073, new_AGEMA_signal_10072, mcs1_mcs_mat1_4_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .c ({new_AGEMA_signal_11033, new_AGEMA_signal_11032, mcs1_mcs_mat1_4_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_9243, new_AGEMA_signal_9242, mcs1_mcs_mat1_4_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7867, new_AGEMA_signal_7866, mcs1_mcs_mat1_4_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_10073, new_AGEMA_signal_10072, mcs1_mcs_mat1_4_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2543], Fresh[2542], Fresh[2541]}), .c ({new_AGEMA_signal_10075, new_AGEMA_signal_10074, mcs1_mcs_mat1_4_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({new_AGEMA_signal_8437, new_AGEMA_signal_8436, mcs1_mcs_mat1_4_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2549], Fresh[2548], Fresh[2547]}), .c ({new_AGEMA_signal_9243, new_AGEMA_signal_9242, mcs1_mcs_mat1_4_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_10077, new_AGEMA_signal_10076, mcs1_mcs_mat1_4_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .c ({new_AGEMA_signal_11035, new_AGEMA_signal_11034, mcs1_mcs_mat1_4_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_9245, new_AGEMA_signal_9244, mcs1_mcs_mat1_4_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8439, new_AGEMA_signal_8438, mcs1_mcs_mat1_4_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_10077, new_AGEMA_signal_10076, mcs1_mcs_mat1_4_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_11037, new_AGEMA_signal_11036, mcs1_mcs_mat1_4_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .c ({new_AGEMA_signal_11997, new_AGEMA_signal_11996, mcs1_mcs_mat1_4_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_10081, new_AGEMA_signal_10080, mcs1_mcs_mat1_4_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8439, new_AGEMA_signal_8438, mcs1_mcs_mat1_4_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_11037, new_AGEMA_signal_11036, mcs1_mcs_mat1_4_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_11999, new_AGEMA_signal_11998, mcs1_mcs_mat1_4_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_12737, new_AGEMA_signal_12736, mcs1_mcs_mat1_4_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_10081, new_AGEMA_signal_10080, mcs1_mcs_mat1_4_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_11039, new_AGEMA_signal_11038, mcs1_mcs_mat1_4_mcs_out[20]}), .c ({new_AGEMA_signal_11999, new_AGEMA_signal_11998, mcs1_mcs_mat1_4_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_10079, new_AGEMA_signal_10078, mcs1_mcs_mat1_4_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_11039, new_AGEMA_signal_11038, mcs1_mcs_mat1_4_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_9245, new_AGEMA_signal_9244, mcs1_mcs_mat1_4_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7869, new_AGEMA_signal_7868, mcs1_mcs_mat1_4_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_10079, new_AGEMA_signal_10078, mcs1_mcs_mat1_4_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({new_AGEMA_signal_10081, new_AGEMA_signal_10080, mcs1_mcs_mat1_4_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2555], Fresh[2554], Fresh[2553]}), .c ({new_AGEMA_signal_8439, new_AGEMA_signal_8438, mcs1_mcs_mat1_4_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({new_AGEMA_signal_9245, new_AGEMA_signal_9244, mcs1_mcs_mat1_4_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_10083, new_AGEMA_signal_10082, mcs1_mcs_mat1_4_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_10089, new_AGEMA_signal_10088, mcs1_mcs_mat1_4_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_11041, new_AGEMA_signal_11040, mcs1_mcs_mat1_4_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_11043, new_AGEMA_signal_11042, mcs1_mcs_mat1_4_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_7871, new_AGEMA_signal_7870, mcs1_mcs_mat1_4_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_12001, new_AGEMA_signal_12000, mcs1_mcs_mat1_4_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_12003, new_AGEMA_signal_12002, mcs1_mcs_mat1_4_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_8441, new_AGEMA_signal_8440, mcs1_mcs_mat1_4_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_12739, new_AGEMA_signal_12738, mcs1_mcs_mat1_4_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_11043, new_AGEMA_signal_11042, mcs1_mcs_mat1_4_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_12003, new_AGEMA_signal_12002, mcs1_mcs_mat1_4_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_10085, new_AGEMA_signal_10084, mcs1_mcs_mat1_4_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .c ({new_AGEMA_signal_11043, new_AGEMA_signal_11042, mcs1_mcs_mat1_4_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_9247, new_AGEMA_signal_9246, mcs1_mcs_mat1_4_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_9249, new_AGEMA_signal_9248, mcs1_mcs_mat1_4_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_10085, new_AGEMA_signal_10084, mcs1_mcs_mat1_4_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_10087, new_AGEMA_signal_10086, mcs1_mcs_mat1_4_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_8441, new_AGEMA_signal_8440, mcs1_mcs_mat1_4_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_11045, new_AGEMA_signal_11044, mcs1_mcs_mat1_4_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2561], Fresh[2560], Fresh[2559]}), .c ({new_AGEMA_signal_10089, new_AGEMA_signal_10088, mcs1_mcs_mat1_4_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2564], Fresh[2563], Fresh[2562]}), .c ({new_AGEMA_signal_8441, new_AGEMA_signal_8440, mcs1_mcs_mat1_4_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2567], Fresh[2566], Fresh[2565]}), .c ({new_AGEMA_signal_9249, new_AGEMA_signal_9248, mcs1_mcs_mat1_4_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_14649, new_AGEMA_signal_14648, mcs1_mcs_mat1_4_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_12741, new_AGEMA_signal_12740, mcs1_mcs_mat1_4_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_15123, new_AGEMA_signal_15122, mcs1_mcs_mat1_4_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_14217, new_AGEMA_signal_14216, mcs1_mcs_mat1_4_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_14213, new_AGEMA_signal_14212, mcs1_mcs_mat1_4_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_14645, new_AGEMA_signal_14644, mcs1_mcs_mat1_4_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_13771, new_AGEMA_signal_13770, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_12005, new_AGEMA_signal_12004, mcs1_mcs_mat1_4_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_14213, new_AGEMA_signal_14212, mcs1_mcs_mat1_4_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_12741, new_AGEMA_signal_12740, mcs1_mcs_mat1_4_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_14215, new_AGEMA_signal_14214, mcs1_mcs_mat1_4_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_14647, new_AGEMA_signal_14646, mcs1_mcs_mat1_4_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_13769, new_AGEMA_signal_13768, mcs1_mcs_mat1_4_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_13771, new_AGEMA_signal_13770, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_14215, new_AGEMA_signal_14214, mcs1_mcs_mat1_4_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_11047, new_AGEMA_signal_11046, mcs1_mcs_mat1_4_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_12005, new_AGEMA_signal_12004, mcs1_mcs_mat1_4_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_12741, new_AGEMA_signal_12740, mcs1_mcs_mat1_4_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_15125, new_AGEMA_signal_15124, mcs1_mcs_mat1_4_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_15659, new_AGEMA_signal_15658, mcs1_mcs_mat1_4_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_14649, new_AGEMA_signal_14648, mcs1_mcs_mat1_4_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_13771, new_AGEMA_signal_13770, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_15125, new_AGEMA_signal_15124, mcs1_mcs_mat1_4_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_14217, new_AGEMA_signal_14216, mcs1_mcs_mat1_4_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_14649, new_AGEMA_signal_14648, mcs1_mcs_mat1_4_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_13769, new_AGEMA_signal_13768, mcs1_mcs_mat1_4_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_14217, new_AGEMA_signal_14216, mcs1_mcs_mat1_4_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_9497, new_AGEMA_signal_9496, shiftr_out[108]}), .b ({new_AGEMA_signal_13309, new_AGEMA_signal_13308, mcs1_mcs_mat1_4_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_13769, new_AGEMA_signal_13768, mcs1_mcs_mat1_4_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({new_AGEMA_signal_13771, new_AGEMA_signal_13770, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10457, new_AGEMA_signal_10456, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2573], Fresh[2572], Fresh[2571]}), .c ({new_AGEMA_signal_12005, new_AGEMA_signal_12004, mcs1_mcs_mat1_4_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2576], Fresh[2575], Fresh[2574]}), .c ({new_AGEMA_signal_13309, new_AGEMA_signal_13308, mcs1_mcs_mat1_4_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_8797, new_AGEMA_signal_8796, mcs1_mcs_mat1_4_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .c ({new_AGEMA_signal_9251, new_AGEMA_signal_9250, mcs1_mcs_mat1_4_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_11051, new_AGEMA_signal_11050, mcs1_mcs_mat1_4_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_12007, new_AGEMA_signal_12006, mcs1_mcs_mat1_4_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_10091, new_AGEMA_signal_10090, mcs1_mcs_mat1_4_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_11049, new_AGEMA_signal_11048, mcs1_mcs_mat1_4_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_9253, new_AGEMA_signal_9252, mcs1_mcs_mat1_4_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_8797, new_AGEMA_signal_8796, mcs1_mcs_mat1_4_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_10091, new_AGEMA_signal_10090, mcs1_mcs_mat1_4_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_7873, new_AGEMA_signal_7872, mcs1_mcs_mat1_4_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8443, new_AGEMA_signal_8442, mcs1_mcs_mat1_4_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_8797, new_AGEMA_signal_8796, mcs1_mcs_mat1_4_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, mcs1_mcs_mat1_4_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, shiftr_out[76]}), .c ({new_AGEMA_signal_12743, new_AGEMA_signal_12742, mcs1_mcs_mat1_4_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_7873, new_AGEMA_signal_7872, mcs1_mcs_mat1_4_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_11051, new_AGEMA_signal_11050, mcs1_mcs_mat1_4_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, mcs1_mcs_mat1_4_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_10093, new_AGEMA_signal_10092, mcs1_mcs_mat1_4_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_9253, new_AGEMA_signal_9252, mcs1_mcs_mat1_4_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_11051, new_AGEMA_signal_11050, mcs1_mcs_mat1_4_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8861, new_AGEMA_signal_8860, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2579], Fresh[2578], Fresh[2577]}), .c ({new_AGEMA_signal_10093, new_AGEMA_signal_10092, mcs1_mcs_mat1_4_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7637, new_AGEMA_signal_7636, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({new_AGEMA_signal_8443, new_AGEMA_signal_8442, mcs1_mcs_mat1_4_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8729, new_AGEMA_signal_8728, shiftr_out[79]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2585], Fresh[2584], Fresh[2583]}), .c ({new_AGEMA_signal_9253, new_AGEMA_signal_9252, mcs1_mcs_mat1_4_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, mcs1_mcs_mat1_4_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_9257, new_AGEMA_signal_9256, mcs1_mcs_mat1_4_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_13773, new_AGEMA_signal_13772, mcs1_mcs_mat1_4_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_12745, new_AGEMA_signal_12744, mcs1_mcs_mat1_4_mcs_out[7]}), .b ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .c ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, mcs1_mcs_mat1_4_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_12011, new_AGEMA_signal_12010, mcs1_mcs_mat1_4_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .c ({new_AGEMA_signal_12745, new_AGEMA_signal_12744, mcs1_mcs_mat1_4_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_11053, new_AGEMA_signal_11052, mcs1_mcs_mat1_4_mcs_out[6]}), .b ({new_AGEMA_signal_8447, new_AGEMA_signal_8446, mcs1_mcs_mat1_4_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_12011, new_AGEMA_signal_12010, mcs1_mcs_mat1_4_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_8445, new_AGEMA_signal_8444, mcs1_mcs_mat1_4_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_10095, new_AGEMA_signal_10094, mcs1_mcs_mat1_4_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_11053, new_AGEMA_signal_11052, mcs1_mcs_mat1_4_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8873, new_AGEMA_signal_8872, shiftr_out[45]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2588], Fresh[2587], Fresh[2586]}), .c ({new_AGEMA_signal_10095, new_AGEMA_signal_10094, mcs1_mcs_mat1_4_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7648, shiftr_out[46]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2591], Fresh[2590], Fresh[2589]}), .c ({new_AGEMA_signal_8447, new_AGEMA_signal_8446, mcs1_mcs_mat1_4_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8741, new_AGEMA_signal_8740, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({new_AGEMA_signal_9257, new_AGEMA_signal_9256, mcs1_mcs_mat1_4_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_9259, new_AGEMA_signal_9258, mcs1_mcs_mat1_4_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_10097, new_AGEMA_signal_10096, mcs1_mcs_mat1_4_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_11057, new_AGEMA_signal_11056, mcs1_mcs_mat1_4_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .b ({new_AGEMA_signal_9261, new_AGEMA_signal_9260, mcs1_mcs_mat1_4_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_10097, new_AGEMA_signal_10096, mcs1_mcs_mat1_4_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_11059, new_AGEMA_signal_11058, mcs1_mcs_mat1_4_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_8449, new_AGEMA_signal_8448, mcs1_mcs_mat1_4_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_12013, new_AGEMA_signal_12012, mcs1_mcs_mat1_4_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_11061, new_AGEMA_signal_11060, mcs1_mcs_mat1_4_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_10101, new_AGEMA_signal_10100, mcs1_mcs_mat1_4_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_12015, new_AGEMA_signal_12014, mcs1_mcs_mat1_4_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_10103, new_AGEMA_signal_10102, mcs1_mcs_mat1_4_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_7877, new_AGEMA_signal_7876, mcs1_mcs_mat1_4_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_11061, new_AGEMA_signal_11060, mcs1_mcs_mat1_4_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8885, new_AGEMA_signal_8884, shiftr_out[13]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2597], Fresh[2596], Fresh[2595]}), .c ({new_AGEMA_signal_10103, new_AGEMA_signal_10102, mcs1_mcs_mat1_4_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7661, new_AGEMA_signal_7660, shiftr_out[14]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2600], Fresh[2599], Fresh[2598]}), .c ({new_AGEMA_signal_8449, new_AGEMA_signal_8448, mcs1_mcs_mat1_4_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8753, new_AGEMA_signal_8752, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2603], Fresh[2602], Fresh[2601]}), .c ({new_AGEMA_signal_9261, new_AGEMA_signal_9260, mcs1_mcs_mat1_4_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U96 ( .a ({new_AGEMA_signal_13313, new_AGEMA_signal_13312, mcs1_mcs_mat1_5_n128}), .b ({new_AGEMA_signal_12747, new_AGEMA_signal_12746, mcs1_mcs_mat1_5_n127}), .c ({temp_next_s2[73], temp_next_s1[73], temp_next_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U95 ( .a ({new_AGEMA_signal_12101, new_AGEMA_signal_12100, mcs1_mcs_mat1_5_mcs_out[41]}), .b ({new_AGEMA_signal_10175, new_AGEMA_signal_10174, mcs1_mcs_mat1_5_mcs_out[45]}), .c ({new_AGEMA_signal_12747, new_AGEMA_signal_12746, mcs1_mcs_mat1_5_n127}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U94 ( .a ({new_AGEMA_signal_12813, new_AGEMA_signal_12812, mcs1_mcs_mat1_5_mcs_out[33]}), .b ({new_AGEMA_signal_12811, new_AGEMA_signal_12810, mcs1_mcs_mat1_5_mcs_out[37]}), .c ({new_AGEMA_signal_13313, new_AGEMA_signal_13312, mcs1_mcs_mat1_5_n128}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U93 ( .a ({new_AGEMA_signal_16095, new_AGEMA_signal_16094, mcs1_mcs_mat1_5_n126}), .b ({new_AGEMA_signal_13777, new_AGEMA_signal_13776, mcs1_mcs_mat1_5_n125}), .c ({temp_next_s2[72], temp_next_s1[72], temp_next_s0[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U92 ( .a ({new_AGEMA_signal_11137, new_AGEMA_signal_11136, mcs1_mcs_mat1_5_mcs_out[40]}), .b ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, mcs1_mcs_mat1_5_mcs_out[44]}), .c ({new_AGEMA_signal_13777, new_AGEMA_signal_13776, mcs1_mcs_mat1_5_n125}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U91 ( .a ({new_AGEMA_signal_15687, new_AGEMA_signal_15686, mcs1_mcs_mat1_5_mcs_out[32]}), .b ({new_AGEMA_signal_11141, new_AGEMA_signal_11140, mcs1_mcs_mat1_5_mcs_out[36]}), .c ({new_AGEMA_signal_16095, new_AGEMA_signal_16094, mcs1_mcs_mat1_5_n126}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U90 ( .a ({new_AGEMA_signal_14651, new_AGEMA_signal_14650, mcs1_mcs_mat1_5_n124}), .b ({new_AGEMA_signal_13315, new_AGEMA_signal_13314, mcs1_mcs_mat1_5_n123}), .c ({temp_next_s2[43], temp_next_s1[43], temp_next_s0[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U89 ( .a ({new_AGEMA_signal_11151, new_AGEMA_signal_11150, mcs1_mcs_mat1_5_mcs_out[27]}), .b ({new_AGEMA_signal_12815, new_AGEMA_signal_12814, mcs1_mcs_mat1_5_mcs_out[31]}), .c ({new_AGEMA_signal_13315, new_AGEMA_signal_13314, mcs1_mcs_mat1_5_n123}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U88 ( .a ({new_AGEMA_signal_14253, new_AGEMA_signal_14252, mcs1_mcs_mat1_5_mcs_out[19]}), .b ({new_AGEMA_signal_11157, new_AGEMA_signal_11156, mcs1_mcs_mat1_5_mcs_out[23]}), .c ({new_AGEMA_signal_14651, new_AGEMA_signal_14650, mcs1_mcs_mat1_5_n124}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U87 ( .a ({new_AGEMA_signal_15129, new_AGEMA_signal_15128, mcs1_mcs_mat1_5_n122}), .b ({new_AGEMA_signal_12749, new_AGEMA_signal_12748, mcs1_mcs_mat1_5_n121}), .c ({temp_next_s2[42], temp_next_s1[42], temp_next_s0[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U86 ( .a ({new_AGEMA_signal_12113, new_AGEMA_signal_12112, mcs1_mcs_mat1_5_mcs_out[26]}), .b ({new_AGEMA_signal_12109, new_AGEMA_signal_12108, mcs1_mcs_mat1_5_mcs_out[30]}), .c ({new_AGEMA_signal_12749, new_AGEMA_signal_12748, mcs1_mcs_mat1_5_n121}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U85 ( .a ({new_AGEMA_signal_14693, new_AGEMA_signal_14692, mcs1_mcs_mat1_5_mcs_out[18]}), .b ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, mcs1_mcs_mat1_5_mcs_out[22]}), .c ({new_AGEMA_signal_15129, new_AGEMA_signal_15128, mcs1_mcs_mat1_5_n122}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U84 ( .a ({new_AGEMA_signal_15663, new_AGEMA_signal_15662, mcs1_mcs_mat1_5_n120}), .b ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, mcs1_mcs_mat1_5_n119}), .c ({temp_next_s2[41], temp_next_s1[41], temp_next_s0[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U83 ( .a ({new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_5_mcs_out[25]}), .b ({new_AGEMA_signal_11147, new_AGEMA_signal_11146, mcs1_mcs_mat1_5_mcs_out[29]}), .c ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, mcs1_mcs_mat1_5_n119}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U82 ( .a ({new_AGEMA_signal_15173, new_AGEMA_signal_15172, mcs1_mcs_mat1_5_mcs_out[17]}), .b ({new_AGEMA_signal_12821, new_AGEMA_signal_12820, mcs1_mcs_mat1_5_mcs_out[21]}), .c ({new_AGEMA_signal_15663, new_AGEMA_signal_15662, mcs1_mcs_mat1_5_n120}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U81 ( .a ({new_AGEMA_signal_14653, new_AGEMA_signal_14652, mcs1_mcs_mat1_5_n118}), .b ({new_AGEMA_signal_13319, new_AGEMA_signal_13318, mcs1_mcs_mat1_5_n117}), .c ({temp_next_s2[40], temp_next_s1[40], temp_next_s0[40]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U80 ( .a ({new_AGEMA_signal_11155, new_AGEMA_signal_11154, mcs1_mcs_mat1_5_mcs_out[24]}), .b ({new_AGEMA_signal_12817, new_AGEMA_signal_12816, mcs1_mcs_mat1_5_mcs_out[28]}), .c ({new_AGEMA_signal_13319, new_AGEMA_signal_13318, mcs1_mcs_mat1_5_n117}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U79 ( .a ({new_AGEMA_signal_14257, new_AGEMA_signal_14256, mcs1_mcs_mat1_5_mcs_out[16]}), .b ({new_AGEMA_signal_11161, new_AGEMA_signal_11160, mcs1_mcs_mat1_5_mcs_out[20]}), .c ({new_AGEMA_signal_14653, new_AGEMA_signal_14652, mcs1_mcs_mat1_5_n118}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U78 ( .a ({new_AGEMA_signal_13321, new_AGEMA_signal_13320, mcs1_mcs_mat1_5_n116}), .b ({new_AGEMA_signal_14655, new_AGEMA_signal_14654, mcs1_mcs_mat1_5_n115}), .c ({temp_next_s2[11], temp_next_s1[11], temp_next_s0[11]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U77 ( .a ({new_AGEMA_signal_14259, new_AGEMA_signal_14258, mcs1_mcs_mat1_5_mcs_out[3]}), .b ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, mcs1_mcs_mat1_5_mcs_out[7]}), .c ({new_AGEMA_signal_14655, new_AGEMA_signal_14654, mcs1_mcs_mat1_5_n115}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U76 ( .a ({new_AGEMA_signal_9331, new_AGEMA_signal_9330, mcs1_mcs_mat1_5_mcs_out[11]}), .b ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, mcs1_mcs_mat1_5_mcs_out[15]}), .c ({new_AGEMA_signal_13321, new_AGEMA_signal_13320, mcs1_mcs_mat1_5_n116}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U75 ( .a ({new_AGEMA_signal_15135, new_AGEMA_signal_15134, mcs1_mcs_mat1_5_n114}), .b ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, mcs1_mcs_mat1_5_n113}), .c ({new_AGEMA_signal_15665, new_AGEMA_signal_15664, mcs_out[235]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U74 ( .a ({new_AGEMA_signal_12771, new_AGEMA_signal_12770, mcs1_mcs_mat1_5_mcs_out[123]}), .b ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, mcs1_mcs_mat1_5_n113}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U73 ( .a ({new_AGEMA_signal_14679, new_AGEMA_signal_14678, mcs1_mcs_mat1_5_mcs_out[115]}), .b ({new_AGEMA_signal_12775, new_AGEMA_signal_12774, mcs1_mcs_mat1_5_mcs_out[119]}), .c ({new_AGEMA_signal_15135, new_AGEMA_signal_15134, mcs1_mcs_mat1_5_n114}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U72 ( .a ({new_AGEMA_signal_14657, new_AGEMA_signal_14656, mcs1_mcs_mat1_5_n112}), .b ({new_AGEMA_signal_11063, new_AGEMA_signal_11062, mcs1_mcs_mat1_5_n111}), .c ({new_AGEMA_signal_15137, new_AGEMA_signal_15136, mcs_out[234]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U71 ( .a ({new_AGEMA_signal_10105, new_AGEMA_signal_10104, mcs1_mcs_mat1_5_mcs_out[122]}), .b ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_11063, new_AGEMA_signal_11062, mcs1_mcs_mat1_5_n111}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U70 ( .a ({new_AGEMA_signal_14229, new_AGEMA_signal_14228, mcs1_mcs_mat1_5_mcs_out[114]}), .b ({new_AGEMA_signal_12777, new_AGEMA_signal_12776, mcs1_mcs_mat1_5_mcs_out[118]}), .c ({new_AGEMA_signal_14657, new_AGEMA_signal_14656, mcs1_mcs_mat1_5_n112}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U69 ( .a ({new_AGEMA_signal_12751, new_AGEMA_signal_12750, mcs1_mcs_mat1_5_n110}), .b ({new_AGEMA_signal_14659, new_AGEMA_signal_14658, mcs1_mcs_mat1_5_n109}), .c ({temp_next_s2[10], temp_next_s1[10], temp_next_s0[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U68 ( .a ({new_AGEMA_signal_14261, new_AGEMA_signal_14260, mcs1_mcs_mat1_5_mcs_out[2]}), .b ({new_AGEMA_signal_11175, new_AGEMA_signal_11174, mcs1_mcs_mat1_5_mcs_out[6]}), .c ({new_AGEMA_signal_14659, new_AGEMA_signal_14658, mcs1_mcs_mat1_5_n109}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U67 ( .a ({new_AGEMA_signal_12129, new_AGEMA_signal_12128, mcs1_mcs_mat1_5_mcs_out[10]}), .b ({new_AGEMA_signal_12123, new_AGEMA_signal_12122, mcs1_mcs_mat1_5_mcs_out[14]}), .c ({new_AGEMA_signal_12751, new_AGEMA_signal_12750, mcs1_mcs_mat1_5_n110}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U66 ( .a ({new_AGEMA_signal_14219, new_AGEMA_signal_14218, mcs1_mcs_mat1_5_n108}), .b ({new_AGEMA_signal_13325, new_AGEMA_signal_13324, mcs1_mcs_mat1_5_n107}), .c ({new_AGEMA_signal_14661, new_AGEMA_signal_14660, mcs_out[233]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U65 ( .a ({new_AGEMA_signal_12773, new_AGEMA_signal_12772, mcs1_mcs_mat1_5_mcs_out[121]}), .b ({new_AGEMA_signal_9263, new_AGEMA_signal_9262, mcs1_mcs_mat1_5_mcs_out[125]}), .c ({new_AGEMA_signal_13325, new_AGEMA_signal_13324, mcs1_mcs_mat1_5_n107}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U64 ( .a ({new_AGEMA_signal_13785, new_AGEMA_signal_13784, mcs1_mcs_mat1_5_mcs_out[113]}), .b ({new_AGEMA_signal_12035, new_AGEMA_signal_12034, mcs1_mcs_mat1_5_mcs_out[117]}), .c ({new_AGEMA_signal_14219, new_AGEMA_signal_14218, mcs1_mcs_mat1_5_n108}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U63 ( .a ({new_AGEMA_signal_15667, new_AGEMA_signal_15666, mcs1_mcs_mat1_5_n106}), .b ({new_AGEMA_signal_12753, new_AGEMA_signal_12752, mcs1_mcs_mat1_5_n105}), .c ({new_AGEMA_signal_16099, new_AGEMA_signal_16098, mcs_out[232]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U62 ( .a ({new_AGEMA_signal_12029, new_AGEMA_signal_12028, mcs1_mcs_mat1_5_mcs_out[120]}), .b ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_12753, new_AGEMA_signal_12752, mcs1_mcs_mat1_5_n105}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U61 ( .a ({new_AGEMA_signal_15163, new_AGEMA_signal_15162, mcs1_mcs_mat1_5_mcs_out[112]}), .b ({new_AGEMA_signal_11075, new_AGEMA_signal_11074, mcs1_mcs_mat1_5_mcs_out[116]}), .c ({new_AGEMA_signal_15667, new_AGEMA_signal_15666, mcs1_mcs_mat1_5_n106}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U60 ( .a ({new_AGEMA_signal_12755, new_AGEMA_signal_12754, mcs1_mcs_mat1_5_n104}), .b ({new_AGEMA_signal_15669, new_AGEMA_signal_15668, mcs1_mcs_mat1_5_n103}), .c ({new_AGEMA_signal_16101, new_AGEMA_signal_16100, mcs_out[203]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U59 ( .a ({new_AGEMA_signal_12779, new_AGEMA_signal_12778, mcs1_mcs_mat1_5_mcs_out[111]}), .b ({new_AGEMA_signal_15165, new_AGEMA_signal_15164, mcs1_mcs_mat1_5_mcs_out[99]}), .c ({new_AGEMA_signal_15669, new_AGEMA_signal_15668, mcs1_mcs_mat1_5_n103}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U58 ( .a ({new_AGEMA_signal_12053, new_AGEMA_signal_12052, mcs1_mcs_mat1_5_mcs_out[103]}), .b ({new_AGEMA_signal_12045, new_AGEMA_signal_12044, mcs1_mcs_mat1_5_mcs_out[107]}), .c ({new_AGEMA_signal_12755, new_AGEMA_signal_12754, mcs1_mcs_mat1_5_n104}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U57 ( .a ({new_AGEMA_signal_12757, new_AGEMA_signal_12756, mcs1_mcs_mat1_5_n102}), .b ({new_AGEMA_signal_14663, new_AGEMA_signal_14662, mcs1_mcs_mat1_5_n101}), .c ({new_AGEMA_signal_15141, new_AGEMA_signal_15140, mcs_out[202]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U56 ( .a ({new_AGEMA_signal_12781, new_AGEMA_signal_12780, mcs1_mcs_mat1_5_mcs_out[110]}), .b ({new_AGEMA_signal_14235, new_AGEMA_signal_14234, mcs1_mcs_mat1_5_mcs_out[98]}), .c ({new_AGEMA_signal_14663, new_AGEMA_signal_14662, mcs1_mcs_mat1_5_n101}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U55 ( .a ({new_AGEMA_signal_10123, new_AGEMA_signal_10122, mcs1_mcs_mat1_5_mcs_out[102]}), .b ({new_AGEMA_signal_12047, new_AGEMA_signal_12046, mcs1_mcs_mat1_5_mcs_out[106]}), .c ({new_AGEMA_signal_12757, new_AGEMA_signal_12756, mcs1_mcs_mat1_5_n102}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U54 ( .a ({new_AGEMA_signal_12759, new_AGEMA_signal_12758, mcs1_mcs_mat1_5_n100}), .b ({new_AGEMA_signal_13779, new_AGEMA_signal_13778, mcs1_mcs_mat1_5_n99}), .c ({new_AGEMA_signal_14221, new_AGEMA_signal_14220, mcs_out[201]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U53 ( .a ({new_AGEMA_signal_12783, new_AGEMA_signal_12782, mcs1_mcs_mat1_5_mcs_out[109]}), .b ({new_AGEMA_signal_13345, new_AGEMA_signal_13344, mcs1_mcs_mat1_5_mcs_out[97]}), .c ({new_AGEMA_signal_13779, new_AGEMA_signal_13778, mcs1_mcs_mat1_5_n99}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U52 ( .a ({new_AGEMA_signal_11089, new_AGEMA_signal_11088, mcs1_mcs_mat1_5_mcs_out[101]}), .b ({new_AGEMA_signal_12049, new_AGEMA_signal_12048, mcs1_mcs_mat1_5_mcs_out[105]}), .c ({new_AGEMA_signal_12759, new_AGEMA_signal_12758, mcs1_mcs_mat1_5_n100}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U51 ( .a ({new_AGEMA_signal_13327, new_AGEMA_signal_13326, mcs1_mcs_mat1_5_n98}), .b ({new_AGEMA_signal_16375, new_AGEMA_signal_16374, mcs1_mcs_mat1_5_n97}), .c ({new_AGEMA_signal_16469, new_AGEMA_signal_16468, mcs_out[200]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U50 ( .a ({new_AGEMA_signal_12785, new_AGEMA_signal_12784, mcs1_mcs_mat1_5_mcs_out[108]}), .b ({new_AGEMA_signal_16107, new_AGEMA_signal_16106, mcs1_mcs_mat1_5_mcs_out[96]}), .c ({new_AGEMA_signal_16375, new_AGEMA_signal_16374, mcs1_mcs_mat1_5_n97}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U49 ( .a ({new_AGEMA_signal_12055, new_AGEMA_signal_12054, mcs1_mcs_mat1_5_mcs_out[100]}), .b ({new_AGEMA_signal_12787, new_AGEMA_signal_12786, mcs1_mcs_mat1_5_mcs_out[104]}), .c ({new_AGEMA_signal_13327, new_AGEMA_signal_13326, mcs1_mcs_mat1_5_n98}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U48 ( .a ({new_AGEMA_signal_14665, new_AGEMA_signal_14664, mcs1_mcs_mat1_5_n96}), .b ({new_AGEMA_signal_12761, new_AGEMA_signal_12760, mcs1_mcs_mat1_5_n95}), .c ({new_AGEMA_signal_15143, new_AGEMA_signal_15142, mcs_out[171]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U47 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_12061, new_AGEMA_signal_12060, mcs1_mcs_mat1_5_mcs_out[95]}), .c ({new_AGEMA_signal_12761, new_AGEMA_signal_12760, mcs1_mcs_mat1_5_n95}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U46 ( .a ({new_AGEMA_signal_14237, new_AGEMA_signal_14236, mcs1_mcs_mat1_5_mcs_out[83]}), .b ({new_AGEMA_signal_10137, new_AGEMA_signal_10136, mcs1_mcs_mat1_5_mcs_out[87]}), .c ({new_AGEMA_signal_14665, new_AGEMA_signal_14664, mcs1_mcs_mat1_5_n96}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U45 ( .a ({new_AGEMA_signal_14667, new_AGEMA_signal_14666, mcs1_mcs_mat1_5_n94}), .b ({new_AGEMA_signal_11065, new_AGEMA_signal_11064, mcs1_mcs_mat1_5_n93}), .c ({new_AGEMA_signal_15145, new_AGEMA_signal_15144, mcs_out[170]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U43 ( .a ({new_AGEMA_signal_14239, new_AGEMA_signal_14238, mcs1_mcs_mat1_5_mcs_out[82]}), .b ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_14667, new_AGEMA_signal_14666, mcs1_mcs_mat1_5_n94}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U42 ( .a ({new_AGEMA_signal_14669, new_AGEMA_signal_14668, mcs1_mcs_mat1_5_n92}), .b ({new_AGEMA_signal_11067, new_AGEMA_signal_11066, mcs1_mcs_mat1_5_n91}), .c ({new_AGEMA_signal_15147, new_AGEMA_signal_15146, mcs_out[169]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U41 ( .a ({new_AGEMA_signal_9293, new_AGEMA_signal_9292, mcs1_mcs_mat1_5_mcs_out[89]}), .b ({new_AGEMA_signal_10133, new_AGEMA_signal_10132, mcs1_mcs_mat1_5_mcs_out[93]}), .c ({new_AGEMA_signal_11067, new_AGEMA_signal_11066, mcs1_mcs_mat1_5_n91}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U40 ( .a ({new_AGEMA_signal_14241, new_AGEMA_signal_14240, mcs1_mcs_mat1_5_mcs_out[81]}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_14669, new_AGEMA_signal_14668, mcs1_mcs_mat1_5_n92}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U39 ( .a ({new_AGEMA_signal_15149, new_AGEMA_signal_15148, mcs1_mcs_mat1_5_n90}), .b ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, mcs1_mcs_mat1_5_n89}), .c ({new_AGEMA_signal_15671, new_AGEMA_signal_15670, mcs_out[168]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U38 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_12789, new_AGEMA_signal_12788, mcs1_mcs_mat1_5_mcs_out[92]}), .c ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, mcs1_mcs_mat1_5_n89}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U37 ( .a ({new_AGEMA_signal_14685, new_AGEMA_signal_14684, mcs1_mcs_mat1_5_mcs_out[80]}), .b ({new_AGEMA_signal_11097, new_AGEMA_signal_11096, mcs1_mcs_mat1_5_mcs_out[84]}), .c ({new_AGEMA_signal_15149, new_AGEMA_signal_15148, mcs1_mcs_mat1_5_n90}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U36 ( .a ({new_AGEMA_signal_15151, new_AGEMA_signal_15150, mcs1_mcs_mat1_5_n88}), .b ({new_AGEMA_signal_12017, new_AGEMA_signal_12016, mcs1_mcs_mat1_5_n87}), .c ({temp_next_s2[9], temp_next_s1[9], temp_next_s0[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U35 ( .a ({new_AGEMA_signal_9335, new_AGEMA_signal_9334, mcs1_mcs_mat1_5_mcs_out[5]}), .b ({new_AGEMA_signal_11171, new_AGEMA_signal_11170, mcs1_mcs_mat1_5_mcs_out[9]}), .c ({new_AGEMA_signal_12017, new_AGEMA_signal_12016, mcs1_mcs_mat1_5_n87}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U34 ( .a ({new_AGEMA_signal_12125, new_AGEMA_signal_12124, mcs1_mcs_mat1_5_mcs_out[13]}), .b ({new_AGEMA_signal_14697, new_AGEMA_signal_14696, mcs1_mcs_mat1_5_mcs_out[1]}), .c ({new_AGEMA_signal_15151, new_AGEMA_signal_15150, mcs1_mcs_mat1_5_n88}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U33 ( .a ({new_AGEMA_signal_15675, new_AGEMA_signal_15674, mcs1_mcs_mat1_5_n86}), .b ({new_AGEMA_signal_12763, new_AGEMA_signal_12762, mcs1_mcs_mat1_5_n85}), .c ({new_AGEMA_signal_16103, new_AGEMA_signal_16102, mcs_out[139]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U32 ( .a ({new_AGEMA_signal_10143, new_AGEMA_signal_10142, mcs1_mcs_mat1_5_mcs_out[75]}), .b ({new_AGEMA_signal_12067, new_AGEMA_signal_12066, mcs1_mcs_mat1_5_mcs_out[79]}), .c ({new_AGEMA_signal_12763, new_AGEMA_signal_12762, mcs1_mcs_mat1_5_n85}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U31 ( .a ({new_AGEMA_signal_15167, new_AGEMA_signal_15166, mcs1_mcs_mat1_5_mcs_out[67]}), .b ({new_AGEMA_signal_12075, new_AGEMA_signal_12074, mcs1_mcs_mat1_5_mcs_out[71]}), .c ({new_AGEMA_signal_15675, new_AGEMA_signal_15674, mcs1_mcs_mat1_5_n86}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U30 ( .a ({new_AGEMA_signal_15153, new_AGEMA_signal_15152, mcs1_mcs_mat1_5_n84}), .b ({new_AGEMA_signal_13331, new_AGEMA_signal_13330, mcs1_mcs_mat1_5_n83}), .c ({new_AGEMA_signal_15677, new_AGEMA_signal_15676, mcs_out[138]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U29 ( .a ({new_AGEMA_signal_12793, new_AGEMA_signal_12792, mcs1_mcs_mat1_5_mcs_out[74]}), .b ({new_AGEMA_signal_8465, new_AGEMA_signal_8464, mcs1_mcs_mat1_5_mcs_out[78]}), .c ({new_AGEMA_signal_13331, new_AGEMA_signal_13330, mcs1_mcs_mat1_5_n83}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U28 ( .a ({new_AGEMA_signal_14687, new_AGEMA_signal_14686, mcs1_mcs_mat1_5_mcs_out[66]}), .b ({new_AGEMA_signal_12797, new_AGEMA_signal_12796, mcs1_mcs_mat1_5_mcs_out[70]}), .c ({new_AGEMA_signal_15153, new_AGEMA_signal_15152, mcs1_mcs_mat1_5_n84}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U27 ( .a ({new_AGEMA_signal_14223, new_AGEMA_signal_14222, mcs1_mcs_mat1_5_n82}), .b ({new_AGEMA_signal_12019, new_AGEMA_signal_12018, mcs1_mcs_mat1_5_n81}), .c ({new_AGEMA_signal_14671, new_AGEMA_signal_14670, mcs_out[137]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U26 ( .a ({new_AGEMA_signal_11103, new_AGEMA_signal_11102, mcs1_mcs_mat1_5_mcs_out[73]}), .b ({new_AGEMA_signal_10139, new_AGEMA_signal_10138, mcs1_mcs_mat1_5_mcs_out[77]}), .c ({new_AGEMA_signal_12019, new_AGEMA_signal_12018, mcs1_mcs_mat1_5_n81}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U25 ( .a ({new_AGEMA_signal_13801, new_AGEMA_signal_13800, mcs1_mcs_mat1_5_mcs_out[65]}), .b ({new_AGEMA_signal_12799, new_AGEMA_signal_12798, mcs1_mcs_mat1_5_mcs_out[69]}), .c ({new_AGEMA_signal_14223, new_AGEMA_signal_14222, mcs1_mcs_mat1_5_n82}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U24 ( .a ({new_AGEMA_signal_16105, new_AGEMA_signal_16104, mcs1_mcs_mat1_5_n80}), .b ({new_AGEMA_signal_13333, new_AGEMA_signal_13332, mcs1_mcs_mat1_5_n79}), .c ({new_AGEMA_signal_16377, new_AGEMA_signal_16376, mcs_out[136]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U23 ( .a ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, mcs1_mcs_mat1_5_mcs_out[72]}), .b ({new_AGEMA_signal_12791, new_AGEMA_signal_12790, mcs1_mcs_mat1_5_mcs_out[76]}), .c ({new_AGEMA_signal_13333, new_AGEMA_signal_13332, mcs1_mcs_mat1_5_n79}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U22 ( .a ({new_AGEMA_signal_15685, new_AGEMA_signal_15684, mcs1_mcs_mat1_5_mcs_out[64]}), .b ({new_AGEMA_signal_12079, new_AGEMA_signal_12078, mcs1_mcs_mat1_5_mcs_out[68]}), .c ({new_AGEMA_signal_16105, new_AGEMA_signal_16104, mcs1_mcs_mat1_5_n80}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U21 ( .a ({new_AGEMA_signal_14225, new_AGEMA_signal_14224, mcs1_mcs_mat1_5_n78}), .b ({new_AGEMA_signal_12765, new_AGEMA_signal_12764, mcs1_mcs_mat1_5_n77}), .c ({temp_next_s2[107], temp_next_s1[107], temp_next_s0[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U20 ( .a ({new_AGEMA_signal_11119, new_AGEMA_signal_11118, mcs1_mcs_mat1_5_mcs_out[59]}), .b ({new_AGEMA_signal_12083, new_AGEMA_signal_12082, mcs1_mcs_mat1_5_mcs_out[63]}), .c ({new_AGEMA_signal_12765, new_AGEMA_signal_12764, mcs1_mcs_mat1_5_n77}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U19 ( .a ({new_AGEMA_signal_13805, new_AGEMA_signal_13804, mcs1_mcs_mat1_5_mcs_out[51]}), .b ({new_AGEMA_signal_12089, new_AGEMA_signal_12088, mcs1_mcs_mat1_5_mcs_out[55]}), .c ({new_AGEMA_signal_14225, new_AGEMA_signal_14224, mcs1_mcs_mat1_5_n78}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U18 ( .a ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, mcs1_mcs_mat1_5_n76}), .b ({new_AGEMA_signal_12021, new_AGEMA_signal_12020, mcs1_mcs_mat1_5_n75}), .c ({temp_next_s2[106], temp_next_s1[106], temp_next_s0[106]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U17 ( .a ({new_AGEMA_signal_10159, new_AGEMA_signal_10158, mcs1_mcs_mat1_5_mcs_out[58]}), .b ({new_AGEMA_signal_11113, new_AGEMA_signal_11112, mcs1_mcs_mat1_5_mcs_out[62]}), .c ({new_AGEMA_signal_12021, new_AGEMA_signal_12020, mcs1_mcs_mat1_5_n75}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U16 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_12803, new_AGEMA_signal_12802, mcs1_mcs_mat1_5_mcs_out[54]}), .c ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, mcs1_mcs_mat1_5_n76}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U15 ( .a ({new_AGEMA_signal_13337, new_AGEMA_signal_13336, mcs1_mcs_mat1_5_n74}), .b ({new_AGEMA_signal_12023, new_AGEMA_signal_12022, mcs1_mcs_mat1_5_n73}), .c ({temp_next_s2[105], temp_next_s1[105], temp_next_s0[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U14 ( .a ({new_AGEMA_signal_11121, new_AGEMA_signal_11120, mcs1_mcs_mat1_5_mcs_out[57]}), .b ({new_AGEMA_signal_11115, new_AGEMA_signal_11114, mcs1_mcs_mat1_5_mcs_out[61]}), .c ({new_AGEMA_signal_12023, new_AGEMA_signal_12022, mcs1_mcs_mat1_5_n73}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U13 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_12805, new_AGEMA_signal_12804, mcs1_mcs_mat1_5_mcs_out[53]}), .c ({new_AGEMA_signal_13337, new_AGEMA_signal_13336, mcs1_mcs_mat1_5_n74}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U12 ( .a ({new_AGEMA_signal_14675, new_AGEMA_signal_14674, mcs1_mcs_mat1_5_n72}), .b ({new_AGEMA_signal_13339, new_AGEMA_signal_13338, mcs1_mcs_mat1_5_n71}), .c ({temp_next_s2[104], temp_next_s1[104], temp_next_s0[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U11 ( .a ({new_AGEMA_signal_12087, new_AGEMA_signal_12086, mcs1_mcs_mat1_5_mcs_out[56]}), .b ({new_AGEMA_signal_12801, new_AGEMA_signal_12800, mcs1_mcs_mat1_5_mcs_out[60]}), .c ({new_AGEMA_signal_13339, new_AGEMA_signal_13338, mcs1_mcs_mat1_5_n71}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U10 ( .a ({new_AGEMA_signal_14247, new_AGEMA_signal_14246, mcs1_mcs_mat1_5_mcs_out[48]}), .b ({new_AGEMA_signal_12093, new_AGEMA_signal_12092, mcs1_mcs_mat1_5_mcs_out[52]}), .c ({new_AGEMA_signal_14675, new_AGEMA_signal_14674, mcs1_mcs_mat1_5_n72}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U9 ( .a ({new_AGEMA_signal_15157, new_AGEMA_signal_15156, mcs1_mcs_mat1_5_n70}), .b ({new_AGEMA_signal_12767, new_AGEMA_signal_12766, mcs1_mcs_mat1_5_n69}), .c ({temp_next_s2[75], temp_next_s1[75], temp_next_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U8 ( .a ({new_AGEMA_signal_12097, new_AGEMA_signal_12096, mcs1_mcs_mat1_5_mcs_out[43]}), .b ({new_AGEMA_signal_12095, new_AGEMA_signal_12094, mcs1_mcs_mat1_5_mcs_out[47]}), .c ({new_AGEMA_signal_12767, new_AGEMA_signal_12766, mcs1_mcs_mat1_5_n69}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U7 ( .a ({new_AGEMA_signal_14691, new_AGEMA_signal_14690, mcs1_mcs_mat1_5_mcs_out[35]}), .b ({new_AGEMA_signal_12809, new_AGEMA_signal_12808, mcs1_mcs_mat1_5_mcs_out[39]}), .c ({new_AGEMA_signal_15157, new_AGEMA_signal_15156, mcs1_mcs_mat1_5_n70}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U6 ( .a ({new_AGEMA_signal_14677, new_AGEMA_signal_14676, mcs1_mcs_mat1_5_n68}), .b ({new_AGEMA_signal_12769, new_AGEMA_signal_12768, mcs1_mcs_mat1_5_n67}), .c ({temp_next_s2[74], temp_next_s1[74], temp_next_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U5 ( .a ({new_AGEMA_signal_12099, new_AGEMA_signal_12098, mcs1_mcs_mat1_5_mcs_out[42]}), .b ({new_AGEMA_signal_9309, new_AGEMA_signal_9308, mcs1_mcs_mat1_5_mcs_out[46]}), .c ({new_AGEMA_signal_12769, new_AGEMA_signal_12768, mcs1_mcs_mat1_5_n67}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U4 ( .a ({new_AGEMA_signal_14249, new_AGEMA_signal_14248, mcs1_mcs_mat1_5_mcs_out[34]}), .b ({new_AGEMA_signal_10185, new_AGEMA_signal_10184, mcs1_mcs_mat1_5_mcs_out[38]}), .c ({new_AGEMA_signal_14677, new_AGEMA_signal_14676, mcs1_mcs_mat1_5_n68}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U3 ( .a ({new_AGEMA_signal_15161, new_AGEMA_signal_15160, mcs1_mcs_mat1_5_n66}), .b ({new_AGEMA_signal_14227, new_AGEMA_signal_14226, mcs1_mcs_mat1_5_n65}), .c ({temp_next_s2[8], temp_next_s1[8], temp_next_s0[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U2 ( .a ({new_AGEMA_signal_13819, new_AGEMA_signal_13818, mcs1_mcs_mat1_5_mcs_out[4]}), .b ({new_AGEMA_signal_12827, new_AGEMA_signal_12826, mcs1_mcs_mat1_5_mcs_out[8]}), .c ({new_AGEMA_signal_14227, new_AGEMA_signal_14226, mcs1_mcs_mat1_5_n65}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_U1 ( .a ({new_AGEMA_signal_14699, new_AGEMA_signal_14698, mcs1_mcs_mat1_5_mcs_out[0]}), .b ({new_AGEMA_signal_13361, new_AGEMA_signal_13360, mcs1_mcs_mat1_5_mcs_out[12]}), .c ({new_AGEMA_signal_15161, new_AGEMA_signal_15160, mcs1_mcs_mat1_5_n66}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_12025, new_AGEMA_signal_12024, mcs1_mcs_mat1_5_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_12771, new_AGEMA_signal_12770, mcs1_mcs_mat1_5_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_11069, new_AGEMA_signal_11068, mcs1_mcs_mat1_5_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_7879, new_AGEMA_signal_7878, mcs1_mcs_mat1_5_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_12025, new_AGEMA_signal_12024, mcs1_mcs_mat1_5_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_8451, new_AGEMA_signal_8450, mcs1_mcs_mat1_5_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_9265, new_AGEMA_signal_9264, mcs1_mcs_mat1_5_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_10105, new_AGEMA_signal_10104, mcs1_mcs_mat1_5_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_8453, new_AGEMA_signal_8452, mcs1_mcs_mat1_5_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .c ({new_AGEMA_signal_9265, new_AGEMA_signal_9264, mcs1_mcs_mat1_5_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_12027, new_AGEMA_signal_12026, mcs1_mcs_mat1_5_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .c ({new_AGEMA_signal_12773, new_AGEMA_signal_12772, mcs1_mcs_mat1_5_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_11069, new_AGEMA_signal_11068, mcs1_mcs_mat1_5_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_12027, new_AGEMA_signal_12026, mcs1_mcs_mat1_5_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_10107, new_AGEMA_signal_10106, mcs1_mcs_mat1_5_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9267, new_AGEMA_signal_9266, mcs1_mcs_mat1_5_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_11069, new_AGEMA_signal_11068, mcs1_mcs_mat1_5_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_11071, new_AGEMA_signal_11070, mcs1_mcs_mat1_5_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_12029, new_AGEMA_signal_12028, mcs1_mcs_mat1_5_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_10107, new_AGEMA_signal_10106, mcs1_mcs_mat1_5_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_8453, new_AGEMA_signal_8452, mcs1_mcs_mat1_5_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_11071, new_AGEMA_signal_11070, mcs1_mcs_mat1_5_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({new_AGEMA_signal_10107, new_AGEMA_signal_10106, mcs1_mcs_mat1_5_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2609], Fresh[2608], Fresh[2607]}), .c ({new_AGEMA_signal_8453, new_AGEMA_signal_8452, mcs1_mcs_mat1_5_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({new_AGEMA_signal_9267, new_AGEMA_signal_9266, mcs1_mcs_mat1_5_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_12031, new_AGEMA_signal_12030, mcs1_mcs_mat1_5_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .c ({new_AGEMA_signal_12775, new_AGEMA_signal_12774, mcs1_mcs_mat1_5_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_11073, new_AGEMA_signal_11072, mcs1_mcs_mat1_5_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9273, new_AGEMA_signal_9272, mcs1_mcs_mat1_5_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_12031, new_AGEMA_signal_12030, mcs1_mcs_mat1_5_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_12033, new_AGEMA_signal_12032, mcs1_mcs_mat1_5_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_10111, new_AGEMA_signal_10110, mcs1_mcs_mat1_5_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_12777, new_AGEMA_signal_12776, mcs1_mcs_mat1_5_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_11073, new_AGEMA_signal_11072, mcs1_mcs_mat1_5_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .c ({new_AGEMA_signal_12033, new_AGEMA_signal_12032, mcs1_mcs_mat1_5_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_11073, new_AGEMA_signal_11072, mcs1_mcs_mat1_5_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10109, new_AGEMA_signal_10108, mcs1_mcs_mat1_5_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_12035, new_AGEMA_signal_12034, mcs1_mcs_mat1_5_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_10113, new_AGEMA_signal_10112, mcs1_mcs_mat1_5_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_8455, new_AGEMA_signal_8454, mcs1_mcs_mat1_5_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_11073, new_AGEMA_signal_11072, mcs1_mcs_mat1_5_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_9271, new_AGEMA_signal_9270, mcs1_mcs_mat1_5_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_10111, new_AGEMA_signal_10110, mcs1_mcs_mat1_5_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_11075, new_AGEMA_signal_11074, mcs1_mcs_mat1_5_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_7881, new_AGEMA_signal_7880, mcs1_mcs_mat1_5_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_9273, new_AGEMA_signal_9272, mcs1_mcs_mat1_5_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_10111, new_AGEMA_signal_10110, mcs1_mcs_mat1_5_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_8455, new_AGEMA_signal_8454, mcs1_mcs_mat1_5_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_9271, new_AGEMA_signal_9270, mcs1_mcs_mat1_5_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2615], Fresh[2614], Fresh[2613]}), .c ({new_AGEMA_signal_10113, new_AGEMA_signal_10112, mcs1_mcs_mat1_5_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({new_AGEMA_signal_8455, new_AGEMA_signal_8454, mcs1_mcs_mat1_5_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2621], Fresh[2620], Fresh[2619]}), .c ({new_AGEMA_signal_9273, new_AGEMA_signal_9272, mcs1_mcs_mat1_5_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_14231, new_AGEMA_signal_14230, mcs1_mcs_mat1_5_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_12037, new_AGEMA_signal_12036, mcs1_mcs_mat1_5_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_14679, new_AGEMA_signal_14678, mcs1_mcs_mat1_5_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, mcs1_mcs_mat1_5_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_13343, new_AGEMA_signal_13342, mcs1_mcs_mat1_5_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_13785, new_AGEMA_signal_13784, mcs1_mcs_mat1_5_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_14233, new_AGEMA_signal_14232, mcs1_mcs_mat1_5_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_14681, new_AGEMA_signal_14680, mcs1_mcs_mat1_5_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_15163, new_AGEMA_signal_15162, mcs1_mcs_mat1_5_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_14231, new_AGEMA_signal_14230, mcs1_mcs_mat1_5_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_14681, new_AGEMA_signal_14680, mcs1_mcs_mat1_5_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_11077, new_AGEMA_signal_11076, mcs1_mcs_mat1_5_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_13789, new_AGEMA_signal_13788, mcs1_mcs_mat1_5_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_14231, new_AGEMA_signal_14230, mcs1_mcs_mat1_5_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_12039, new_AGEMA_signal_12038, mcs1_mcs_mat1_5_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_13787, new_AGEMA_signal_13786, mcs1_mcs_mat1_5_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_14233, new_AGEMA_signal_14232, mcs1_mcs_mat1_5_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2624], Fresh[2623], Fresh[2622]}), .c ({new_AGEMA_signal_13789, new_AGEMA_signal_13788, mcs1_mcs_mat1_5_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2627], Fresh[2626], Fresh[2625]}), .c ({new_AGEMA_signal_12039, new_AGEMA_signal_12038, mcs1_mcs_mat1_5_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({new_AGEMA_signal_13343, new_AGEMA_signal_13342, mcs1_mcs_mat1_5_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({new_AGEMA_signal_12041, new_AGEMA_signal_12040, mcs1_mcs_mat1_5_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12779, new_AGEMA_signal_12778, mcs1_mcs_mat1_5_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({new_AGEMA_signal_12043, new_AGEMA_signal_12042, mcs1_mcs_mat1_5_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12781, new_AGEMA_signal_12780, mcs1_mcs_mat1_5_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_9275, new_AGEMA_signal_9274, mcs1_mcs_mat1_5_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_12041, new_AGEMA_signal_12040, mcs1_mcs_mat1_5_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12783, new_AGEMA_signal_12782, mcs1_mcs_mat1_5_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_8457, new_AGEMA_signal_8456, mcs1_mcs_mat1_5_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_11079, new_AGEMA_signal_11078, mcs1_mcs_mat1_5_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_12041, new_AGEMA_signal_12040, mcs1_mcs_mat1_5_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_10115, new_AGEMA_signal_10114, mcs1_mcs_mat1_5_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_12043, new_AGEMA_signal_12042, mcs1_mcs_mat1_5_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12785, new_AGEMA_signal_12784, mcs1_mcs_mat1_5_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_11081, new_AGEMA_signal_11080, mcs1_mcs_mat1_5_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_12043, new_AGEMA_signal_12042, mcs1_mcs_mat1_5_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_9275, new_AGEMA_signal_9274, mcs1_mcs_mat1_5_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_10117, new_AGEMA_signal_10116, mcs1_mcs_mat1_5_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_11081, new_AGEMA_signal_11080, mcs1_mcs_mat1_5_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2633], Fresh[2632], Fresh[2631]}), .c ({new_AGEMA_signal_10117, new_AGEMA_signal_10116, mcs1_mcs_mat1_5_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2636], Fresh[2635], Fresh[2634]}), .c ({new_AGEMA_signal_8457, new_AGEMA_signal_8456, mcs1_mcs_mat1_5_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2639], Fresh[2638], Fresh[2637]}), .c ({new_AGEMA_signal_9275, new_AGEMA_signal_9274, mcs1_mcs_mat1_5_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_11085, new_AGEMA_signal_11084, mcs1_mcs_mat1_5_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_11083, new_AGEMA_signal_11082, mcs1_mcs_mat1_5_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_12045, new_AGEMA_signal_12044, mcs1_mcs_mat1_5_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_11083, new_AGEMA_signal_11082, mcs1_mcs_mat1_5_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_9277, new_AGEMA_signal_9276, mcs1_mcs_mat1_5_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_12047, new_AGEMA_signal_12046, mcs1_mcs_mat1_5_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_8459, new_AGEMA_signal_8458, mcs1_mcs_mat1_5_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .c ({new_AGEMA_signal_9277, new_AGEMA_signal_9276, mcs1_mcs_mat1_5_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_11083, new_AGEMA_signal_11082, mcs1_mcs_mat1_5_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_12049, new_AGEMA_signal_12048, mcs1_mcs_mat1_5_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_10121, new_AGEMA_signal_10120, mcs1_mcs_mat1_5_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_7885, new_AGEMA_signal_7884, mcs1_mcs_mat1_5_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_11083, new_AGEMA_signal_11082, mcs1_mcs_mat1_5_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_12051, new_AGEMA_signal_12050, mcs1_mcs_mat1_5_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_12787, new_AGEMA_signal_12786, mcs1_mcs_mat1_5_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_11085, new_AGEMA_signal_11084, mcs1_mcs_mat1_5_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_10121, new_AGEMA_signal_10120, mcs1_mcs_mat1_5_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_12051, new_AGEMA_signal_12050, mcs1_mcs_mat1_5_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_10119, new_AGEMA_signal_10118, mcs1_mcs_mat1_5_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .c ({new_AGEMA_signal_11085, new_AGEMA_signal_11084, mcs1_mcs_mat1_5_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_8459, new_AGEMA_signal_8458, mcs1_mcs_mat1_5_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_9279, new_AGEMA_signal_9278, mcs1_mcs_mat1_5_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_10119, new_AGEMA_signal_10118, mcs1_mcs_mat1_5_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({new_AGEMA_signal_10121, new_AGEMA_signal_10120, mcs1_mcs_mat1_5_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2645], Fresh[2644], Fresh[2643]}), .c ({new_AGEMA_signal_8459, new_AGEMA_signal_8458, mcs1_mcs_mat1_5_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2648], Fresh[2647], Fresh[2646]}), .c ({new_AGEMA_signal_9279, new_AGEMA_signal_9278, mcs1_mcs_mat1_5_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_9281, new_AGEMA_signal_9280, mcs1_mcs_mat1_5_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_11087, new_AGEMA_signal_11086, mcs1_mcs_mat1_5_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_12053, new_AGEMA_signal_12052, mcs1_mcs_mat1_5_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_10129, new_AGEMA_signal_10128, mcs1_mcs_mat1_5_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_11087, new_AGEMA_signal_11086, mcs1_mcs_mat1_5_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_10125, new_AGEMA_signal_10124, mcs1_mcs_mat1_5_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_9283, new_AGEMA_signal_9282, mcs1_mcs_mat1_5_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_11089, new_AGEMA_signal_11088, mcs1_mcs_mat1_5_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_10127, new_AGEMA_signal_10126, mcs1_mcs_mat1_5_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_11091, new_AGEMA_signal_11090, mcs1_mcs_mat1_5_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_12055, new_AGEMA_signal_12054, mcs1_mcs_mat1_5_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_7887, new_AGEMA_signal_7886, mcs1_mcs_mat1_5_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_10129, new_AGEMA_signal_10128, mcs1_mcs_mat1_5_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_11091, new_AGEMA_signal_11090, mcs1_mcs_mat1_5_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_8461, new_AGEMA_signal_8460, mcs1_mcs_mat1_5_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .c ({new_AGEMA_signal_10127, new_AGEMA_signal_10126, mcs1_mcs_mat1_5_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2651], Fresh[2650], Fresh[2649]}), .c ({new_AGEMA_signal_10129, new_AGEMA_signal_10128, mcs1_mcs_mat1_5_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2654], Fresh[2653], Fresh[2652]}), .c ({new_AGEMA_signal_8461, new_AGEMA_signal_8460, mcs1_mcs_mat1_5_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2657], Fresh[2656], Fresh[2655]}), .c ({new_AGEMA_signal_9283, new_AGEMA_signal_9282, mcs1_mcs_mat1_5_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_15683, new_AGEMA_signal_15682, mcs1_mcs_mat1_5_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, mcs1_mcs_mat1_5_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_16107, new_AGEMA_signal_16106, mcs1_mcs_mat1_5_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_15165, new_AGEMA_signal_15164, mcs1_mcs_mat1_5_mcs_out[99]}), .b ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .c ({new_AGEMA_signal_15683, new_AGEMA_signal_15682, mcs1_mcs_mat1_5_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_14683, new_AGEMA_signal_14682, mcs1_mcs_mat1_5_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .c ({new_AGEMA_signal_15165, new_AGEMA_signal_15164, mcs1_mcs_mat1_5_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_14235, new_AGEMA_signal_14234, mcs1_mcs_mat1_5_mcs_out[98]}), .b ({new_AGEMA_signal_12059, new_AGEMA_signal_12058, mcs1_mcs_mat1_5_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_14683, new_AGEMA_signal_14682, mcs1_mcs_mat1_5_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_12057, new_AGEMA_signal_12056, mcs1_mcs_mat1_5_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_13791, new_AGEMA_signal_13790, mcs1_mcs_mat1_5_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_14235, new_AGEMA_signal_14234, mcs1_mcs_mat1_5_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2660], Fresh[2659], Fresh[2658]}), .c ({new_AGEMA_signal_13791, new_AGEMA_signal_13790, mcs1_mcs_mat1_5_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2663], Fresh[2662], Fresh[2661]}), .c ({new_AGEMA_signal_12059, new_AGEMA_signal_12058, mcs1_mcs_mat1_5_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2666], Fresh[2665], Fresh[2664]}), .c ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, mcs1_mcs_mat1_5_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_11095, new_AGEMA_signal_11094, mcs1_mcs_mat1_5_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_12061, new_AGEMA_signal_12060, mcs1_mcs_mat1_5_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_9287, new_AGEMA_signal_9286, mcs1_mcs_mat1_5_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_9289, new_AGEMA_signal_9288, mcs1_mcs_mat1_5_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_10133, new_AGEMA_signal_10132, mcs1_mcs_mat1_5_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, mcs1_mcs_mat1_5_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_8463, new_AGEMA_signal_8462, mcs1_mcs_mat1_5_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_12789, new_AGEMA_signal_12788, mcs1_mcs_mat1_5_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_11095, new_AGEMA_signal_11094, mcs1_mcs_mat1_5_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, mcs1_mcs_mat1_5_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_7889, new_AGEMA_signal_7888, mcs1_mcs_mat1_5_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_10135, new_AGEMA_signal_10134, mcs1_mcs_mat1_5_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_11095, new_AGEMA_signal_11094, mcs1_mcs_mat1_5_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2669], Fresh[2668], Fresh[2667]}), .c ({new_AGEMA_signal_10135, new_AGEMA_signal_10134, mcs1_mcs_mat1_5_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({new_AGEMA_signal_8463, new_AGEMA_signal_8462, mcs1_mcs_mat1_5_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2675], Fresh[2674], Fresh[2673]}), .c ({new_AGEMA_signal_9289, new_AGEMA_signal_9288, mcs1_mcs_mat1_5_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_13797, new_AGEMA_signal_13796, mcs1_mcs_mat1_5_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_13799, new_AGEMA_signal_13798, mcs1_mcs_mat1_5_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_14237, new_AGEMA_signal_14236, mcs1_mcs_mat1_5_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_13793, new_AGEMA_signal_13792, mcs1_mcs_mat1_5_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_11099, new_AGEMA_signal_11098, mcs1_mcs_mat1_5_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_14239, new_AGEMA_signal_14238, mcs1_mcs_mat1_5_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_13349, new_AGEMA_signal_13348, mcs1_mcs_mat1_5_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_13793, new_AGEMA_signal_13792, mcs1_mcs_mat1_5_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_13795, new_AGEMA_signal_13794, mcs1_mcs_mat1_5_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_14241, new_AGEMA_signal_14240, mcs1_mcs_mat1_5_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_12065, new_AGEMA_signal_12064, mcs1_mcs_mat1_5_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_13349, new_AGEMA_signal_13348, mcs1_mcs_mat1_5_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_13795, new_AGEMA_signal_13794, mcs1_mcs_mat1_5_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_14243, new_AGEMA_signal_14242, mcs1_mcs_mat1_5_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .c ({new_AGEMA_signal_14685, new_AGEMA_signal_14684, mcs1_mcs_mat1_5_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_13797, new_AGEMA_signal_13796, mcs1_mcs_mat1_5_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_12065, new_AGEMA_signal_12064, mcs1_mcs_mat1_5_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_14243, new_AGEMA_signal_14242, mcs1_mcs_mat1_5_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2678], Fresh[2677], Fresh[2676]}), .c ({new_AGEMA_signal_13799, new_AGEMA_signal_13798, mcs1_mcs_mat1_5_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2681], Fresh[2680], Fresh[2679]}), .c ({new_AGEMA_signal_12065, new_AGEMA_signal_12064, mcs1_mcs_mat1_5_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2684], Fresh[2683], Fresh[2682]}), .c ({new_AGEMA_signal_13349, new_AGEMA_signal_13348, mcs1_mcs_mat1_5_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_11101, new_AGEMA_signal_11100, mcs1_mcs_mat1_5_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_12067, new_AGEMA_signal_12066, mcs1_mcs_mat1_5_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_9295, new_AGEMA_signal_9294, mcs1_mcs_mat1_5_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_10139, new_AGEMA_signal_10138, mcs1_mcs_mat1_5_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_12069, new_AGEMA_signal_12068, mcs1_mcs_mat1_5_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_8467, new_AGEMA_signal_8466, mcs1_mcs_mat1_5_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_12791, new_AGEMA_signal_12790, mcs1_mcs_mat1_5_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_11101, new_AGEMA_signal_11100, mcs1_mcs_mat1_5_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .c ({new_AGEMA_signal_12069, new_AGEMA_signal_12068, mcs1_mcs_mat1_5_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_7891, new_AGEMA_signal_7890, mcs1_mcs_mat1_5_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_10141, new_AGEMA_signal_10140, mcs1_mcs_mat1_5_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_11101, new_AGEMA_signal_11100, mcs1_mcs_mat1_5_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2687], Fresh[2686], Fresh[2685]}), .c ({new_AGEMA_signal_10141, new_AGEMA_signal_10140, mcs1_mcs_mat1_5_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2690], Fresh[2689], Fresh[2688]}), .c ({new_AGEMA_signal_8467, new_AGEMA_signal_8466, mcs1_mcs_mat1_5_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2693], Fresh[2692], Fresh[2691]}), .c ({new_AGEMA_signal_9295, new_AGEMA_signal_9294, mcs1_mcs_mat1_5_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_12071, new_AGEMA_signal_12070, mcs1_mcs_mat1_5_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_12793, new_AGEMA_signal_12792, mcs1_mcs_mat1_5_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_11105, new_AGEMA_signal_11104, mcs1_mcs_mat1_5_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_10145, new_AGEMA_signal_10144, mcs1_mcs_mat1_5_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_12071, new_AGEMA_signal_12070, mcs1_mcs_mat1_5_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, mcs1_mcs_mat1_5_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_10143, new_AGEMA_signal_10142, mcs1_mcs_mat1_5_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_10145, new_AGEMA_signal_10144, mcs1_mcs_mat1_5_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, mcs1_mcs_mat1_5_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_11103, new_AGEMA_signal_11102, mcs1_mcs_mat1_5_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, mcs1_mcs_mat1_5_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_8471, new_AGEMA_signal_8470, mcs1_mcs_mat1_5_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, mcs1_mcs_mat1_5_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_9297, new_AGEMA_signal_9296, mcs1_mcs_mat1_5_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .c ({new_AGEMA_signal_10145, new_AGEMA_signal_10144, mcs1_mcs_mat1_5_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_12073, new_AGEMA_signal_12072, mcs1_mcs_mat1_5_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, mcs1_mcs_mat1_5_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, mcs1_mcs_mat1_5_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_11105, new_AGEMA_signal_11104, mcs1_mcs_mat1_5_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9297, new_AGEMA_signal_9296, mcs1_mcs_mat1_5_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_12073, new_AGEMA_signal_12072, mcs1_mcs_mat1_5_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .b ({new_AGEMA_signal_10147, new_AGEMA_signal_10146, mcs1_mcs_mat1_5_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_11105, new_AGEMA_signal_11104, mcs1_mcs_mat1_5_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2696], Fresh[2695], Fresh[2694]}), .c ({new_AGEMA_signal_10147, new_AGEMA_signal_10146, mcs1_mcs_mat1_5_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2699], Fresh[2698], Fresh[2697]}), .c ({new_AGEMA_signal_8471, new_AGEMA_signal_8470, mcs1_mcs_mat1_5_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({new_AGEMA_signal_9297, new_AGEMA_signal_9296, mcs1_mcs_mat1_5_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_11107, new_AGEMA_signal_11106, mcs1_mcs_mat1_5_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_9299, new_AGEMA_signal_9298, mcs1_mcs_mat1_5_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_12075, new_AGEMA_signal_12074, mcs1_mcs_mat1_5_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_10151, new_AGEMA_signal_10150, mcs1_mcs_mat1_5_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_12077, new_AGEMA_signal_12076, mcs1_mcs_mat1_5_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12797, new_AGEMA_signal_12796, mcs1_mcs_mat1_5_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_11107, new_AGEMA_signal_11106, mcs1_mcs_mat1_5_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_12077, new_AGEMA_signal_12076, mcs1_mcs_mat1_5_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12799, new_AGEMA_signal_12798, mcs1_mcs_mat1_5_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_9299, new_AGEMA_signal_9298, mcs1_mcs_mat1_5_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_11109, new_AGEMA_signal_11108, mcs1_mcs_mat1_5_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_12077, new_AGEMA_signal_12076, mcs1_mcs_mat1_5_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({new_AGEMA_signal_8473, new_AGEMA_signal_8472, mcs1_mcs_mat1_5_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_9299, new_AGEMA_signal_9298, mcs1_mcs_mat1_5_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_10149, new_AGEMA_signal_10148, mcs1_mcs_mat1_5_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .c ({new_AGEMA_signal_11107, new_AGEMA_signal_11106, mcs1_mcs_mat1_5_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_9301, new_AGEMA_signal_9300, mcs1_mcs_mat1_5_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7895, new_AGEMA_signal_7894, mcs1_mcs_mat1_5_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_10149, new_AGEMA_signal_10148, mcs1_mcs_mat1_5_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_11109, new_AGEMA_signal_11108, mcs1_mcs_mat1_5_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_10151, new_AGEMA_signal_10150, mcs1_mcs_mat1_5_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_12079, new_AGEMA_signal_12078, mcs1_mcs_mat1_5_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_9301, new_AGEMA_signal_9300, mcs1_mcs_mat1_5_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_10151, new_AGEMA_signal_10150, mcs1_mcs_mat1_5_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({new_AGEMA_signal_10153, new_AGEMA_signal_10152, mcs1_mcs_mat1_5_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_11109, new_AGEMA_signal_11108, mcs1_mcs_mat1_5_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2705], Fresh[2704], Fresh[2703]}), .c ({new_AGEMA_signal_10153, new_AGEMA_signal_10152, mcs1_mcs_mat1_5_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2708], Fresh[2707], Fresh[2706]}), .c ({new_AGEMA_signal_8473, new_AGEMA_signal_8472, mcs1_mcs_mat1_5_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2711], Fresh[2710], Fresh[2709]}), .c ({new_AGEMA_signal_9301, new_AGEMA_signal_9300, mcs1_mcs_mat1_5_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_14689, new_AGEMA_signal_14688, mcs1_mcs_mat1_5_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_15167, new_AGEMA_signal_15166, mcs1_mcs_mat1_5_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({new_AGEMA_signal_14245, new_AGEMA_signal_14244, mcs1_mcs_mat1_5_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_14687, new_AGEMA_signal_14686, mcs1_mcs_mat1_5_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_15169, new_AGEMA_signal_15168, mcs1_mcs_mat1_5_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_13351, new_AGEMA_signal_13350, mcs1_mcs_mat1_5_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_15685, new_AGEMA_signal_15684, mcs1_mcs_mat1_5_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_14689, new_AGEMA_signal_14688, mcs1_mcs_mat1_5_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .c ({new_AGEMA_signal_15169, new_AGEMA_signal_15168, mcs1_mcs_mat1_5_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_12081, new_AGEMA_signal_12080, mcs1_mcs_mat1_5_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_14245, new_AGEMA_signal_14244, mcs1_mcs_mat1_5_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_14689, new_AGEMA_signal_14688, mcs1_mcs_mat1_5_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_11111, new_AGEMA_signal_11110, mcs1_mcs_mat1_5_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_13803, new_AGEMA_signal_13802, mcs1_mcs_mat1_5_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_14245, new_AGEMA_signal_14244, mcs1_mcs_mat1_5_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2714], Fresh[2713], Fresh[2712]}), .c ({new_AGEMA_signal_13803, new_AGEMA_signal_13802, mcs1_mcs_mat1_5_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2717], Fresh[2716], Fresh[2715]}), .c ({new_AGEMA_signal_12081, new_AGEMA_signal_12080, mcs1_mcs_mat1_5_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2720], Fresh[2719], Fresh[2718]}), .c ({new_AGEMA_signal_13351, new_AGEMA_signal_13350, mcs1_mcs_mat1_5_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_11117, new_AGEMA_signal_11116, mcs1_mcs_mat1_5_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_9303, new_AGEMA_signal_9302, mcs1_mcs_mat1_5_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_12083, new_AGEMA_signal_12082, mcs1_mcs_mat1_5_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_8475, new_AGEMA_signal_8474, mcs1_mcs_mat1_5_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, mcs1_mcs_mat1_5_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_11113, new_AGEMA_signal_11112, mcs1_mcs_mat1_5_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({new_AGEMA_signal_10157, new_AGEMA_signal_10156, mcs1_mcs_mat1_5_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_11115, new_AGEMA_signal_11114, mcs1_mcs_mat1_5_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2723], Fresh[2722], Fresh[2721]}), .c ({new_AGEMA_signal_10157, new_AGEMA_signal_10156, mcs1_mcs_mat1_5_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2726], Fresh[2725], Fresh[2724]}), .c ({new_AGEMA_signal_8475, new_AGEMA_signal_8474, mcs1_mcs_mat1_5_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2729], Fresh[2728], Fresh[2727]}), .c ({new_AGEMA_signal_9303, new_AGEMA_signal_9302, mcs1_mcs_mat1_5_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_8479, new_AGEMA_signal_8478, mcs1_mcs_mat1_5_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_9305, new_AGEMA_signal_9304, mcs1_mcs_mat1_5_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_10159, new_AGEMA_signal_10158, mcs1_mcs_mat1_5_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_8481, new_AGEMA_signal_8480, mcs1_mcs_mat1_5_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_10161, new_AGEMA_signal_10160, mcs1_mcs_mat1_5_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_11121, new_AGEMA_signal_11120, mcs1_mcs_mat1_5_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_11123, new_AGEMA_signal_11122, mcs1_mcs_mat1_5_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_10163, new_AGEMA_signal_10162, mcs1_mcs_mat1_5_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_12087, new_AGEMA_signal_12086, mcs1_mcs_mat1_5_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_10165, new_AGEMA_signal_10164, mcs1_mcs_mat1_5_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_11123, new_AGEMA_signal_11122, mcs1_mcs_mat1_5_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({new_AGEMA_signal_10165, new_AGEMA_signal_10164, mcs1_mcs_mat1_5_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2735], Fresh[2734], Fresh[2733]}), .c ({new_AGEMA_signal_8481, new_AGEMA_signal_8480, mcs1_mcs_mat1_5_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2738], Fresh[2737], Fresh[2736]}), .c ({new_AGEMA_signal_9305, new_AGEMA_signal_9304, mcs1_mcs_mat1_5_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_10169, new_AGEMA_signal_10168, mcs1_mcs_mat1_5_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_11125, new_AGEMA_signal_11124, mcs1_mcs_mat1_5_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_12089, new_AGEMA_signal_12088, mcs1_mcs_mat1_5_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_12091, new_AGEMA_signal_12090, mcs1_mcs_mat1_5_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_10167, new_AGEMA_signal_10166, mcs1_mcs_mat1_5_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_12803, new_AGEMA_signal_12802, mcs1_mcs_mat1_5_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_9307, new_AGEMA_signal_9306, mcs1_mcs_mat1_5_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_10167, new_AGEMA_signal_10166, mcs1_mcs_mat1_5_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({new_AGEMA_signal_12091, new_AGEMA_signal_12090, mcs1_mcs_mat1_5_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_12805, new_AGEMA_signal_12804, mcs1_mcs_mat1_5_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_7901, new_AGEMA_signal_7900, mcs1_mcs_mat1_5_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_11125, new_AGEMA_signal_11124, mcs1_mcs_mat1_5_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_12091, new_AGEMA_signal_12090, mcs1_mcs_mat1_5_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_8483, new_AGEMA_signal_8482, mcs1_mcs_mat1_5_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_10173, new_AGEMA_signal_10172, mcs1_mcs_mat1_5_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_11125, new_AGEMA_signal_11124, mcs1_mcs_mat1_5_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_10171, new_AGEMA_signal_10170, mcs1_mcs_mat1_5_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_11127, new_AGEMA_signal_11126, mcs1_mcs_mat1_5_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_12093, new_AGEMA_signal_12092, mcs1_mcs_mat1_5_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_10169, new_AGEMA_signal_10168, mcs1_mcs_mat1_5_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8483, new_AGEMA_signal_8482, mcs1_mcs_mat1_5_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_11127, new_AGEMA_signal_11126, mcs1_mcs_mat1_5_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_9307, new_AGEMA_signal_9306, mcs1_mcs_mat1_5_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_10169, new_AGEMA_signal_10168, mcs1_mcs_mat1_5_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2741], Fresh[2740], Fresh[2739]}), .c ({new_AGEMA_signal_10173, new_AGEMA_signal_10172, mcs1_mcs_mat1_5_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2744], Fresh[2743], Fresh[2742]}), .c ({new_AGEMA_signal_8483, new_AGEMA_signal_8482, mcs1_mcs_mat1_5_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2747], Fresh[2746], Fresh[2745]}), .c ({new_AGEMA_signal_9307, new_AGEMA_signal_9306, mcs1_mcs_mat1_5_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_9311, new_AGEMA_signal_9310, mcs1_mcs_mat1_5_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_10175, new_AGEMA_signal_10174, mcs1_mcs_mat1_5_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_12807, new_AGEMA_signal_12806, mcs1_mcs_mat1_5_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_8485, new_AGEMA_signal_8484, mcs1_mcs_mat1_5_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, mcs1_mcs_mat1_5_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_12095, new_AGEMA_signal_12094, mcs1_mcs_mat1_5_mcs_out[47]}), .b ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_12807, new_AGEMA_signal_12806, mcs1_mcs_mat1_5_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_11129, new_AGEMA_signal_11128, mcs1_mcs_mat1_5_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .c ({new_AGEMA_signal_12095, new_AGEMA_signal_12094, mcs1_mcs_mat1_5_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_7903, new_AGEMA_signal_7902, mcs1_mcs_mat1_5_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_10177, new_AGEMA_signal_10176, mcs1_mcs_mat1_5_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_11129, new_AGEMA_signal_11128, mcs1_mcs_mat1_5_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2750], Fresh[2749], Fresh[2748]}), .c ({new_AGEMA_signal_10177, new_AGEMA_signal_10176, mcs1_mcs_mat1_5_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2753], Fresh[2752], Fresh[2751]}), .c ({new_AGEMA_signal_8485, new_AGEMA_signal_8484, mcs1_mcs_mat1_5_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2756], Fresh[2755], Fresh[2754]}), .c ({new_AGEMA_signal_9311, new_AGEMA_signal_9310, mcs1_mcs_mat1_5_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_11131, new_AGEMA_signal_11130, mcs1_mcs_mat1_5_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_9313, new_AGEMA_signal_9312, mcs1_mcs_mat1_5_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_12097, new_AGEMA_signal_12096, mcs1_mcs_mat1_5_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_10179, new_AGEMA_signal_10178, mcs1_mcs_mat1_5_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8487, new_AGEMA_signal_8486, mcs1_mcs_mat1_5_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_11131, new_AGEMA_signal_11130, mcs1_mcs_mat1_5_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_11133, new_AGEMA_signal_11132, mcs1_mcs_mat1_5_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_10183, new_AGEMA_signal_10182, mcs1_mcs_mat1_5_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_12099, new_AGEMA_signal_12098, mcs1_mcs_mat1_5_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_11135, new_AGEMA_signal_11134, mcs1_mcs_mat1_5_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_7905, new_AGEMA_signal_7904, mcs1_mcs_mat1_5_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_12101, new_AGEMA_signal_12100, mcs1_mcs_mat1_5_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_10179, new_AGEMA_signal_10178, mcs1_mcs_mat1_5_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9315, new_AGEMA_signal_9314, mcs1_mcs_mat1_5_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_11135, new_AGEMA_signal_11134, mcs1_mcs_mat1_5_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_10181, new_AGEMA_signal_10180, mcs1_mcs_mat1_5_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_9315, new_AGEMA_signal_9314, mcs1_mcs_mat1_5_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_11137, new_AGEMA_signal_11136, mcs1_mcs_mat1_5_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2759], Fresh[2758], Fresh[2757]}), .c ({new_AGEMA_signal_10183, new_AGEMA_signal_10182, mcs1_mcs_mat1_5_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({new_AGEMA_signal_8487, new_AGEMA_signal_8486, mcs1_mcs_mat1_5_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2765], Fresh[2764], Fresh[2763]}), .c ({new_AGEMA_signal_9315, new_AGEMA_signal_9314, mcs1_mcs_mat1_5_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_12103, new_AGEMA_signal_12102, mcs1_mcs_mat1_5_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_7907, new_AGEMA_signal_7906, mcs1_mcs_mat1_5_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_12809, new_AGEMA_signal_12808, mcs1_mcs_mat1_5_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_9319, new_AGEMA_signal_9318, mcs1_mcs_mat1_5_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_9317, new_AGEMA_signal_9316, mcs1_mcs_mat1_5_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_10185, new_AGEMA_signal_10184, mcs1_mcs_mat1_5_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({new_AGEMA_signal_12103, new_AGEMA_signal_12102, mcs1_mcs_mat1_5_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_12811, new_AGEMA_signal_12810, mcs1_mcs_mat1_5_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_10187, new_AGEMA_signal_10186, mcs1_mcs_mat1_5_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_11139, new_AGEMA_signal_11138, mcs1_mcs_mat1_5_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_12103, new_AGEMA_signal_12102, mcs1_mcs_mat1_5_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_10189, new_AGEMA_signal_10188, mcs1_mcs_mat1_5_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9321, new_AGEMA_signal_9320, mcs1_mcs_mat1_5_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_11139, new_AGEMA_signal_11138, mcs1_mcs_mat1_5_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_10189, new_AGEMA_signal_10188, mcs1_mcs_mat1_5_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9319, new_AGEMA_signal_9318, mcs1_mcs_mat1_5_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_11141, new_AGEMA_signal_11140, mcs1_mcs_mat1_5_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_8801, new_AGEMA_signal_8800, mcs1_mcs_mat1_5_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_9319, new_AGEMA_signal_9318, mcs1_mcs_mat1_5_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({new_AGEMA_signal_8489, new_AGEMA_signal_8488, mcs1_mcs_mat1_5_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_8801, new_AGEMA_signal_8800, mcs1_mcs_mat1_5_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2768], Fresh[2767], Fresh[2766]}), .c ({new_AGEMA_signal_10189, new_AGEMA_signal_10188, mcs1_mcs_mat1_5_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2771], Fresh[2770], Fresh[2769]}), .c ({new_AGEMA_signal_8489, new_AGEMA_signal_8488, mcs1_mcs_mat1_5_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2774], Fresh[2773], Fresh[2772]}), .c ({new_AGEMA_signal_9321, new_AGEMA_signal_9320, mcs1_mcs_mat1_5_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_13807, new_AGEMA_signal_13806, mcs1_mcs_mat1_5_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_13355, new_AGEMA_signal_13354, mcs1_mcs_mat1_5_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_14249, new_AGEMA_signal_14248, mcs1_mcs_mat1_5_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_12105, new_AGEMA_signal_12104, mcs1_mcs_mat1_5_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_12813, new_AGEMA_signal_12812, mcs1_mcs_mat1_5_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_15171, new_AGEMA_signal_15170, mcs1_mcs_mat1_5_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_13809, new_AGEMA_signal_13808, mcs1_mcs_mat1_5_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_15687, new_AGEMA_signal_15686, mcs1_mcs_mat1_5_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2777], Fresh[2776], Fresh[2775]}), .c ({new_AGEMA_signal_13809, new_AGEMA_signal_13808, mcs1_mcs_mat1_5_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2780], Fresh[2779], Fresh[2778]}), .c ({new_AGEMA_signal_12105, new_AGEMA_signal_12104, mcs1_mcs_mat1_5_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2783], Fresh[2782], Fresh[2781]}), .c ({new_AGEMA_signal_13355, new_AGEMA_signal_13354, mcs1_mcs_mat1_5_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_12107, new_AGEMA_signal_12106, mcs1_mcs_mat1_5_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_11145, new_AGEMA_signal_11144, mcs1_mcs_mat1_5_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_12815, new_AGEMA_signal_12814, mcs1_mcs_mat1_5_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, mcs1_mcs_mat1_5_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_11147, new_AGEMA_signal_11146, mcs1_mcs_mat1_5_mcs_out[29]}), .c ({new_AGEMA_signal_12107, new_AGEMA_signal_12106, mcs1_mcs_mat1_5_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_8491, new_AGEMA_signal_8490, mcs1_mcs_mat1_5_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_11145, new_AGEMA_signal_11144, mcs1_mcs_mat1_5_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_12109, new_AGEMA_signal_12108, mcs1_mcs_mat1_5_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_10195, new_AGEMA_signal_10194, mcs1_mcs_mat1_5_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .c ({new_AGEMA_signal_11145, new_AGEMA_signal_11144, mcs1_mcs_mat1_5_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_12111, new_AGEMA_signal_12110, mcs1_mcs_mat1_5_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, mcs1_mcs_mat1_5_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_12817, new_AGEMA_signal_12816, mcs1_mcs_mat1_5_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_11149, new_AGEMA_signal_11148, mcs1_mcs_mat1_5_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_10193, new_AGEMA_signal_10192, mcs1_mcs_mat1_5_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_12111, new_AGEMA_signal_12110, mcs1_mcs_mat1_5_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_9323, new_AGEMA_signal_9322, mcs1_mcs_mat1_5_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_10193, new_AGEMA_signal_10192, mcs1_mcs_mat1_5_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_10195, new_AGEMA_signal_10194, mcs1_mcs_mat1_5_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, mcs1_mcs_mat1_5_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_11149, new_AGEMA_signal_11148, mcs1_mcs_mat1_5_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2786], Fresh[2785], Fresh[2784]}), .c ({new_AGEMA_signal_10195, new_AGEMA_signal_10194, mcs1_mcs_mat1_5_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2789], Fresh[2788], Fresh[2787]}), .c ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, mcs1_mcs_mat1_5_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({new_AGEMA_signal_9323, new_AGEMA_signal_9322, mcs1_mcs_mat1_5_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_10197, new_AGEMA_signal_10196, mcs1_mcs_mat1_5_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_11151, new_AGEMA_signal_11150, mcs1_mcs_mat1_5_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_9325, new_AGEMA_signal_9324, mcs1_mcs_mat1_5_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8495, new_AGEMA_signal_8494, mcs1_mcs_mat1_5_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_10197, new_AGEMA_signal_10196, mcs1_mcs_mat1_5_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_11153, new_AGEMA_signal_11152, mcs1_mcs_mat1_5_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_12113, new_AGEMA_signal_12112, mcs1_mcs_mat1_5_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_10201, new_AGEMA_signal_10200, mcs1_mcs_mat1_5_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8495, new_AGEMA_signal_8494, mcs1_mcs_mat1_5_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_11153, new_AGEMA_signal_11152, mcs1_mcs_mat1_5_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_12115, new_AGEMA_signal_12114, mcs1_mcs_mat1_5_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .c ({new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_5_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_10201, new_AGEMA_signal_10200, mcs1_mcs_mat1_5_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_11155, new_AGEMA_signal_11154, mcs1_mcs_mat1_5_mcs_out[24]}), .c ({new_AGEMA_signal_12115, new_AGEMA_signal_12114, mcs1_mcs_mat1_5_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_10199, new_AGEMA_signal_10198, mcs1_mcs_mat1_5_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .c ({new_AGEMA_signal_11155, new_AGEMA_signal_11154, mcs1_mcs_mat1_5_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_9325, new_AGEMA_signal_9324, mcs1_mcs_mat1_5_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7911, new_AGEMA_signal_7910, mcs1_mcs_mat1_5_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_10199, new_AGEMA_signal_10198, mcs1_mcs_mat1_5_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2795], Fresh[2794], Fresh[2793]}), .c ({new_AGEMA_signal_10201, new_AGEMA_signal_10200, mcs1_mcs_mat1_5_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2798], Fresh[2797], Fresh[2796]}), .c ({new_AGEMA_signal_8495, new_AGEMA_signal_8494, mcs1_mcs_mat1_5_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2801], Fresh[2800], Fresh[2799]}), .c ({new_AGEMA_signal_9325, new_AGEMA_signal_9324, mcs1_mcs_mat1_5_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_5_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .c ({new_AGEMA_signal_11157, new_AGEMA_signal_11156, mcs1_mcs_mat1_5_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_9327, new_AGEMA_signal_9326, mcs1_mcs_mat1_5_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8497, new_AGEMA_signal_8496, mcs1_mcs_mat1_5_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_5_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_11159, new_AGEMA_signal_11158, mcs1_mcs_mat1_5_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .c ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, mcs1_mcs_mat1_5_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, mcs1_mcs_mat1_5_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8497, new_AGEMA_signal_8496, mcs1_mcs_mat1_5_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_11159, new_AGEMA_signal_11158, mcs1_mcs_mat1_5_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_12119, new_AGEMA_signal_12118, mcs1_mcs_mat1_5_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_7511, new_AGEMA_signal_7510, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_12821, new_AGEMA_signal_12820, mcs1_mcs_mat1_5_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, mcs1_mcs_mat1_5_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_11161, new_AGEMA_signal_11160, mcs1_mcs_mat1_5_mcs_out[20]}), .c ({new_AGEMA_signal_12119, new_AGEMA_signal_12118, mcs1_mcs_mat1_5_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_10205, new_AGEMA_signal_10204, mcs1_mcs_mat1_5_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_11161, new_AGEMA_signal_11160, mcs1_mcs_mat1_5_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_9327, new_AGEMA_signal_9326, mcs1_mcs_mat1_5_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7913, new_AGEMA_signal_7912, mcs1_mcs_mat1_5_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_10205, new_AGEMA_signal_10204, mcs1_mcs_mat1_5_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2804], Fresh[2803], Fresh[2802]}), .c ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, mcs1_mcs_mat1_5_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2807], Fresh[2806], Fresh[2805]}), .c ({new_AGEMA_signal_8497, new_AGEMA_signal_8496, mcs1_mcs_mat1_5_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2810], Fresh[2809], Fresh[2808]}), .c ({new_AGEMA_signal_9327, new_AGEMA_signal_9326, mcs1_mcs_mat1_5_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_13811, new_AGEMA_signal_13810, mcs1_mcs_mat1_5_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_13817, new_AGEMA_signal_13816, mcs1_mcs_mat1_5_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_14253, new_AGEMA_signal_14252, mcs1_mcs_mat1_5_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_14255, new_AGEMA_signal_14254, mcs1_mcs_mat1_5_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_11163, new_AGEMA_signal_11162, mcs1_mcs_mat1_5_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_14693, new_AGEMA_signal_14692, mcs1_mcs_mat1_5_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_14695, new_AGEMA_signal_14694, mcs1_mcs_mat1_5_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_12121, new_AGEMA_signal_12120, mcs1_mcs_mat1_5_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_15173, new_AGEMA_signal_15172, mcs1_mcs_mat1_5_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_9509, new_AGEMA_signal_9508, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_14255, new_AGEMA_signal_14254, mcs1_mcs_mat1_5_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_14695, new_AGEMA_signal_14694, mcs1_mcs_mat1_5_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_13813, new_AGEMA_signal_13812, mcs1_mcs_mat1_5_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .c ({new_AGEMA_signal_14255, new_AGEMA_signal_14254, mcs1_mcs_mat1_5_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_13357, new_AGEMA_signal_13356, mcs1_mcs_mat1_5_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, mcs1_mcs_mat1_5_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_13813, new_AGEMA_signal_13812, mcs1_mcs_mat1_5_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_13815, new_AGEMA_signal_13814, mcs1_mcs_mat1_5_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_12121, new_AGEMA_signal_12120, mcs1_mcs_mat1_5_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_14257, new_AGEMA_signal_14256, mcs1_mcs_mat1_5_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2813], Fresh[2812], Fresh[2811]}), .c ({new_AGEMA_signal_13817, new_AGEMA_signal_13816, mcs1_mcs_mat1_5_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2816], Fresh[2815], Fresh[2814]}), .c ({new_AGEMA_signal_12121, new_AGEMA_signal_12120, mcs1_mcs_mat1_5_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2819], Fresh[2818], Fresh[2817]}), .c ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, mcs1_mcs_mat1_5_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_12127, new_AGEMA_signal_12126, mcs1_mcs_mat1_5_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_8803, new_AGEMA_signal_8802, mcs1_mcs_mat1_5_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, mcs1_mcs_mat1_5_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_11169, new_AGEMA_signal_11168, mcs1_mcs_mat1_5_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_11165, new_AGEMA_signal_11164, mcs1_mcs_mat1_5_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_12123, new_AGEMA_signal_12122, mcs1_mcs_mat1_5_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_10211, new_AGEMA_signal_10210, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_8499, new_AGEMA_signal_8498, mcs1_mcs_mat1_5_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_11165, new_AGEMA_signal_11164, mcs1_mcs_mat1_5_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_8803, new_AGEMA_signal_8802, mcs1_mcs_mat1_5_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_11167, new_AGEMA_signal_11166, mcs1_mcs_mat1_5_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_12125, new_AGEMA_signal_12124, mcs1_mcs_mat1_5_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_10211, new_AGEMA_signal_10210, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_11167, new_AGEMA_signal_11166, mcs1_mcs_mat1_5_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_7915, new_AGEMA_signal_7914, mcs1_mcs_mat1_5_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_8499, new_AGEMA_signal_8498, mcs1_mcs_mat1_5_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8803, new_AGEMA_signal_8802, mcs1_mcs_mat1_5_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_5_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_13361, new_AGEMA_signal_13360, mcs1_mcs_mat1_5_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_12127, new_AGEMA_signal_12126, mcs1_mcs_mat1_5_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_10211, new_AGEMA_signal_10210, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_5_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_11169, new_AGEMA_signal_11168, mcs1_mcs_mat1_5_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_12127, new_AGEMA_signal_12126, mcs1_mcs_mat1_5_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_11169, new_AGEMA_signal_11168, mcs1_mcs_mat1_5_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, shiftr_out[104]}), .b ({new_AGEMA_signal_9329, new_AGEMA_signal_9328, mcs1_mcs_mat1_5_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8849, new_AGEMA_signal_8848, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({new_AGEMA_signal_10211, new_AGEMA_signal_10210, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7624, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2825], Fresh[2824], Fresh[2823]}), .c ({new_AGEMA_signal_8499, new_AGEMA_signal_8498, mcs1_mcs_mat1_5_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8717, new_AGEMA_signal_8716, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2828], Fresh[2827], Fresh[2826]}), .c ({new_AGEMA_signal_9329, new_AGEMA_signal_9328, mcs1_mcs_mat1_5_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_8805, new_AGEMA_signal_8804, mcs1_mcs_mat1_5_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .c ({new_AGEMA_signal_9331, new_AGEMA_signal_9330, mcs1_mcs_mat1_5_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_11173, new_AGEMA_signal_11172, mcs1_mcs_mat1_5_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_12129, new_AGEMA_signal_12128, mcs1_mcs_mat1_5_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, mcs1_mcs_mat1_5_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_11171, new_AGEMA_signal_11170, mcs1_mcs_mat1_5_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_9333, new_AGEMA_signal_9332, mcs1_mcs_mat1_5_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_8805, new_AGEMA_signal_8804, mcs1_mcs_mat1_5_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, mcs1_mcs_mat1_5_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_7917, new_AGEMA_signal_7916, mcs1_mcs_mat1_5_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8501, new_AGEMA_signal_8500, mcs1_mcs_mat1_5_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_8805, new_AGEMA_signal_8804, mcs1_mcs_mat1_5_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_12131, new_AGEMA_signal_12130, mcs1_mcs_mat1_5_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_7499, new_AGEMA_signal_7498, shiftr_out[72]}), .c ({new_AGEMA_signal_12827, new_AGEMA_signal_12826, mcs1_mcs_mat1_5_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_7917, new_AGEMA_signal_7916, mcs1_mcs_mat1_5_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_11173, new_AGEMA_signal_11172, mcs1_mcs_mat1_5_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_12131, new_AGEMA_signal_12130, mcs1_mcs_mat1_5_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_5_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_9333, new_AGEMA_signal_9332, mcs1_mcs_mat1_5_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_11173, new_AGEMA_signal_11172, mcs1_mcs_mat1_5_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2831], Fresh[2830], Fresh[2829]}), .c ({new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_5_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2834], Fresh[2833], Fresh[2832]}), .c ({new_AGEMA_signal_8501, new_AGEMA_signal_8500, mcs1_mcs_mat1_5_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, shiftr_out[75]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2837], Fresh[2836], Fresh[2835]}), .c ({new_AGEMA_signal_9333, new_AGEMA_signal_9332, mcs1_mcs_mat1_5_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_13363, new_AGEMA_signal_13362, mcs1_mcs_mat1_5_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_9337, new_AGEMA_signal_9336, mcs1_mcs_mat1_5_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_13819, new_AGEMA_signal_13818, mcs1_mcs_mat1_5_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, mcs1_mcs_mat1_5_mcs_out[7]}), .b ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .c ({new_AGEMA_signal_13363, new_AGEMA_signal_13362, mcs1_mcs_mat1_5_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_12133, new_AGEMA_signal_12132, mcs1_mcs_mat1_5_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .c ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, mcs1_mcs_mat1_5_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_11175, new_AGEMA_signal_11174, mcs1_mcs_mat1_5_mcs_out[6]}), .b ({new_AGEMA_signal_8505, new_AGEMA_signal_8504, mcs1_mcs_mat1_5_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_12133, new_AGEMA_signal_12132, mcs1_mcs_mat1_5_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_8503, new_AGEMA_signal_8502, mcs1_mcs_mat1_5_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_10217, new_AGEMA_signal_10216, mcs1_mcs_mat1_5_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_11175, new_AGEMA_signal_11174, mcs1_mcs_mat1_5_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, shiftr_out[41]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2840], Fresh[2839], Fresh[2838]}), .c ({new_AGEMA_signal_10217, new_AGEMA_signal_10216, mcs1_mcs_mat1_5_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, shiftr_out[42]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2843], Fresh[2842], Fresh[2841]}), .c ({new_AGEMA_signal_8505, new_AGEMA_signal_8504, mcs1_mcs_mat1_5_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2846], Fresh[2845], Fresh[2844]}), .c ({new_AGEMA_signal_9337, new_AGEMA_signal_9336, mcs1_mcs_mat1_5_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, mcs1_mcs_mat1_5_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_13821, new_AGEMA_signal_13820, mcs1_mcs_mat1_5_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_14261, new_AGEMA_signal_14260, mcs1_mcs_mat1_5_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .b ({new_AGEMA_signal_13367, new_AGEMA_signal_13366, mcs1_mcs_mat1_5_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_13821, new_AGEMA_signal_13820, mcs1_mcs_mat1_5_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_14263, new_AGEMA_signal_14262, mcs1_mcs_mat1_5_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_12135, new_AGEMA_signal_12134, mcs1_mcs_mat1_5_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_14697, new_AGEMA_signal_14696, mcs1_mcs_mat1_5_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_14265, new_AGEMA_signal_14264, mcs1_mcs_mat1_5_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_13825, new_AGEMA_signal_13824, mcs1_mcs_mat1_5_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_14699, new_AGEMA_signal_14698, mcs1_mcs_mat1_5_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_13827, new_AGEMA_signal_13826, mcs1_mcs_mat1_5_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_11177, new_AGEMA_signal_11176, mcs1_mcs_mat1_5_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_14265, new_AGEMA_signal_14264, mcs1_mcs_mat1_5_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, shiftr_out[9]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2849], Fresh[2848], Fresh[2847]}), .c ({new_AGEMA_signal_13827, new_AGEMA_signal_13826, mcs1_mcs_mat1_5_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10469, new_AGEMA_signal_10468, shiftr_out[10]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({new_AGEMA_signal_12135, new_AGEMA_signal_12134, mcs1_mcs_mat1_5_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2855], Fresh[2854], Fresh[2853]}), .c ({new_AGEMA_signal_13367, new_AGEMA_signal_13366, mcs1_mcs_mat1_5_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U96 ( .a ({new_AGEMA_signal_15689, new_AGEMA_signal_15688, mcs1_mcs_mat1_6_n128}), .b ({new_AGEMA_signal_12831, new_AGEMA_signal_12830, mcs1_mcs_mat1_6_n127}), .c ({temp_next_s2[69], temp_next_s1[69], temp_next_s0[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U95 ( .a ({new_AGEMA_signal_12207, new_AGEMA_signal_12206, mcs1_mcs_mat1_6_mcs_out[41]}), .b ({new_AGEMA_signal_10281, new_AGEMA_signal_10280, mcs1_mcs_mat1_6_mcs_out[45]}), .c ({new_AGEMA_signal_12831, new_AGEMA_signal_12830, mcs1_mcs_mat1_6_n127}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U94 ( .a ({new_AGEMA_signal_8809, new_AGEMA_signal_8808, mcs1_mcs_mat1_6_mcs_out[33]}), .b ({new_AGEMA_signal_15219, new_AGEMA_signal_15218, mcs1_mcs_mat1_6_mcs_out[37]}), .c ({new_AGEMA_signal_15689, new_AGEMA_signal_15688, mcs1_mcs_mat1_6_n128}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U93 ( .a ({new_AGEMA_signal_14701, new_AGEMA_signal_14700, mcs1_mcs_mat1_6_n126}), .b ({new_AGEMA_signal_13829, new_AGEMA_signal_13828, mcs1_mcs_mat1_6_n125}), .c ({temp_next_s2[68], temp_next_s1[68], temp_next_s0[68]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U92 ( .a ({new_AGEMA_signal_11253, new_AGEMA_signal_11252, mcs1_mcs_mat1_6_mcs_out[40]}), .b ({new_AGEMA_signal_13417, new_AGEMA_signal_13416, mcs1_mcs_mat1_6_mcs_out[44]}), .c ({new_AGEMA_signal_13829, new_AGEMA_signal_13828, mcs1_mcs_mat1_6_n125}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U91 ( .a ({new_AGEMA_signal_13425, new_AGEMA_signal_13424, mcs1_mcs_mat1_6_mcs_out[32]}), .b ({new_AGEMA_signal_14299, new_AGEMA_signal_14298, mcs1_mcs_mat1_6_mcs_out[36]}), .c ({new_AGEMA_signal_14701, new_AGEMA_signal_14700, mcs1_mcs_mat1_6_n126}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U90 ( .a ({new_AGEMA_signal_14703, new_AGEMA_signal_14702, mcs1_mcs_mat1_6_n124}), .b ({new_AGEMA_signal_13369, new_AGEMA_signal_13368, mcs1_mcs_mat1_6_n123}), .c ({temp_next_s2[39], temp_next_s1[39], temp_next_s0[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U89 ( .a ({new_AGEMA_signal_11267, new_AGEMA_signal_11266, mcs1_mcs_mat1_6_mcs_out[27]}), .b ({new_AGEMA_signal_12891, new_AGEMA_signal_12890, mcs1_mcs_mat1_6_mcs_out[31]}), .c ({new_AGEMA_signal_13369, new_AGEMA_signal_13368, mcs1_mcs_mat1_6_n123}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U88 ( .a ({new_AGEMA_signal_11275, new_AGEMA_signal_11274, mcs1_mcs_mat1_6_mcs_out[19]}), .b ({new_AGEMA_signal_14301, new_AGEMA_signal_14300, mcs1_mcs_mat1_6_mcs_out[23]}), .c ({new_AGEMA_signal_14703, new_AGEMA_signal_14702, mcs1_mcs_mat1_6_n124}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U87 ( .a ({new_AGEMA_signal_15179, new_AGEMA_signal_15178, mcs1_mcs_mat1_6_n122}), .b ({new_AGEMA_signal_12833, new_AGEMA_signal_12832, mcs1_mcs_mat1_6_n121}), .c ({temp_next_s2[38], temp_next_s1[38], temp_next_s0[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U86 ( .a ({new_AGEMA_signal_12219, new_AGEMA_signal_12218, mcs1_mcs_mat1_6_mcs_out[26]}), .b ({new_AGEMA_signal_12215, new_AGEMA_signal_12214, mcs1_mcs_mat1_6_mcs_out[30]}), .c ({new_AGEMA_signal_12833, new_AGEMA_signal_12832, mcs1_mcs_mat1_6_n121}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U85 ( .a ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, mcs1_mcs_mat1_6_mcs_out[18]}), .b ({new_AGEMA_signal_14745, new_AGEMA_signal_14744, mcs1_mcs_mat1_6_mcs_out[22]}), .c ({new_AGEMA_signal_15179, new_AGEMA_signal_15178, mcs1_mcs_mat1_6_n122}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U84 ( .a ({new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_6_n120}), .b ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, mcs1_mcs_mat1_6_n119}), .c ({temp_next_s2[37], temp_next_s1[37], temp_next_s0[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U83 ( .a ({new_AGEMA_signal_12895, new_AGEMA_signal_12894, mcs1_mcs_mat1_6_mcs_out[25]}), .b ({new_AGEMA_signal_11263, new_AGEMA_signal_11262, mcs1_mcs_mat1_6_mcs_out[29]}), .c ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, mcs1_mcs_mat1_6_n119}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U82 ( .a ({new_AGEMA_signal_12897, new_AGEMA_signal_12896, mcs1_mcs_mat1_6_mcs_out[17]}), .b ({new_AGEMA_signal_15221, new_AGEMA_signal_15220, mcs1_mcs_mat1_6_mcs_out[21]}), .c ({new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_6_n120}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U81 ( .a ({new_AGEMA_signal_14705, new_AGEMA_signal_14704, mcs1_mcs_mat1_6_n118}), .b ({new_AGEMA_signal_13373, new_AGEMA_signal_13372, mcs1_mcs_mat1_6_n117}), .c ({temp_next_s2[36], temp_next_s1[36], temp_next_s0[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U80 ( .a ({new_AGEMA_signal_11271, new_AGEMA_signal_11270, mcs1_mcs_mat1_6_mcs_out[24]}), .b ({new_AGEMA_signal_12893, new_AGEMA_signal_12892, mcs1_mcs_mat1_6_mcs_out[28]}), .c ({new_AGEMA_signal_13373, new_AGEMA_signal_13372, mcs1_mcs_mat1_6_n117}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U79 ( .a ({new_AGEMA_signal_11279, new_AGEMA_signal_11278, mcs1_mcs_mat1_6_mcs_out[16]}), .b ({new_AGEMA_signal_14305, new_AGEMA_signal_14304, mcs1_mcs_mat1_6_mcs_out[20]}), .c ({new_AGEMA_signal_14705, new_AGEMA_signal_14704, mcs1_mcs_mat1_6_n118}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U78 ( .a ({new_AGEMA_signal_13375, new_AGEMA_signal_13374, mcs1_mcs_mat1_6_n116}), .b ({new_AGEMA_signal_15695, new_AGEMA_signal_15694, mcs1_mcs_mat1_6_n115}), .c ({temp_next_s2[7], temp_next_s1[7], temp_next_s0[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U77 ( .a ({new_AGEMA_signal_11293, new_AGEMA_signal_11292, mcs1_mcs_mat1_6_mcs_out[3]}), .b ({new_AGEMA_signal_15223, new_AGEMA_signal_15222, mcs1_mcs_mat1_6_mcs_out[7]}), .c ({new_AGEMA_signal_15695, new_AGEMA_signal_15694, mcs1_mcs_mat1_6_n115}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U76 ( .a ({new_AGEMA_signal_9401, new_AGEMA_signal_9400, mcs1_mcs_mat1_6_mcs_out[11]}), .b ({new_AGEMA_signal_12899, new_AGEMA_signal_12898, mcs1_mcs_mat1_6_mcs_out[15]}), .c ({new_AGEMA_signal_13375, new_AGEMA_signal_13374, mcs1_mcs_mat1_6_n116}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U75 ( .a ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, mcs1_mcs_mat1_6_n114}), .b ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, mcs1_mcs_mat1_6_n113}), .c ({new_AGEMA_signal_16115, new_AGEMA_signal_16114, mcs_out[231]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U74 ( .a ({new_AGEMA_signal_12853, new_AGEMA_signal_12852, mcs1_mcs_mat1_6_mcs_out[123]}), .b ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, mcs1_mcs_mat1_6_n113}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U73 ( .a ({new_AGEMA_signal_12153, new_AGEMA_signal_12152, mcs1_mcs_mat1_6_mcs_out[115]}), .b ({new_AGEMA_signal_15205, new_AGEMA_signal_15204, mcs1_mcs_mat1_6_mcs_out[119]}), .c ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, mcs1_mcs_mat1_6_n114}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U72 ( .a ({new_AGEMA_signal_15699, new_AGEMA_signal_15698, mcs1_mcs_mat1_6_n112}), .b ({new_AGEMA_signal_11179, new_AGEMA_signal_11178, mcs1_mcs_mat1_6_n111}), .c ({new_AGEMA_signal_16117, new_AGEMA_signal_16116, mcs_out[230]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U71 ( .a ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, mcs1_mcs_mat1_6_mcs_out[122]}), .b ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_11179, new_AGEMA_signal_11178, mcs1_mcs_mat1_6_n111}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U70 ( .a ({new_AGEMA_signal_11191, new_AGEMA_signal_11190, mcs1_mcs_mat1_6_mcs_out[114]}), .b ({new_AGEMA_signal_15207, new_AGEMA_signal_15206, mcs1_mcs_mat1_6_mcs_out[118]}), .c ({new_AGEMA_signal_15699, new_AGEMA_signal_15698, mcs1_mcs_mat1_6_n112}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U69 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, mcs1_mcs_mat1_6_n110}), .b ({new_AGEMA_signal_14707, new_AGEMA_signal_14706, mcs1_mcs_mat1_6_n109}), .c ({temp_next_s2[6], temp_next_s1[6], temp_next_s0[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U68 ( .a ({new_AGEMA_signal_11295, new_AGEMA_signal_11294, mcs1_mcs_mat1_6_mcs_out[2]}), .b ({new_AGEMA_signal_14307, new_AGEMA_signal_14306, mcs1_mcs_mat1_6_mcs_out[6]}), .c ({new_AGEMA_signal_14707, new_AGEMA_signal_14706, mcs1_mcs_mat1_6_n109}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U67 ( .a ({new_AGEMA_signal_12235, new_AGEMA_signal_12234, mcs1_mcs_mat1_6_mcs_out[10]}), .b ({new_AGEMA_signal_12229, new_AGEMA_signal_12228, mcs1_mcs_mat1_6_mcs_out[14]}), .c ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, mcs1_mcs_mat1_6_n110}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U66 ( .a ({new_AGEMA_signal_15185, new_AGEMA_signal_15184, mcs1_mcs_mat1_6_n108}), .b ({new_AGEMA_signal_13379, new_AGEMA_signal_13378, mcs1_mcs_mat1_6_n107}), .c ({new_AGEMA_signal_15701, new_AGEMA_signal_15700, mcs_out[229]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U65 ( .a ({new_AGEMA_signal_12855, new_AGEMA_signal_12854, mcs1_mcs_mat1_6_mcs_out[121]}), .b ({new_AGEMA_signal_9339, new_AGEMA_signal_9338, mcs1_mcs_mat1_6_mcs_out[125]}), .c ({new_AGEMA_signal_13379, new_AGEMA_signal_13378, mcs1_mcs_mat1_6_n107}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U64 ( .a ({new_AGEMA_signal_10223, new_AGEMA_signal_10222, mcs1_mcs_mat1_6_mcs_out[113]}), .b ({new_AGEMA_signal_14725, new_AGEMA_signal_14724, mcs1_mcs_mat1_6_mcs_out[117]}), .c ({new_AGEMA_signal_15185, new_AGEMA_signal_15184, mcs1_mcs_mat1_6_n108}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U63 ( .a ({new_AGEMA_signal_14709, new_AGEMA_signal_14708, mcs1_mcs_mat1_6_n106}), .b ({new_AGEMA_signal_12837, new_AGEMA_signal_12836, mcs1_mcs_mat1_6_n105}), .c ({new_AGEMA_signal_15187, new_AGEMA_signal_15186, mcs_out[228]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U62 ( .a ({new_AGEMA_signal_12149, new_AGEMA_signal_12148, mcs1_mcs_mat1_6_mcs_out[120]}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_12837, new_AGEMA_signal_12836, mcs1_mcs_mat1_6_n105}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U61 ( .a ({new_AGEMA_signal_12857, new_AGEMA_signal_12856, mcs1_mcs_mat1_6_mcs_out[112]}), .b ({new_AGEMA_signal_14279, new_AGEMA_signal_14278, mcs1_mcs_mat1_6_mcs_out[116]}), .c ({new_AGEMA_signal_14709, new_AGEMA_signal_14708, mcs1_mcs_mat1_6_n106}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U60 ( .a ({new_AGEMA_signal_15189, new_AGEMA_signal_15188, mcs1_mcs_mat1_6_n104}), .b ({new_AGEMA_signal_13381, new_AGEMA_signal_13380, mcs1_mcs_mat1_6_n103}), .c ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, mcs_out[199]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U59 ( .a ({new_AGEMA_signal_12859, new_AGEMA_signal_12858, mcs1_mcs_mat1_6_mcs_out[111]}), .b ({new_AGEMA_signal_12869, new_AGEMA_signal_12868, mcs1_mcs_mat1_6_mcs_out[99]}), .c ({new_AGEMA_signal_13381, new_AGEMA_signal_13380, mcs1_mcs_mat1_6_n103}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U58 ( .a ({new_AGEMA_signal_14727, new_AGEMA_signal_14726, mcs1_mcs_mat1_6_mcs_out[103]}), .b ({new_AGEMA_signal_12161, new_AGEMA_signal_12160, mcs1_mcs_mat1_6_mcs_out[107]}), .c ({new_AGEMA_signal_15189, new_AGEMA_signal_15188, mcs1_mcs_mat1_6_n104}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U57 ( .a ({new_AGEMA_signal_14267, new_AGEMA_signal_14266, mcs1_mcs_mat1_6_n102}), .b ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, mcs1_mcs_mat1_6_n101}), .c ({new_AGEMA_signal_14711, new_AGEMA_signal_14710, mcs_out[198]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U56 ( .a ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, mcs1_mcs_mat1_6_mcs_out[110]}), .b ({new_AGEMA_signal_11207, new_AGEMA_signal_11206, mcs1_mcs_mat1_6_mcs_out[98]}), .c ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, mcs1_mcs_mat1_6_n101}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U55 ( .a ({new_AGEMA_signal_13843, new_AGEMA_signal_13842, mcs1_mcs_mat1_6_mcs_out[102]}), .b ({new_AGEMA_signal_12163, new_AGEMA_signal_12162, mcs1_mcs_mat1_6_mcs_out[106]}), .c ({new_AGEMA_signal_14267, new_AGEMA_signal_14266, mcs1_mcs_mat1_6_n102}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U54 ( .a ({new_AGEMA_signal_14713, new_AGEMA_signal_14712, mcs1_mcs_mat1_6_n100}), .b ({new_AGEMA_signal_13385, new_AGEMA_signal_13384, mcs1_mcs_mat1_6_n99}), .c ({new_AGEMA_signal_15191, new_AGEMA_signal_15190, mcs_out[197]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U53 ( .a ({new_AGEMA_signal_12863, new_AGEMA_signal_12862, mcs1_mcs_mat1_6_mcs_out[109]}), .b ({new_AGEMA_signal_9355, new_AGEMA_signal_9354, mcs1_mcs_mat1_6_mcs_out[97]}), .c ({new_AGEMA_signal_13385, new_AGEMA_signal_13384, mcs1_mcs_mat1_6_n99}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U52 ( .a ({new_AGEMA_signal_14283, new_AGEMA_signal_14282, mcs1_mcs_mat1_6_mcs_out[101]}), .b ({new_AGEMA_signal_12165, new_AGEMA_signal_12164, mcs1_mcs_mat1_6_mcs_out[105]}), .c ({new_AGEMA_signal_14713, new_AGEMA_signal_14712, mcs1_mcs_mat1_6_n100}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U51 ( .a ({new_AGEMA_signal_15193, new_AGEMA_signal_15192, mcs1_mcs_mat1_6_n98}), .b ({new_AGEMA_signal_14269, new_AGEMA_signal_14268, mcs1_mcs_mat1_6_n97}), .c ({new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs_out[196]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U50 ( .a ({new_AGEMA_signal_12865, new_AGEMA_signal_12864, mcs1_mcs_mat1_6_mcs_out[108]}), .b ({new_AGEMA_signal_13851, new_AGEMA_signal_13850, mcs1_mcs_mat1_6_mcs_out[96]}), .c ({new_AGEMA_signal_14269, new_AGEMA_signal_14268, mcs1_mcs_mat1_6_n97}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U49 ( .a ({new_AGEMA_signal_14729, new_AGEMA_signal_14728, mcs1_mcs_mat1_6_mcs_out[100]}), .b ({new_AGEMA_signal_12867, new_AGEMA_signal_12866, mcs1_mcs_mat1_6_mcs_out[104]}), .c ({new_AGEMA_signal_15193, new_AGEMA_signal_15192, mcs1_mcs_mat1_6_n98}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U48 ( .a ({new_AGEMA_signal_14271, new_AGEMA_signal_14270, mcs1_mcs_mat1_6_n96}), .b ({new_AGEMA_signal_12839, new_AGEMA_signal_12838, mcs1_mcs_mat1_6_n95}), .c ({new_AGEMA_signal_14715, new_AGEMA_signal_14714, mcs_out[167]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U47 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_12173, new_AGEMA_signal_12172, mcs1_mcs_mat1_6_mcs_out[95]}), .c ({new_AGEMA_signal_12839, new_AGEMA_signal_12838, mcs1_mcs_mat1_6_n95}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U46 ( .a ({new_AGEMA_signal_11211, new_AGEMA_signal_11210, mcs1_mcs_mat1_6_mcs_out[83]}), .b ({new_AGEMA_signal_13853, new_AGEMA_signal_13852, mcs1_mcs_mat1_6_mcs_out[87]}), .c ({new_AGEMA_signal_14271, new_AGEMA_signal_14270, mcs1_mcs_mat1_6_n96}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U45 ( .a ({new_AGEMA_signal_12137, new_AGEMA_signal_12136, mcs1_mcs_mat1_6_n94}), .b ({new_AGEMA_signal_11181, new_AGEMA_signal_11180, mcs1_mcs_mat1_6_n93}), .c ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, mcs_out[166]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U43 ( .a ({new_AGEMA_signal_11213, new_AGEMA_signal_11212, mcs1_mcs_mat1_6_mcs_out[82]}), .b ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_12137, new_AGEMA_signal_12136, mcs1_mcs_mat1_6_n94}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U42 ( .a ({new_AGEMA_signal_13387, new_AGEMA_signal_13386, mcs1_mcs_mat1_6_n92}), .b ({new_AGEMA_signal_11183, new_AGEMA_signal_11182, mcs1_mcs_mat1_6_n91}), .c ({new_AGEMA_signal_13831, new_AGEMA_signal_13830, mcs_out[165]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U41 ( .a ({new_AGEMA_signal_9367, new_AGEMA_signal_9366, mcs1_mcs_mat1_6_mcs_out[89]}), .b ({new_AGEMA_signal_10241, new_AGEMA_signal_10240, mcs1_mcs_mat1_6_mcs_out[93]}), .c ({new_AGEMA_signal_11183, new_AGEMA_signal_11182, mcs1_mcs_mat1_6_n91}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U40 ( .a ({new_AGEMA_signal_11215, new_AGEMA_signal_11214, mcs1_mcs_mat1_6_mcs_out[81]}), .b ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_13387, new_AGEMA_signal_13386, mcs1_mcs_mat1_6_n92}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U39 ( .a ({new_AGEMA_signal_14717, new_AGEMA_signal_14716, mcs1_mcs_mat1_6_n90}), .b ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, mcs1_mcs_mat1_6_n89}), .c ({new_AGEMA_signal_15195, new_AGEMA_signal_15194, mcs_out[164]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U38 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_12871, new_AGEMA_signal_12870, mcs1_mcs_mat1_6_mcs_out[92]}), .c ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, mcs1_mcs_mat1_6_n89}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U37 ( .a ({new_AGEMA_signal_12177, new_AGEMA_signal_12176, mcs1_mcs_mat1_6_mcs_out[80]}), .b ({new_AGEMA_signal_14287, new_AGEMA_signal_14286, mcs1_mcs_mat1_6_mcs_out[84]}), .c ({new_AGEMA_signal_14717, new_AGEMA_signal_14716, mcs1_mcs_mat1_6_n90}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U36 ( .a ({new_AGEMA_signal_12843, new_AGEMA_signal_12842, mcs1_mcs_mat1_6_n88}), .b ({new_AGEMA_signal_13833, new_AGEMA_signal_13832, mcs1_mcs_mat1_6_n87}), .c ({temp_next_s2[5], temp_next_s1[5], temp_next_s0[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U35 ( .a ({new_AGEMA_signal_13431, new_AGEMA_signal_13430, mcs1_mcs_mat1_6_mcs_out[5]}), .b ({new_AGEMA_signal_11287, new_AGEMA_signal_11286, mcs1_mcs_mat1_6_mcs_out[9]}), .c ({new_AGEMA_signal_13833, new_AGEMA_signal_13832, mcs1_mcs_mat1_6_n87}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U34 ( .a ({new_AGEMA_signal_12231, new_AGEMA_signal_12230, mcs1_mcs_mat1_6_mcs_out[13]}), .b ({new_AGEMA_signal_12243, new_AGEMA_signal_12242, mcs1_mcs_mat1_6_mcs_out[1]}), .c ({new_AGEMA_signal_12843, new_AGEMA_signal_12842, mcs1_mcs_mat1_6_n88}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U33 ( .a ({new_AGEMA_signal_15197, new_AGEMA_signal_15196, mcs1_mcs_mat1_6_n86}), .b ({new_AGEMA_signal_12845, new_AGEMA_signal_12844, mcs1_mcs_mat1_6_n85}), .c ({new_AGEMA_signal_15707, new_AGEMA_signal_15706, mcs_out[135]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U32 ( .a ({new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_6_mcs_out[75]}), .b ({new_AGEMA_signal_12179, new_AGEMA_signal_12178, mcs1_mcs_mat1_6_mcs_out[79]}), .c ({new_AGEMA_signal_12845, new_AGEMA_signal_12844, mcs1_mcs_mat1_6_n85}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U31 ( .a ({new_AGEMA_signal_12879, new_AGEMA_signal_12878, mcs1_mcs_mat1_6_mcs_out[67]}), .b ({new_AGEMA_signal_14731, new_AGEMA_signal_14730, mcs1_mcs_mat1_6_mcs_out[71]}), .c ({new_AGEMA_signal_15197, new_AGEMA_signal_15196, mcs1_mcs_mat1_6_n86}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U30 ( .a ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, mcs1_mcs_mat1_6_n84}), .b ({new_AGEMA_signal_13391, new_AGEMA_signal_13390, mcs1_mcs_mat1_6_n83}), .c ({new_AGEMA_signal_16119, new_AGEMA_signal_16118, mcs_out[134]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U29 ( .a ({new_AGEMA_signal_12875, new_AGEMA_signal_12874, mcs1_mcs_mat1_6_mcs_out[74]}), .b ({new_AGEMA_signal_8527, new_AGEMA_signal_8526, mcs1_mcs_mat1_6_mcs_out[78]}), .c ({new_AGEMA_signal_13391, new_AGEMA_signal_13390, mcs1_mcs_mat1_6_n83}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U28 ( .a ({new_AGEMA_signal_12189, new_AGEMA_signal_12188, mcs1_mcs_mat1_6_mcs_out[66]}), .b ({new_AGEMA_signal_15209, new_AGEMA_signal_15208, mcs1_mcs_mat1_6_mcs_out[70]}), .c ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, mcs1_mcs_mat1_6_n84}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U27 ( .a ({new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_6_n82}), .b ({new_AGEMA_signal_12139, new_AGEMA_signal_12138, mcs1_mcs_mat1_6_n81}), .c ({new_AGEMA_signal_16121, new_AGEMA_signal_16120, mcs_out[133]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U26 ( .a ({new_AGEMA_signal_11221, new_AGEMA_signal_11220, mcs1_mcs_mat1_6_mcs_out[73]}), .b ({new_AGEMA_signal_10253, new_AGEMA_signal_10252, mcs1_mcs_mat1_6_mcs_out[77]}), .c ({new_AGEMA_signal_12139, new_AGEMA_signal_12138, mcs1_mcs_mat1_6_n81}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U25 ( .a ({new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_6_mcs_out[65]}), .b ({new_AGEMA_signal_15211, new_AGEMA_signal_15210, mcs1_mcs_mat1_6_mcs_out[69]}), .c ({new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_6_n82}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U24 ( .a ({new_AGEMA_signal_15199, new_AGEMA_signal_15198, mcs1_mcs_mat1_6_n80}), .b ({new_AGEMA_signal_13393, new_AGEMA_signal_13392, mcs1_mcs_mat1_6_n79}), .c ({new_AGEMA_signal_15713, new_AGEMA_signal_15712, mcs_out[132]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U23 ( .a ({new_AGEMA_signal_12877, new_AGEMA_signal_12876, mcs1_mcs_mat1_6_mcs_out[72]}), .b ({new_AGEMA_signal_12873, new_AGEMA_signal_12872, mcs1_mcs_mat1_6_mcs_out[76]}), .c ({new_AGEMA_signal_13393, new_AGEMA_signal_13392, mcs1_mcs_mat1_6_n79}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U22 ( .a ({new_AGEMA_signal_13413, new_AGEMA_signal_13412, mcs1_mcs_mat1_6_mcs_out[64]}), .b ({new_AGEMA_signal_14735, new_AGEMA_signal_14734, mcs1_mcs_mat1_6_mcs_out[68]}), .c ({new_AGEMA_signal_15199, new_AGEMA_signal_15198, mcs1_mcs_mat1_6_n80}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U21 ( .a ({new_AGEMA_signal_15201, new_AGEMA_signal_15200, mcs1_mcs_mat1_6_n78}), .b ({new_AGEMA_signal_12847, new_AGEMA_signal_12846, mcs1_mcs_mat1_6_n77}), .c ({temp_next_s2[103], temp_next_s1[103], temp_next_s0[103]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U20 ( .a ({new_AGEMA_signal_11235, new_AGEMA_signal_11234, mcs1_mcs_mat1_6_mcs_out[59]}), .b ({new_AGEMA_signal_12193, new_AGEMA_signal_12192, mcs1_mcs_mat1_6_mcs_out[63]}), .c ({new_AGEMA_signal_12847, new_AGEMA_signal_12846, mcs1_mcs_mat1_6_n77}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U19 ( .a ({new_AGEMA_signal_10279, new_AGEMA_signal_10278, mcs1_mcs_mat1_6_mcs_out[51]}), .b ({new_AGEMA_signal_14737, new_AGEMA_signal_14736, mcs1_mcs_mat1_6_mcs_out[55]}), .c ({new_AGEMA_signal_15201, new_AGEMA_signal_15200, mcs1_mcs_mat1_6_n78}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U18 ( .a ({new_AGEMA_signal_15717, new_AGEMA_signal_15716, mcs1_mcs_mat1_6_n76}), .b ({new_AGEMA_signal_12141, new_AGEMA_signal_12140, mcs1_mcs_mat1_6_n75}), .c ({temp_next_s2[102], temp_next_s1[102], temp_next_s0[102]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U17 ( .a ({new_AGEMA_signal_10271, new_AGEMA_signal_10270, mcs1_mcs_mat1_6_mcs_out[58]}), .b ({new_AGEMA_signal_11229, new_AGEMA_signal_11228, mcs1_mcs_mat1_6_mcs_out[62]}), .c ({new_AGEMA_signal_12141, new_AGEMA_signal_12140, mcs1_mcs_mat1_6_n75}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U16 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_15213, new_AGEMA_signal_15212, mcs1_mcs_mat1_6_mcs_out[54]}), .c ({new_AGEMA_signal_15717, new_AGEMA_signal_15716, mcs1_mcs_mat1_6_n76}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U15 ( .a ({new_AGEMA_signal_15719, new_AGEMA_signal_15718, mcs1_mcs_mat1_6_n74}), .b ({new_AGEMA_signal_12143, new_AGEMA_signal_12142, mcs1_mcs_mat1_6_n73}), .c ({temp_next_s2[101], temp_next_s1[101], temp_next_s0[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U14 ( .a ({new_AGEMA_signal_11237, new_AGEMA_signal_11236, mcs1_mcs_mat1_6_mcs_out[57]}), .b ({new_AGEMA_signal_11231, new_AGEMA_signal_11230, mcs1_mcs_mat1_6_mcs_out[61]}), .c ({new_AGEMA_signal_12143, new_AGEMA_signal_12142, mcs1_mcs_mat1_6_n73}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U13 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_15215, new_AGEMA_signal_15214, mcs1_mcs_mat1_6_mcs_out[53]}), .c ({new_AGEMA_signal_15719, new_AGEMA_signal_15718, mcs1_mcs_mat1_6_n74}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U12 ( .a ({new_AGEMA_signal_15203, new_AGEMA_signal_15202, mcs1_mcs_mat1_6_n72}), .b ({new_AGEMA_signal_13395, new_AGEMA_signal_13394, mcs1_mcs_mat1_6_n71}), .c ({temp_next_s2[100], temp_next_s1[100], temp_next_s0[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U11 ( .a ({new_AGEMA_signal_12197, new_AGEMA_signal_12196, mcs1_mcs_mat1_6_mcs_out[56]}), .b ({new_AGEMA_signal_12883, new_AGEMA_signal_12882, mcs1_mcs_mat1_6_mcs_out[60]}), .c ({new_AGEMA_signal_13395, new_AGEMA_signal_13394, mcs1_mcs_mat1_6_n71}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U10 ( .a ({new_AGEMA_signal_11243, new_AGEMA_signal_11242, mcs1_mcs_mat1_6_mcs_out[48]}), .b ({new_AGEMA_signal_14741, new_AGEMA_signal_14740, mcs1_mcs_mat1_6_mcs_out[52]}), .c ({new_AGEMA_signal_15203, new_AGEMA_signal_15202, mcs1_mcs_mat1_6_n72}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U9 ( .a ({new_AGEMA_signal_15723, new_AGEMA_signal_15722, mcs1_mcs_mat1_6_n70}), .b ({new_AGEMA_signal_12849, new_AGEMA_signal_12848, mcs1_mcs_mat1_6_n69}), .c ({temp_next_s2[71], temp_next_s1[71], temp_next_s0[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U8 ( .a ({new_AGEMA_signal_12203, new_AGEMA_signal_12202, mcs1_mcs_mat1_6_mcs_out[43]}), .b ({new_AGEMA_signal_12201, new_AGEMA_signal_12200, mcs1_mcs_mat1_6_mcs_out[47]}), .c ({new_AGEMA_signal_12849, new_AGEMA_signal_12848, mcs1_mcs_mat1_6_n69}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U7 ( .a ({new_AGEMA_signal_12211, new_AGEMA_signal_12210, mcs1_mcs_mat1_6_mcs_out[35]}), .b ({new_AGEMA_signal_15217, new_AGEMA_signal_15216, mcs1_mcs_mat1_6_mcs_out[39]}), .c ({new_AGEMA_signal_15723, new_AGEMA_signal_15722, mcs1_mcs_mat1_6_n70}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U6 ( .a ({new_AGEMA_signal_14275, new_AGEMA_signal_14274, mcs1_mcs_mat1_6_n68}), .b ({new_AGEMA_signal_12851, new_AGEMA_signal_12850, mcs1_mcs_mat1_6_n67}), .c ({temp_next_s2[70], temp_next_s1[70], temp_next_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U5 ( .a ({new_AGEMA_signal_12205, new_AGEMA_signal_12204, mcs1_mcs_mat1_6_mcs_out[42]}), .b ({new_AGEMA_signal_9381, new_AGEMA_signal_9380, mcs1_mcs_mat1_6_mcs_out[46]}), .c ({new_AGEMA_signal_12851, new_AGEMA_signal_12850, mcs1_mcs_mat1_6_n67}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U4 ( .a ({new_AGEMA_signal_11257, new_AGEMA_signal_11256, mcs1_mcs_mat1_6_mcs_out[34]}), .b ({new_AGEMA_signal_13869, new_AGEMA_signal_13868, mcs1_mcs_mat1_6_mcs_out[38]}), .c ({new_AGEMA_signal_14275, new_AGEMA_signal_14274, mcs1_mcs_mat1_6_n68}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U3 ( .a ({new_AGEMA_signal_13835, new_AGEMA_signal_13834, mcs1_mcs_mat1_6_n66}), .b ({new_AGEMA_signal_16379, new_AGEMA_signal_16378, mcs1_mcs_mat1_6_n65}), .c ({temp_next_s2[4], temp_next_s1[4], temp_next_s0[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U2 ( .a ({new_AGEMA_signal_16129, new_AGEMA_signal_16128, mcs1_mcs_mat1_6_mcs_out[4]}), .b ({new_AGEMA_signal_12903, new_AGEMA_signal_12902, mcs1_mcs_mat1_6_mcs_out[8]}), .c ({new_AGEMA_signal_16379, new_AGEMA_signal_16378, mcs1_mcs_mat1_6_n65}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_U1 ( .a ({new_AGEMA_signal_12245, new_AGEMA_signal_12244, mcs1_mcs_mat1_6_mcs_out[0]}), .b ({new_AGEMA_signal_13429, new_AGEMA_signal_13428, mcs1_mcs_mat1_6_mcs_out[12]}), .c ({new_AGEMA_signal_13835, new_AGEMA_signal_13834, mcs1_mcs_mat1_6_n66}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_12145, new_AGEMA_signal_12144, mcs1_mcs_mat1_6_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_12853, new_AGEMA_signal_12852, mcs1_mcs_mat1_6_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_11185, new_AGEMA_signal_11184, mcs1_mcs_mat1_6_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_7921, new_AGEMA_signal_7920, mcs1_mcs_mat1_6_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_12145, new_AGEMA_signal_12144, mcs1_mcs_mat1_6_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_8507, new_AGEMA_signal_8506, mcs1_mcs_mat1_6_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_9341, new_AGEMA_signal_9340, mcs1_mcs_mat1_6_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, mcs1_mcs_mat1_6_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_8509, new_AGEMA_signal_8508, mcs1_mcs_mat1_6_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .c ({new_AGEMA_signal_9341, new_AGEMA_signal_9340, mcs1_mcs_mat1_6_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_12147, new_AGEMA_signal_12146, mcs1_mcs_mat1_6_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .c ({new_AGEMA_signal_12855, new_AGEMA_signal_12854, mcs1_mcs_mat1_6_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_11185, new_AGEMA_signal_11184, mcs1_mcs_mat1_6_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_12147, new_AGEMA_signal_12146, mcs1_mcs_mat1_6_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_10221, new_AGEMA_signal_10220, mcs1_mcs_mat1_6_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9343, new_AGEMA_signal_9342, mcs1_mcs_mat1_6_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_11185, new_AGEMA_signal_11184, mcs1_mcs_mat1_6_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_11187, new_AGEMA_signal_11186, mcs1_mcs_mat1_6_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_12149, new_AGEMA_signal_12148, mcs1_mcs_mat1_6_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_10221, new_AGEMA_signal_10220, mcs1_mcs_mat1_6_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_8509, new_AGEMA_signal_8508, mcs1_mcs_mat1_6_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_11187, new_AGEMA_signal_11186, mcs1_mcs_mat1_6_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2858], Fresh[2857], Fresh[2856]}), .c ({new_AGEMA_signal_10221, new_AGEMA_signal_10220, mcs1_mcs_mat1_6_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2861], Fresh[2860], Fresh[2859]}), .c ({new_AGEMA_signal_8509, new_AGEMA_signal_8508, mcs1_mcs_mat1_6_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2864], Fresh[2863], Fresh[2862]}), .c ({new_AGEMA_signal_9343, new_AGEMA_signal_9342, mcs1_mcs_mat1_6_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_14721, new_AGEMA_signal_14720, mcs1_mcs_mat1_6_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .c ({new_AGEMA_signal_15205, new_AGEMA_signal_15204, mcs1_mcs_mat1_6_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_14277, new_AGEMA_signal_14276, mcs1_mcs_mat1_6_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_13401, new_AGEMA_signal_13400, mcs1_mcs_mat1_6_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_14721, new_AGEMA_signal_14720, mcs1_mcs_mat1_6_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_14723, new_AGEMA_signal_14722, mcs1_mcs_mat1_6_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_13839, new_AGEMA_signal_13838, mcs1_mcs_mat1_6_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_15207, new_AGEMA_signal_15206, mcs1_mcs_mat1_6_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_14277, new_AGEMA_signal_14276, mcs1_mcs_mat1_6_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .c ({new_AGEMA_signal_14723, new_AGEMA_signal_14722, mcs1_mcs_mat1_6_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_14277, new_AGEMA_signal_14276, mcs1_mcs_mat1_6_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_13837, new_AGEMA_signal_13836, mcs1_mcs_mat1_6_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_14725, new_AGEMA_signal_14724, mcs1_mcs_mat1_6_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_13841, new_AGEMA_signal_13840, mcs1_mcs_mat1_6_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_12151, new_AGEMA_signal_12150, mcs1_mcs_mat1_6_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_14277, new_AGEMA_signal_14276, mcs1_mcs_mat1_6_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_13399, new_AGEMA_signal_13398, mcs1_mcs_mat1_6_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_13839, new_AGEMA_signal_13838, mcs1_mcs_mat1_6_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_14279, new_AGEMA_signal_14278, mcs1_mcs_mat1_6_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_11189, new_AGEMA_signal_11188, mcs1_mcs_mat1_6_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_13401, new_AGEMA_signal_13400, mcs1_mcs_mat1_6_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_13839, new_AGEMA_signal_13838, mcs1_mcs_mat1_6_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_12151, new_AGEMA_signal_12150, mcs1_mcs_mat1_6_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_13399, new_AGEMA_signal_13398, mcs1_mcs_mat1_6_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2867], Fresh[2866], Fresh[2865]}), .c ({new_AGEMA_signal_13841, new_AGEMA_signal_13840, mcs1_mcs_mat1_6_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2870], Fresh[2869], Fresh[2868]}), .c ({new_AGEMA_signal_12151, new_AGEMA_signal_12150, mcs1_mcs_mat1_6_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2873], Fresh[2872], Fresh[2871]}), .c ({new_AGEMA_signal_13401, new_AGEMA_signal_13400, mcs1_mcs_mat1_6_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_11193, new_AGEMA_signal_11192, mcs1_mcs_mat1_6_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_8511, new_AGEMA_signal_8510, mcs1_mcs_mat1_6_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_12153, new_AGEMA_signal_12152, mcs1_mcs_mat1_6_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_9345, new_AGEMA_signal_9344, mcs1_mcs_mat1_6_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_9347, new_AGEMA_signal_9346, mcs1_mcs_mat1_6_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_10223, new_AGEMA_signal_10222, mcs1_mcs_mat1_6_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_11195, new_AGEMA_signal_11194, mcs1_mcs_mat1_6_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_12155, new_AGEMA_signal_12154, mcs1_mcs_mat1_6_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_12857, new_AGEMA_signal_12856, mcs1_mcs_mat1_6_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_11193, new_AGEMA_signal_11192, mcs1_mcs_mat1_6_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_12155, new_AGEMA_signal_12154, mcs1_mcs_mat1_6_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_7923, new_AGEMA_signal_7922, mcs1_mcs_mat1_6_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_10227, new_AGEMA_signal_10226, mcs1_mcs_mat1_6_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_11193, new_AGEMA_signal_11192, mcs1_mcs_mat1_6_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_8513, new_AGEMA_signal_8512, mcs1_mcs_mat1_6_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, mcs1_mcs_mat1_6_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_11195, new_AGEMA_signal_11194, mcs1_mcs_mat1_6_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2876], Fresh[2875], Fresh[2874]}), .c ({new_AGEMA_signal_10227, new_AGEMA_signal_10226, mcs1_mcs_mat1_6_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2879], Fresh[2878], Fresh[2877]}), .c ({new_AGEMA_signal_8513, new_AGEMA_signal_8512, mcs1_mcs_mat1_6_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({new_AGEMA_signal_9347, new_AGEMA_signal_9346, mcs1_mcs_mat1_6_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({new_AGEMA_signal_12157, new_AGEMA_signal_12156, mcs1_mcs_mat1_6_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12859, new_AGEMA_signal_12858, mcs1_mcs_mat1_6_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({new_AGEMA_signal_12159, new_AGEMA_signal_12158, mcs1_mcs_mat1_6_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, mcs1_mcs_mat1_6_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_9349, new_AGEMA_signal_9348, mcs1_mcs_mat1_6_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_12157, new_AGEMA_signal_12156, mcs1_mcs_mat1_6_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12863, new_AGEMA_signal_12862, mcs1_mcs_mat1_6_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_8515, new_AGEMA_signal_8514, mcs1_mcs_mat1_6_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_11197, new_AGEMA_signal_11196, mcs1_mcs_mat1_6_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_12157, new_AGEMA_signal_12156, mcs1_mcs_mat1_6_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_10229, new_AGEMA_signal_10228, mcs1_mcs_mat1_6_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_12159, new_AGEMA_signal_12158, mcs1_mcs_mat1_6_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12865, new_AGEMA_signal_12864, mcs1_mcs_mat1_6_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_11199, new_AGEMA_signal_11198, mcs1_mcs_mat1_6_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_12159, new_AGEMA_signal_12158, mcs1_mcs_mat1_6_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_9349, new_AGEMA_signal_9348, mcs1_mcs_mat1_6_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, mcs1_mcs_mat1_6_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_11199, new_AGEMA_signal_11198, mcs1_mcs_mat1_6_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2885], Fresh[2884], Fresh[2883]}), .c ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, mcs1_mcs_mat1_6_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2888], Fresh[2887], Fresh[2886]}), .c ({new_AGEMA_signal_8515, new_AGEMA_signal_8514, mcs1_mcs_mat1_6_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2891], Fresh[2890], Fresh[2889]}), .c ({new_AGEMA_signal_9349, new_AGEMA_signal_9348, mcs1_mcs_mat1_6_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_11203, new_AGEMA_signal_11202, mcs1_mcs_mat1_6_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_11201, new_AGEMA_signal_11200, mcs1_mcs_mat1_6_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_12161, new_AGEMA_signal_12160, mcs1_mcs_mat1_6_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_11201, new_AGEMA_signal_11200, mcs1_mcs_mat1_6_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_9351, new_AGEMA_signal_9350, mcs1_mcs_mat1_6_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_12163, new_AGEMA_signal_12162, mcs1_mcs_mat1_6_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, mcs1_mcs_mat1_6_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .c ({new_AGEMA_signal_9351, new_AGEMA_signal_9350, mcs1_mcs_mat1_6_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_11201, new_AGEMA_signal_11200, mcs1_mcs_mat1_6_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_12165, new_AGEMA_signal_12164, mcs1_mcs_mat1_6_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_10235, new_AGEMA_signal_10234, mcs1_mcs_mat1_6_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_7927, new_AGEMA_signal_7926, mcs1_mcs_mat1_6_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_11201, new_AGEMA_signal_11200, mcs1_mcs_mat1_6_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_12167, new_AGEMA_signal_12166, mcs1_mcs_mat1_6_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_12867, new_AGEMA_signal_12866, mcs1_mcs_mat1_6_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_11203, new_AGEMA_signal_11202, mcs1_mcs_mat1_6_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_10235, new_AGEMA_signal_10234, mcs1_mcs_mat1_6_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_12167, new_AGEMA_signal_12166, mcs1_mcs_mat1_6_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_10233, new_AGEMA_signal_10232, mcs1_mcs_mat1_6_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .c ({new_AGEMA_signal_11203, new_AGEMA_signal_11202, mcs1_mcs_mat1_6_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, mcs1_mcs_mat1_6_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_9353, new_AGEMA_signal_9352, mcs1_mcs_mat1_6_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_10233, new_AGEMA_signal_10232, mcs1_mcs_mat1_6_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2894], Fresh[2893], Fresh[2892]}), .c ({new_AGEMA_signal_10235, new_AGEMA_signal_10234, mcs1_mcs_mat1_6_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2897], Fresh[2896], Fresh[2895]}), .c ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, mcs1_mcs_mat1_6_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2900], Fresh[2899], Fresh[2898]}), .c ({new_AGEMA_signal_9353, new_AGEMA_signal_9352, mcs1_mcs_mat1_6_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_13403, new_AGEMA_signal_13402, mcs1_mcs_mat1_6_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_14281, new_AGEMA_signal_14280, mcs1_mcs_mat1_6_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_14727, new_AGEMA_signal_14726, mcs1_mcs_mat1_6_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_13849, new_AGEMA_signal_13848, mcs1_mcs_mat1_6_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_14281, new_AGEMA_signal_14280, mcs1_mcs_mat1_6_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_13845, new_AGEMA_signal_13844, mcs1_mcs_mat1_6_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_13405, new_AGEMA_signal_13404, mcs1_mcs_mat1_6_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_14283, new_AGEMA_signal_14282, mcs1_mcs_mat1_6_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_13847, new_AGEMA_signal_13846, mcs1_mcs_mat1_6_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_14285, new_AGEMA_signal_14284, mcs1_mcs_mat1_6_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_14729, new_AGEMA_signal_14728, mcs1_mcs_mat1_6_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_11205, new_AGEMA_signal_11204, mcs1_mcs_mat1_6_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_13849, new_AGEMA_signal_13848, mcs1_mcs_mat1_6_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_14285, new_AGEMA_signal_14284, mcs1_mcs_mat1_6_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_12169, new_AGEMA_signal_12168, mcs1_mcs_mat1_6_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .c ({new_AGEMA_signal_13847, new_AGEMA_signal_13846, mcs1_mcs_mat1_6_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2903], Fresh[2902], Fresh[2901]}), .c ({new_AGEMA_signal_13849, new_AGEMA_signal_13848, mcs1_mcs_mat1_6_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2906], Fresh[2905], Fresh[2904]}), .c ({new_AGEMA_signal_12169, new_AGEMA_signal_12168, mcs1_mcs_mat1_6_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2909], Fresh[2908], Fresh[2907]}), .c ({new_AGEMA_signal_13405, new_AGEMA_signal_13404, mcs1_mcs_mat1_6_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_13407, new_AGEMA_signal_13406, mcs1_mcs_mat1_6_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_9357, new_AGEMA_signal_9356, mcs1_mcs_mat1_6_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_13851, new_AGEMA_signal_13850, mcs1_mcs_mat1_6_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_12869, new_AGEMA_signal_12868, mcs1_mcs_mat1_6_mcs_out[99]}), .b ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .c ({new_AGEMA_signal_13407, new_AGEMA_signal_13406, mcs1_mcs_mat1_6_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, mcs1_mcs_mat1_6_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .c ({new_AGEMA_signal_12869, new_AGEMA_signal_12868, mcs1_mcs_mat1_6_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_11207, new_AGEMA_signal_11206, mcs1_mcs_mat1_6_mcs_out[98]}), .b ({new_AGEMA_signal_8521, new_AGEMA_signal_8520, mcs1_mcs_mat1_6_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, mcs1_mcs_mat1_6_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_8519, new_AGEMA_signal_8518, mcs1_mcs_mat1_6_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, mcs1_mcs_mat1_6_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_11207, new_AGEMA_signal_11206, mcs1_mcs_mat1_6_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, mcs1_mcs_mat1_6_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2915], Fresh[2914], Fresh[2913]}), .c ({new_AGEMA_signal_8521, new_AGEMA_signal_8520, mcs1_mcs_mat1_6_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2918], Fresh[2917], Fresh[2916]}), .c ({new_AGEMA_signal_9357, new_AGEMA_signal_9356, mcs1_mcs_mat1_6_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_11209, new_AGEMA_signal_11208, mcs1_mcs_mat1_6_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_12173, new_AGEMA_signal_12172, mcs1_mcs_mat1_6_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_9361, new_AGEMA_signal_9360, mcs1_mcs_mat1_6_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_9363, new_AGEMA_signal_9362, mcs1_mcs_mat1_6_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_10241, new_AGEMA_signal_10240, mcs1_mcs_mat1_6_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_12175, new_AGEMA_signal_12174, mcs1_mcs_mat1_6_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_8523, new_AGEMA_signal_8522, mcs1_mcs_mat1_6_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_12871, new_AGEMA_signal_12870, mcs1_mcs_mat1_6_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_11209, new_AGEMA_signal_11208, mcs1_mcs_mat1_6_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_12175, new_AGEMA_signal_12174, mcs1_mcs_mat1_6_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_7931, new_AGEMA_signal_7930, mcs1_mcs_mat1_6_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, mcs1_mcs_mat1_6_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_11209, new_AGEMA_signal_11208, mcs1_mcs_mat1_6_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2921], Fresh[2920], Fresh[2919]}), .c ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, mcs1_mcs_mat1_6_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2924], Fresh[2923], Fresh[2922]}), .c ({new_AGEMA_signal_8523, new_AGEMA_signal_8522, mcs1_mcs_mat1_6_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2927], Fresh[2926], Fresh[2925]}), .c ({new_AGEMA_signal_9363, new_AGEMA_signal_9362, mcs1_mcs_mat1_6_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, mcs1_mcs_mat1_6_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_6_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_11211, new_AGEMA_signal_11210, mcs1_mcs_mat1_6_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_6_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_7933, new_AGEMA_signal_7932, mcs1_mcs_mat1_6_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_11213, new_AGEMA_signal_11212, mcs1_mcs_mat1_6_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_9369, new_AGEMA_signal_9368, mcs1_mcs_mat1_6_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_6_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_10247, new_AGEMA_signal_10246, mcs1_mcs_mat1_6_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_11215, new_AGEMA_signal_11214, mcs1_mcs_mat1_6_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_8525, new_AGEMA_signal_8524, mcs1_mcs_mat1_6_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_9369, new_AGEMA_signal_9368, mcs1_mcs_mat1_6_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_10247, new_AGEMA_signal_10246, mcs1_mcs_mat1_6_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_11217, new_AGEMA_signal_11216, mcs1_mcs_mat1_6_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .c ({new_AGEMA_signal_12177, new_AGEMA_signal_12176, mcs1_mcs_mat1_6_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, mcs1_mcs_mat1_6_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_8525, new_AGEMA_signal_8524, mcs1_mcs_mat1_6_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_11217, new_AGEMA_signal_11216, mcs1_mcs_mat1_6_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2930], Fresh[2929], Fresh[2928]}), .c ({new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_6_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2933], Fresh[2932], Fresh[2931]}), .c ({new_AGEMA_signal_8525, new_AGEMA_signal_8524, mcs1_mcs_mat1_6_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2936], Fresh[2935], Fresh[2934]}), .c ({new_AGEMA_signal_9369, new_AGEMA_signal_9368, mcs1_mcs_mat1_6_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_11219, new_AGEMA_signal_11218, mcs1_mcs_mat1_6_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_12179, new_AGEMA_signal_12178, mcs1_mcs_mat1_6_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_9371, new_AGEMA_signal_9370, mcs1_mcs_mat1_6_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_10253, new_AGEMA_signal_10252, mcs1_mcs_mat1_6_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_12181, new_AGEMA_signal_12180, mcs1_mcs_mat1_6_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_8529, new_AGEMA_signal_8528, mcs1_mcs_mat1_6_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_12873, new_AGEMA_signal_12872, mcs1_mcs_mat1_6_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_11219, new_AGEMA_signal_11218, mcs1_mcs_mat1_6_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .c ({new_AGEMA_signal_12181, new_AGEMA_signal_12180, mcs1_mcs_mat1_6_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, mcs1_mcs_mat1_6_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, mcs1_mcs_mat1_6_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_11219, new_AGEMA_signal_11218, mcs1_mcs_mat1_6_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2939], Fresh[2938], Fresh[2937]}), .c ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, mcs1_mcs_mat1_6_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({new_AGEMA_signal_8529, new_AGEMA_signal_8528, mcs1_mcs_mat1_6_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2945], Fresh[2944], Fresh[2943]}), .c ({new_AGEMA_signal_9371, new_AGEMA_signal_9370, mcs1_mcs_mat1_6_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_12183, new_AGEMA_signal_12182, mcs1_mcs_mat1_6_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_12875, new_AGEMA_signal_12874, mcs1_mcs_mat1_6_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_11223, new_AGEMA_signal_11222, mcs1_mcs_mat1_6_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_10259, new_AGEMA_signal_10258, mcs1_mcs_mat1_6_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_12183, new_AGEMA_signal_12182, mcs1_mcs_mat1_6_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_8807, new_AGEMA_signal_8806, mcs1_mcs_mat1_6_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_6_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_10259, new_AGEMA_signal_10258, mcs1_mcs_mat1_6_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_8807, new_AGEMA_signal_8806, mcs1_mcs_mat1_6_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_11221, new_AGEMA_signal_11220, mcs1_mcs_mat1_6_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_8531, new_AGEMA_signal_8530, mcs1_mcs_mat1_6_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_8533, new_AGEMA_signal_8532, mcs1_mcs_mat1_6_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_8807, new_AGEMA_signal_8806, mcs1_mcs_mat1_6_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_9373, new_AGEMA_signal_9372, mcs1_mcs_mat1_6_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .c ({new_AGEMA_signal_10259, new_AGEMA_signal_10258, mcs1_mcs_mat1_6_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_12185, new_AGEMA_signal_12184, mcs1_mcs_mat1_6_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_8531, new_AGEMA_signal_8530, mcs1_mcs_mat1_6_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_12877, new_AGEMA_signal_12876, mcs1_mcs_mat1_6_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_11223, new_AGEMA_signal_11222, mcs1_mcs_mat1_6_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_9373, new_AGEMA_signal_9372, mcs1_mcs_mat1_6_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_12185, new_AGEMA_signal_12184, mcs1_mcs_mat1_6_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .b ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, mcs1_mcs_mat1_6_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_11223, new_AGEMA_signal_11222, mcs1_mcs_mat1_6_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2948], Fresh[2947], Fresh[2946]}), .c ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, mcs1_mcs_mat1_6_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2951], Fresh[2950], Fresh[2949]}), .c ({new_AGEMA_signal_8533, new_AGEMA_signal_8532, mcs1_mcs_mat1_6_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2954], Fresh[2953], Fresh[2952]}), .c ({new_AGEMA_signal_9373, new_AGEMA_signal_9372, mcs1_mcs_mat1_6_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_14289, new_AGEMA_signal_14288, mcs1_mcs_mat1_6_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_13409, new_AGEMA_signal_13408, mcs1_mcs_mat1_6_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_14731, new_AGEMA_signal_14730, mcs1_mcs_mat1_6_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_13857, new_AGEMA_signal_13856, mcs1_mcs_mat1_6_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_14733, new_AGEMA_signal_14732, mcs1_mcs_mat1_6_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_15209, new_AGEMA_signal_15208, mcs1_mcs_mat1_6_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_14289, new_AGEMA_signal_14288, mcs1_mcs_mat1_6_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_14733, new_AGEMA_signal_14732, mcs1_mcs_mat1_6_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_15211, new_AGEMA_signal_15210, mcs1_mcs_mat1_6_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_13409, new_AGEMA_signal_13408, mcs1_mcs_mat1_6_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_14291, new_AGEMA_signal_14290, mcs1_mcs_mat1_6_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_14733, new_AGEMA_signal_14732, mcs1_mcs_mat1_6_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({new_AGEMA_signal_12187, new_AGEMA_signal_12186, mcs1_mcs_mat1_6_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_13409, new_AGEMA_signal_13408, mcs1_mcs_mat1_6_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_13855, new_AGEMA_signal_13854, mcs1_mcs_mat1_6_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .c ({new_AGEMA_signal_14289, new_AGEMA_signal_14288, mcs1_mcs_mat1_6_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_13411, new_AGEMA_signal_13410, mcs1_mcs_mat1_6_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_11225, new_AGEMA_signal_11224, mcs1_mcs_mat1_6_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_13855, new_AGEMA_signal_13854, mcs1_mcs_mat1_6_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_14291, new_AGEMA_signal_14290, mcs1_mcs_mat1_6_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_13857, new_AGEMA_signal_13856, mcs1_mcs_mat1_6_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_14735, new_AGEMA_signal_14734, mcs1_mcs_mat1_6_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_13411, new_AGEMA_signal_13410, mcs1_mcs_mat1_6_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_13857, new_AGEMA_signal_13856, mcs1_mcs_mat1_6_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({new_AGEMA_signal_13859, new_AGEMA_signal_13858, mcs1_mcs_mat1_6_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_14291, new_AGEMA_signal_14290, mcs1_mcs_mat1_6_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2957], Fresh[2956], Fresh[2955]}), .c ({new_AGEMA_signal_13859, new_AGEMA_signal_13858, mcs1_mcs_mat1_6_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2960], Fresh[2959], Fresh[2958]}), .c ({new_AGEMA_signal_12187, new_AGEMA_signal_12186, mcs1_mcs_mat1_6_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2963], Fresh[2962], Fresh[2961]}), .c ({new_AGEMA_signal_13411, new_AGEMA_signal_13410, mcs1_mcs_mat1_6_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_12191, new_AGEMA_signal_12190, mcs1_mcs_mat1_6_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_12879, new_AGEMA_signal_12878, mcs1_mcs_mat1_6_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({new_AGEMA_signal_11227, new_AGEMA_signal_11226, mcs1_mcs_mat1_6_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_12189, new_AGEMA_signal_12188, mcs1_mcs_mat1_6_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_12881, new_AGEMA_signal_12880, mcs1_mcs_mat1_6_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_9375, new_AGEMA_signal_9374, mcs1_mcs_mat1_6_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_13413, new_AGEMA_signal_13412, mcs1_mcs_mat1_6_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_12191, new_AGEMA_signal_12190, mcs1_mcs_mat1_6_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .c ({new_AGEMA_signal_12881, new_AGEMA_signal_12880, mcs1_mcs_mat1_6_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_8535, new_AGEMA_signal_8534, mcs1_mcs_mat1_6_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_11227, new_AGEMA_signal_11226, mcs1_mcs_mat1_6_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_12191, new_AGEMA_signal_12190, mcs1_mcs_mat1_6_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_7939, new_AGEMA_signal_7938, mcs1_mcs_mat1_6_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_10265, new_AGEMA_signal_10264, mcs1_mcs_mat1_6_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_11227, new_AGEMA_signal_11226, mcs1_mcs_mat1_6_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2966], Fresh[2965], Fresh[2964]}), .c ({new_AGEMA_signal_10265, new_AGEMA_signal_10264, mcs1_mcs_mat1_6_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2969], Fresh[2968], Fresh[2967]}), .c ({new_AGEMA_signal_8535, new_AGEMA_signal_8534, mcs1_mcs_mat1_6_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({new_AGEMA_signal_9375, new_AGEMA_signal_9374, mcs1_mcs_mat1_6_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_11233, new_AGEMA_signal_11232, mcs1_mcs_mat1_6_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_9377, new_AGEMA_signal_9376, mcs1_mcs_mat1_6_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_12193, new_AGEMA_signal_12192, mcs1_mcs_mat1_6_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_8537, new_AGEMA_signal_8536, mcs1_mcs_mat1_6_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, mcs1_mcs_mat1_6_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_11229, new_AGEMA_signal_11228, mcs1_mcs_mat1_6_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_6_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_11231, new_AGEMA_signal_11230, mcs1_mcs_mat1_6_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2975], Fresh[2974], Fresh[2973]}), .c ({new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_6_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2978], Fresh[2977], Fresh[2976]}), .c ({new_AGEMA_signal_8537, new_AGEMA_signal_8536, mcs1_mcs_mat1_6_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2981], Fresh[2980], Fresh[2979]}), .c ({new_AGEMA_signal_9377, new_AGEMA_signal_9376, mcs1_mcs_mat1_6_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_8541, new_AGEMA_signal_8540, mcs1_mcs_mat1_6_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_9379, new_AGEMA_signal_9378, mcs1_mcs_mat1_6_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_10271, new_AGEMA_signal_10270, mcs1_mcs_mat1_6_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_8543, new_AGEMA_signal_8542, mcs1_mcs_mat1_6_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, mcs1_mcs_mat1_6_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_11237, new_AGEMA_signal_11236, mcs1_mcs_mat1_6_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_11239, new_AGEMA_signal_11238, mcs1_mcs_mat1_6_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_10275, new_AGEMA_signal_10274, mcs1_mcs_mat1_6_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_12197, new_AGEMA_signal_12196, mcs1_mcs_mat1_6_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_10277, new_AGEMA_signal_10276, mcs1_mcs_mat1_6_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_11239, new_AGEMA_signal_11238, mcs1_mcs_mat1_6_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2984], Fresh[2983], Fresh[2982]}), .c ({new_AGEMA_signal_10277, new_AGEMA_signal_10276, mcs1_mcs_mat1_6_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2987], Fresh[2986], Fresh[2985]}), .c ({new_AGEMA_signal_8543, new_AGEMA_signal_8542, mcs1_mcs_mat1_6_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2990], Fresh[2989], Fresh[2988]}), .c ({new_AGEMA_signal_9379, new_AGEMA_signal_9378, mcs1_mcs_mat1_6_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_13863, new_AGEMA_signal_13862, mcs1_mcs_mat1_6_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_14293, new_AGEMA_signal_14292, mcs1_mcs_mat1_6_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_14737, new_AGEMA_signal_14736, mcs1_mcs_mat1_6_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_14739, new_AGEMA_signal_14738, mcs1_mcs_mat1_6_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_13861, new_AGEMA_signal_13860, mcs1_mcs_mat1_6_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_15213, new_AGEMA_signal_15212, mcs1_mcs_mat1_6_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_13415, new_AGEMA_signal_13414, mcs1_mcs_mat1_6_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_13861, new_AGEMA_signal_13860, mcs1_mcs_mat1_6_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({new_AGEMA_signal_14739, new_AGEMA_signal_14738, mcs1_mcs_mat1_6_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_15215, new_AGEMA_signal_15214, mcs1_mcs_mat1_6_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_11241, new_AGEMA_signal_11240, mcs1_mcs_mat1_6_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_14293, new_AGEMA_signal_14292, mcs1_mcs_mat1_6_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_14739, new_AGEMA_signal_14738, mcs1_mcs_mat1_6_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_12199, new_AGEMA_signal_12198, mcs1_mcs_mat1_6_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_13867, new_AGEMA_signal_13866, mcs1_mcs_mat1_6_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_14293, new_AGEMA_signal_14292, mcs1_mcs_mat1_6_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_13865, new_AGEMA_signal_13864, mcs1_mcs_mat1_6_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_14295, new_AGEMA_signal_14294, mcs1_mcs_mat1_6_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_14741, new_AGEMA_signal_14740, mcs1_mcs_mat1_6_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_13863, new_AGEMA_signal_13862, mcs1_mcs_mat1_6_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_12199, new_AGEMA_signal_12198, mcs1_mcs_mat1_6_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_14295, new_AGEMA_signal_14294, mcs1_mcs_mat1_6_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_13415, new_AGEMA_signal_13414, mcs1_mcs_mat1_6_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_13863, new_AGEMA_signal_13862, mcs1_mcs_mat1_6_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2993], Fresh[2992], Fresh[2991]}), .c ({new_AGEMA_signal_13867, new_AGEMA_signal_13866, mcs1_mcs_mat1_6_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2996], Fresh[2995], Fresh[2994]}), .c ({new_AGEMA_signal_12199, new_AGEMA_signal_12198, mcs1_mcs_mat1_6_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2999], Fresh[2998], Fresh[2997]}), .c ({new_AGEMA_signal_13415, new_AGEMA_signal_13414, mcs1_mcs_mat1_6_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_9383, new_AGEMA_signal_9382, mcs1_mcs_mat1_6_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_10281, new_AGEMA_signal_10280, mcs1_mcs_mat1_6_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_12885, new_AGEMA_signal_12884, mcs1_mcs_mat1_6_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_8545, new_AGEMA_signal_8544, mcs1_mcs_mat1_6_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_13417, new_AGEMA_signal_13416, mcs1_mcs_mat1_6_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_12201, new_AGEMA_signal_12200, mcs1_mcs_mat1_6_mcs_out[47]}), .b ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_12885, new_AGEMA_signal_12884, mcs1_mcs_mat1_6_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_11245, new_AGEMA_signal_11244, mcs1_mcs_mat1_6_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .c ({new_AGEMA_signal_12201, new_AGEMA_signal_12200, mcs1_mcs_mat1_6_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_7945, new_AGEMA_signal_7944, mcs1_mcs_mat1_6_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_10283, new_AGEMA_signal_10282, mcs1_mcs_mat1_6_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_11245, new_AGEMA_signal_11244, mcs1_mcs_mat1_6_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({new_AGEMA_signal_10283, new_AGEMA_signal_10282, mcs1_mcs_mat1_6_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3005], Fresh[3004], Fresh[3003]}), .c ({new_AGEMA_signal_8545, new_AGEMA_signal_8544, mcs1_mcs_mat1_6_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3008], Fresh[3007], Fresh[3006]}), .c ({new_AGEMA_signal_9383, new_AGEMA_signal_9382, mcs1_mcs_mat1_6_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_11247, new_AGEMA_signal_11246, mcs1_mcs_mat1_6_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_9385, new_AGEMA_signal_9384, mcs1_mcs_mat1_6_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_12203, new_AGEMA_signal_12202, mcs1_mcs_mat1_6_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_10285, new_AGEMA_signal_10284, mcs1_mcs_mat1_6_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8547, new_AGEMA_signal_8546, mcs1_mcs_mat1_6_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_11247, new_AGEMA_signal_11246, mcs1_mcs_mat1_6_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_11249, new_AGEMA_signal_11248, mcs1_mcs_mat1_6_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_10289, new_AGEMA_signal_10288, mcs1_mcs_mat1_6_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_12205, new_AGEMA_signal_12204, mcs1_mcs_mat1_6_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_11251, new_AGEMA_signal_11250, mcs1_mcs_mat1_6_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_7947, new_AGEMA_signal_7946, mcs1_mcs_mat1_6_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_12207, new_AGEMA_signal_12206, mcs1_mcs_mat1_6_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_10285, new_AGEMA_signal_10284, mcs1_mcs_mat1_6_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9387, new_AGEMA_signal_9386, mcs1_mcs_mat1_6_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_11251, new_AGEMA_signal_11250, mcs1_mcs_mat1_6_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_10287, new_AGEMA_signal_10286, mcs1_mcs_mat1_6_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_9387, new_AGEMA_signal_9386, mcs1_mcs_mat1_6_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_11253, new_AGEMA_signal_11252, mcs1_mcs_mat1_6_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3011], Fresh[3010], Fresh[3009]}), .c ({new_AGEMA_signal_10289, new_AGEMA_signal_10288, mcs1_mcs_mat1_6_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3014], Fresh[3013], Fresh[3012]}), .c ({new_AGEMA_signal_8547, new_AGEMA_signal_8546, mcs1_mcs_mat1_6_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3017], Fresh[3016], Fresh[3015]}), .c ({new_AGEMA_signal_9387, new_AGEMA_signal_9386, mcs1_mcs_mat1_6_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_14743, new_AGEMA_signal_14742, mcs1_mcs_mat1_6_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_11255, new_AGEMA_signal_11254, mcs1_mcs_mat1_6_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_15217, new_AGEMA_signal_15216, mcs1_mcs_mat1_6_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_13421, new_AGEMA_signal_13420, mcs1_mcs_mat1_6_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_13419, new_AGEMA_signal_13418, mcs1_mcs_mat1_6_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_13869, new_AGEMA_signal_13868, mcs1_mcs_mat1_6_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({new_AGEMA_signal_14743, new_AGEMA_signal_14742, mcs1_mcs_mat1_6_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_15219, new_AGEMA_signal_15218, mcs1_mcs_mat1_6_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_13871, new_AGEMA_signal_13870, mcs1_mcs_mat1_6_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_14297, new_AGEMA_signal_14296, mcs1_mcs_mat1_6_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_14743, new_AGEMA_signal_14742, mcs1_mcs_mat1_6_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_13873, new_AGEMA_signal_13872, mcs1_mcs_mat1_6_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_13423, new_AGEMA_signal_13422, mcs1_mcs_mat1_6_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_14297, new_AGEMA_signal_14296, mcs1_mcs_mat1_6_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_13873, new_AGEMA_signal_13872, mcs1_mcs_mat1_6_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_13421, new_AGEMA_signal_13420, mcs1_mcs_mat1_6_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_14299, new_AGEMA_signal_14298, mcs1_mcs_mat1_6_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_12887, new_AGEMA_signal_12886, mcs1_mcs_mat1_6_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_13421, new_AGEMA_signal_13420, mcs1_mcs_mat1_6_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({new_AGEMA_signal_12209, new_AGEMA_signal_12208, mcs1_mcs_mat1_6_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_12887, new_AGEMA_signal_12886, mcs1_mcs_mat1_6_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3020], Fresh[3019], Fresh[3018]}), .c ({new_AGEMA_signal_13873, new_AGEMA_signal_13872, mcs1_mcs_mat1_6_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3023], Fresh[3022], Fresh[3021]}), .c ({new_AGEMA_signal_12209, new_AGEMA_signal_12208, mcs1_mcs_mat1_6_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3026], Fresh[3025], Fresh[3024]}), .c ({new_AGEMA_signal_13423, new_AGEMA_signal_13422, mcs1_mcs_mat1_6_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_10291, new_AGEMA_signal_10290, mcs1_mcs_mat1_6_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_9389, new_AGEMA_signal_9388, mcs1_mcs_mat1_6_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_11257, new_AGEMA_signal_11256, mcs1_mcs_mat1_6_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_8549, new_AGEMA_signal_8548, mcs1_mcs_mat1_6_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_8809, new_AGEMA_signal_8808, mcs1_mcs_mat1_6_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_12889, new_AGEMA_signal_12888, mcs1_mcs_mat1_6_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_10293, new_AGEMA_signal_10292, mcs1_mcs_mat1_6_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_13425, new_AGEMA_signal_13424, mcs1_mcs_mat1_6_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3029], Fresh[3028], Fresh[3027]}), .c ({new_AGEMA_signal_10293, new_AGEMA_signal_10292, mcs1_mcs_mat1_6_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({new_AGEMA_signal_8549, new_AGEMA_signal_8548, mcs1_mcs_mat1_6_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3035], Fresh[3034], Fresh[3033]}), .c ({new_AGEMA_signal_9389, new_AGEMA_signal_9388, mcs1_mcs_mat1_6_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_12213, new_AGEMA_signal_12212, mcs1_mcs_mat1_6_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_11261, new_AGEMA_signal_11260, mcs1_mcs_mat1_6_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_12891, new_AGEMA_signal_12890, mcs1_mcs_mat1_6_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, mcs1_mcs_mat1_6_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_11263, new_AGEMA_signal_11262, mcs1_mcs_mat1_6_mcs_out[29]}), .c ({new_AGEMA_signal_12213, new_AGEMA_signal_12212, mcs1_mcs_mat1_6_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_8551, new_AGEMA_signal_8550, mcs1_mcs_mat1_6_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_11261, new_AGEMA_signal_11260, mcs1_mcs_mat1_6_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_12215, new_AGEMA_signal_12214, mcs1_mcs_mat1_6_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, mcs1_mcs_mat1_6_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .c ({new_AGEMA_signal_11261, new_AGEMA_signal_11260, mcs1_mcs_mat1_6_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_12217, new_AGEMA_signal_12216, mcs1_mcs_mat1_6_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_10295, new_AGEMA_signal_10294, mcs1_mcs_mat1_6_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_12893, new_AGEMA_signal_12892, mcs1_mcs_mat1_6_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_11265, new_AGEMA_signal_11264, mcs1_mcs_mat1_6_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_10297, new_AGEMA_signal_10296, mcs1_mcs_mat1_6_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_12217, new_AGEMA_signal_12216, mcs1_mcs_mat1_6_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_9391, new_AGEMA_signal_9390, mcs1_mcs_mat1_6_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_10297, new_AGEMA_signal_10296, mcs1_mcs_mat1_6_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, mcs1_mcs_mat1_6_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, mcs1_mcs_mat1_6_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_11265, new_AGEMA_signal_11264, mcs1_mcs_mat1_6_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3038], Fresh[3037], Fresh[3036]}), .c ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, mcs1_mcs_mat1_6_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3041], Fresh[3040], Fresh[3039]}), .c ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, mcs1_mcs_mat1_6_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3044], Fresh[3043], Fresh[3042]}), .c ({new_AGEMA_signal_9391, new_AGEMA_signal_9390, mcs1_mcs_mat1_6_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_10301, new_AGEMA_signal_10300, mcs1_mcs_mat1_6_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_11267, new_AGEMA_signal_11266, mcs1_mcs_mat1_6_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_9393, new_AGEMA_signal_9392, mcs1_mcs_mat1_6_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8555, new_AGEMA_signal_8554, mcs1_mcs_mat1_6_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_10301, new_AGEMA_signal_10300, mcs1_mcs_mat1_6_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_11269, new_AGEMA_signal_11268, mcs1_mcs_mat1_6_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_12219, new_AGEMA_signal_12218, mcs1_mcs_mat1_6_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_10305, new_AGEMA_signal_10304, mcs1_mcs_mat1_6_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_8555, new_AGEMA_signal_8554, mcs1_mcs_mat1_6_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_11269, new_AGEMA_signal_11268, mcs1_mcs_mat1_6_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_12221, new_AGEMA_signal_12220, mcs1_mcs_mat1_6_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .c ({new_AGEMA_signal_12895, new_AGEMA_signal_12894, mcs1_mcs_mat1_6_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_10305, new_AGEMA_signal_10304, mcs1_mcs_mat1_6_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_11271, new_AGEMA_signal_11270, mcs1_mcs_mat1_6_mcs_out[24]}), .c ({new_AGEMA_signal_12221, new_AGEMA_signal_12220, mcs1_mcs_mat1_6_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_10303, new_AGEMA_signal_10302, mcs1_mcs_mat1_6_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .c ({new_AGEMA_signal_11271, new_AGEMA_signal_11270, mcs1_mcs_mat1_6_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_9393, new_AGEMA_signal_9392, mcs1_mcs_mat1_6_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_7953, new_AGEMA_signal_7952, mcs1_mcs_mat1_6_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_10303, new_AGEMA_signal_10302, mcs1_mcs_mat1_6_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3047], Fresh[3046], Fresh[3045]}), .c ({new_AGEMA_signal_10305, new_AGEMA_signal_10304, mcs1_mcs_mat1_6_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3050], Fresh[3049], Fresh[3048]}), .c ({new_AGEMA_signal_8555, new_AGEMA_signal_8554, mcs1_mcs_mat1_6_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3053], Fresh[3052], Fresh[3051]}), .c ({new_AGEMA_signal_9393, new_AGEMA_signal_9392, mcs1_mcs_mat1_6_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_13875, new_AGEMA_signal_13874, mcs1_mcs_mat1_6_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .c ({new_AGEMA_signal_14301, new_AGEMA_signal_14300, mcs1_mcs_mat1_6_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_13427, new_AGEMA_signal_13426, mcs1_mcs_mat1_6_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_12223, new_AGEMA_signal_12222, mcs1_mcs_mat1_6_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_13875, new_AGEMA_signal_13874, mcs1_mcs_mat1_6_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_14303, new_AGEMA_signal_14302, mcs1_mcs_mat1_6_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .c ({new_AGEMA_signal_14745, new_AGEMA_signal_14744, mcs1_mcs_mat1_6_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_13879, new_AGEMA_signal_13878, mcs1_mcs_mat1_6_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_12223, new_AGEMA_signal_12222, mcs1_mcs_mat1_6_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_14303, new_AGEMA_signal_14302, mcs1_mcs_mat1_6_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_14747, new_AGEMA_signal_14746, mcs1_mcs_mat1_6_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_15221, new_AGEMA_signal_15220, mcs1_mcs_mat1_6_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_13879, new_AGEMA_signal_13878, mcs1_mcs_mat1_6_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_14305, new_AGEMA_signal_14304, mcs1_mcs_mat1_6_mcs_out[20]}), .c ({new_AGEMA_signal_14747, new_AGEMA_signal_14746, mcs1_mcs_mat1_6_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_13877, new_AGEMA_signal_13876, mcs1_mcs_mat1_6_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_14305, new_AGEMA_signal_14304, mcs1_mcs_mat1_6_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_13427, new_AGEMA_signal_13426, mcs1_mcs_mat1_6_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_11273, new_AGEMA_signal_11272, mcs1_mcs_mat1_6_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_13877, new_AGEMA_signal_13876, mcs1_mcs_mat1_6_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3056], Fresh[3055], Fresh[3054]}), .c ({new_AGEMA_signal_13879, new_AGEMA_signal_13878, mcs1_mcs_mat1_6_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3059], Fresh[3058], Fresh[3057]}), .c ({new_AGEMA_signal_12223, new_AGEMA_signal_12222, mcs1_mcs_mat1_6_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({new_AGEMA_signal_13427, new_AGEMA_signal_13426, mcs1_mcs_mat1_6_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_10307, new_AGEMA_signal_10306, mcs1_mcs_mat1_6_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_10313, new_AGEMA_signal_10312, mcs1_mcs_mat1_6_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_11275, new_AGEMA_signal_11274, mcs1_mcs_mat1_6_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_11277, new_AGEMA_signal_11276, mcs1_mcs_mat1_6_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_7955, new_AGEMA_signal_7954, mcs1_mcs_mat1_6_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, mcs1_mcs_mat1_6_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_12227, new_AGEMA_signal_12226, mcs1_mcs_mat1_6_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_8557, new_AGEMA_signal_8556, mcs1_mcs_mat1_6_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_12897, new_AGEMA_signal_12896, mcs1_mcs_mat1_6_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_7523, new_AGEMA_signal_7522, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_11277, new_AGEMA_signal_11276, mcs1_mcs_mat1_6_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_12227, new_AGEMA_signal_12226, mcs1_mcs_mat1_6_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_10309, new_AGEMA_signal_10308, mcs1_mcs_mat1_6_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .c ({new_AGEMA_signal_11277, new_AGEMA_signal_11276, mcs1_mcs_mat1_6_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_9395, new_AGEMA_signal_9394, mcs1_mcs_mat1_6_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_9397, new_AGEMA_signal_9396, mcs1_mcs_mat1_6_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_10309, new_AGEMA_signal_10308, mcs1_mcs_mat1_6_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_10311, new_AGEMA_signal_10310, mcs1_mcs_mat1_6_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_8557, new_AGEMA_signal_8556, mcs1_mcs_mat1_6_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_11279, new_AGEMA_signal_11278, mcs1_mcs_mat1_6_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3065], Fresh[3064], Fresh[3063]}), .c ({new_AGEMA_signal_10313, new_AGEMA_signal_10312, mcs1_mcs_mat1_6_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3068], Fresh[3067], Fresh[3066]}), .c ({new_AGEMA_signal_8557, new_AGEMA_signal_8556, mcs1_mcs_mat1_6_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3071], Fresh[3070], Fresh[3069]}), .c ({new_AGEMA_signal_9397, new_AGEMA_signal_9396, mcs1_mcs_mat1_6_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_12233, new_AGEMA_signal_12232, mcs1_mcs_mat1_6_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, mcs1_mcs_mat1_6_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_12899, new_AGEMA_signal_12898, mcs1_mcs_mat1_6_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_11285, new_AGEMA_signal_11284, mcs1_mcs_mat1_6_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_11281, new_AGEMA_signal_11280, mcs1_mcs_mat1_6_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_12229, new_AGEMA_signal_12228, mcs1_mcs_mat1_6_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_10317, new_AGEMA_signal_10316, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_8559, new_AGEMA_signal_8558, mcs1_mcs_mat1_6_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_11281, new_AGEMA_signal_11280, mcs1_mcs_mat1_6_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, mcs1_mcs_mat1_6_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_11283, new_AGEMA_signal_11282, mcs1_mcs_mat1_6_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_12231, new_AGEMA_signal_12230, mcs1_mcs_mat1_6_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_10315, new_AGEMA_signal_10314, mcs1_mcs_mat1_6_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_10317, new_AGEMA_signal_10316, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_11283, new_AGEMA_signal_11282, mcs1_mcs_mat1_6_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_7957, new_AGEMA_signal_7956, mcs1_mcs_mat1_6_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_8559, new_AGEMA_signal_8558, mcs1_mcs_mat1_6_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, mcs1_mcs_mat1_6_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_12901, new_AGEMA_signal_12900, mcs1_mcs_mat1_6_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_13429, new_AGEMA_signal_13428, mcs1_mcs_mat1_6_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_12233, new_AGEMA_signal_12232, mcs1_mcs_mat1_6_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_10317, new_AGEMA_signal_10316, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_12901, new_AGEMA_signal_12900, mcs1_mcs_mat1_6_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_11285, new_AGEMA_signal_11284, mcs1_mcs_mat1_6_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_12233, new_AGEMA_signal_12232, mcs1_mcs_mat1_6_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_10315, new_AGEMA_signal_10314, mcs1_mcs_mat1_6_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_11285, new_AGEMA_signal_11284, mcs1_mcs_mat1_6_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_7487, new_AGEMA_signal_7486, shiftr_out[100]}), .b ({new_AGEMA_signal_9399, new_AGEMA_signal_9398, mcs1_mcs_mat1_6_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_10315, new_AGEMA_signal_10314, mcs1_mcs_mat1_6_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3074], Fresh[3073], Fresh[3072]}), .c ({new_AGEMA_signal_10317, new_AGEMA_signal_10316, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3077], Fresh[3076], Fresh[3075]}), .c ({new_AGEMA_signal_8559, new_AGEMA_signal_8558, mcs1_mcs_mat1_6_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3080], Fresh[3079], Fresh[3078]}), .c ({new_AGEMA_signal_9399, new_AGEMA_signal_9398, mcs1_mcs_mat1_6_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_8813, new_AGEMA_signal_8812, mcs1_mcs_mat1_6_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .c ({new_AGEMA_signal_9401, new_AGEMA_signal_9400, mcs1_mcs_mat1_6_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_11289, new_AGEMA_signal_11288, mcs1_mcs_mat1_6_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_12235, new_AGEMA_signal_12234, mcs1_mcs_mat1_6_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_10319, new_AGEMA_signal_10318, mcs1_mcs_mat1_6_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_11287, new_AGEMA_signal_11286, mcs1_mcs_mat1_6_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_9403, new_AGEMA_signal_9402, mcs1_mcs_mat1_6_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_8813, new_AGEMA_signal_8812, mcs1_mcs_mat1_6_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_10319, new_AGEMA_signal_10318, mcs1_mcs_mat1_6_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_7959, new_AGEMA_signal_7958, mcs1_mcs_mat1_6_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_8561, new_AGEMA_signal_8560, mcs1_mcs_mat1_6_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_8813, new_AGEMA_signal_8812, mcs1_mcs_mat1_6_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_12237, new_AGEMA_signal_12236, mcs1_mcs_mat1_6_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, shiftr_out[68]}), .c ({new_AGEMA_signal_12903, new_AGEMA_signal_12902, mcs1_mcs_mat1_6_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_7959, new_AGEMA_signal_7958, mcs1_mcs_mat1_6_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_11289, new_AGEMA_signal_11288, mcs1_mcs_mat1_6_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_12237, new_AGEMA_signal_12236, mcs1_mcs_mat1_6_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_10321, new_AGEMA_signal_10320, mcs1_mcs_mat1_6_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_9403, new_AGEMA_signal_9402, mcs1_mcs_mat1_6_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_11289, new_AGEMA_signal_11288, mcs1_mcs_mat1_6_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3083], Fresh[3082], Fresh[3081]}), .c ({new_AGEMA_signal_10321, new_AGEMA_signal_10320, mcs1_mcs_mat1_6_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3086], Fresh[3085], Fresh[3084]}), .c ({new_AGEMA_signal_8561, new_AGEMA_signal_8560, mcs1_mcs_mat1_6_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, shiftr_out[71]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3089], Fresh[3088], Fresh[3087]}), .c ({new_AGEMA_signal_9403, new_AGEMA_signal_9402, mcs1_mcs_mat1_6_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_15725, new_AGEMA_signal_15724, mcs1_mcs_mat1_6_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_13433, new_AGEMA_signal_13432, mcs1_mcs_mat1_6_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_16129, new_AGEMA_signal_16128, mcs1_mcs_mat1_6_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_15223, new_AGEMA_signal_15222, mcs1_mcs_mat1_6_mcs_out[7]}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .c ({new_AGEMA_signal_15725, new_AGEMA_signal_15724, mcs1_mcs_mat1_6_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_14749, new_AGEMA_signal_14748, mcs1_mcs_mat1_6_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .c ({new_AGEMA_signal_15223, new_AGEMA_signal_15222, mcs1_mcs_mat1_6_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_14307, new_AGEMA_signal_14306, mcs1_mcs_mat1_6_mcs_out[6]}), .b ({new_AGEMA_signal_12241, new_AGEMA_signal_12240, mcs1_mcs_mat1_6_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_14749, new_AGEMA_signal_14748, mcs1_mcs_mat1_6_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_12239, new_AGEMA_signal_12238, mcs1_mcs_mat1_6_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_13881, new_AGEMA_signal_13880, mcs1_mcs_mat1_6_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_14307, new_AGEMA_signal_14306, mcs1_mcs_mat1_6_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12989, new_AGEMA_signal_12988, shiftr_out[37]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({new_AGEMA_signal_13881, new_AGEMA_signal_13880, mcs1_mcs_mat1_6_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, shiftr_out[38]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3095], Fresh[3094], Fresh[3093]}), .c ({new_AGEMA_signal_12241, new_AGEMA_signal_12240, mcs1_mcs_mat1_6_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3098], Fresh[3097], Fresh[3096]}), .c ({new_AGEMA_signal_13433, new_AGEMA_signal_13432, mcs1_mcs_mat1_6_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_9405, new_AGEMA_signal_9404, mcs1_mcs_mat1_6_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_10323, new_AGEMA_signal_10322, mcs1_mcs_mat1_6_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_11295, new_AGEMA_signal_11294, mcs1_mcs_mat1_6_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .b ({new_AGEMA_signal_9407, new_AGEMA_signal_9406, mcs1_mcs_mat1_6_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_10323, new_AGEMA_signal_10322, mcs1_mcs_mat1_6_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_11297, new_AGEMA_signal_11296, mcs1_mcs_mat1_6_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_8563, new_AGEMA_signal_8562, mcs1_mcs_mat1_6_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_12243, new_AGEMA_signal_12242, mcs1_mcs_mat1_6_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_11299, new_AGEMA_signal_11298, mcs1_mcs_mat1_6_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_10327, new_AGEMA_signal_10326, mcs1_mcs_mat1_6_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_12245, new_AGEMA_signal_12244, mcs1_mcs_mat1_6_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_10329, new_AGEMA_signal_10328, mcs1_mcs_mat1_6_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_7961, new_AGEMA_signal_7960, mcs1_mcs_mat1_6_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_11299, new_AGEMA_signal_11298, mcs1_mcs_mat1_6_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, shiftr_out[5]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3101], Fresh[3100], Fresh[3099]}), .c ({new_AGEMA_signal_10329, new_AGEMA_signal_10328, mcs1_mcs_mat1_6_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, shiftr_out[6]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3104], Fresh[3103], Fresh[3102]}), .c ({new_AGEMA_signal_8563, new_AGEMA_signal_8562, mcs1_mcs_mat1_6_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3107], Fresh[3106], Fresh[3105]}), .c ({new_AGEMA_signal_9407, new_AGEMA_signal_9406, mcs1_mcs_mat1_6_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U96 ( .a ({new_AGEMA_signal_13435, new_AGEMA_signal_13434, mcs1_mcs_mat1_7_n128}), .b ({new_AGEMA_signal_15225, new_AGEMA_signal_15224, mcs1_mcs_mat1_7_n127}), .c ({temp_next_s2[65], temp_next_s1[65], temp_next_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U95 ( .a ({new_AGEMA_signal_14795, new_AGEMA_signal_14794, mcs1_mcs_mat1_7_mcs_out[41]}), .b ({new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[45]}), .c ({new_AGEMA_signal_15225, new_AGEMA_signal_15224, mcs1_mcs_mat1_7_n127}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U94 ( .a ({new_AGEMA_signal_8817, new_AGEMA_signal_8816, mcs1_mcs_mat1_7_mcs_out[33]}), .b ({new_AGEMA_signal_12957, new_AGEMA_signal_12956, mcs1_mcs_mat1_7_mcs_out[37]}), .c ({new_AGEMA_signal_13435, new_AGEMA_signal_13434, mcs1_mcs_mat1_7_n128}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U93 ( .a ({new_AGEMA_signal_13883, new_AGEMA_signal_13882, mcs1_mcs_mat1_7_n126}), .b ({new_AGEMA_signal_14751, new_AGEMA_signal_14750, mcs1_mcs_mat1_7_n125}), .c ({temp_next_s2[64], temp_next_s1[64], temp_next_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U92 ( .a ({new_AGEMA_signal_14349, new_AGEMA_signal_14348, mcs1_mcs_mat1_7_mcs_out[40]}), .b ({new_AGEMA_signal_13487, new_AGEMA_signal_13486, mcs1_mcs_mat1_7_mcs_out[44]}), .c ({new_AGEMA_signal_14751, new_AGEMA_signal_14750, mcs1_mcs_mat1_7_n125}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U91 ( .a ({new_AGEMA_signal_13493, new_AGEMA_signal_13492, mcs1_mcs_mat1_7_mcs_out[32]}), .b ({new_AGEMA_signal_11369, new_AGEMA_signal_11368, mcs1_mcs_mat1_7_mcs_out[36]}), .c ({new_AGEMA_signal_13883, new_AGEMA_signal_13882, mcs1_mcs_mat1_7_n126}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U90 ( .a ({new_AGEMA_signal_12247, new_AGEMA_signal_12246, mcs1_mcs_mat1_7_n124}), .b ({new_AGEMA_signal_14753, new_AGEMA_signal_14752, mcs1_mcs_mat1_7_n123}), .c ({temp_next_s2[35], temp_next_s1[35], temp_next_s0[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U89 ( .a ({new_AGEMA_signal_14351, new_AGEMA_signal_14350, mcs1_mcs_mat1_7_mcs_out[27]}), .b ({new_AGEMA_signal_12961, new_AGEMA_signal_12960, mcs1_mcs_mat1_7_mcs_out[31]}), .c ({new_AGEMA_signal_14753, new_AGEMA_signal_14752, mcs1_mcs_mat1_7_n123}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U88 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, mcs1_mcs_mat1_7_mcs_out[19]}), .b ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, mcs1_mcs_mat1_7_mcs_out[23]}), .c ({new_AGEMA_signal_12247, new_AGEMA_signal_12246, mcs1_mcs_mat1_7_n124}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U87 ( .a ({new_AGEMA_signal_12905, new_AGEMA_signal_12904, mcs1_mcs_mat1_7_n122}), .b ({new_AGEMA_signal_15231, new_AGEMA_signal_15230, mcs1_mcs_mat1_7_n121}), .c ({temp_next_s2[34], temp_next_s1[34], temp_next_s0[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U86 ( .a ({new_AGEMA_signal_14797, new_AGEMA_signal_14796, mcs1_mcs_mat1_7_mcs_out[26]}), .b ({new_AGEMA_signal_12337, new_AGEMA_signal_12336, mcs1_mcs_mat1_7_mcs_out[30]}), .c ({new_AGEMA_signal_15231, new_AGEMA_signal_15230, mcs1_mcs_mat1_7_n121}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U85 ( .a ({new_AGEMA_signal_12347, new_AGEMA_signal_12346, mcs1_mcs_mat1_7_mcs_out[18]}), .b ({new_AGEMA_signal_12343, new_AGEMA_signal_12342, mcs1_mcs_mat1_7_mcs_out[22]}), .c ({new_AGEMA_signal_12905, new_AGEMA_signal_12904, mcs1_mcs_mat1_7_n122}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U84 ( .a ({new_AGEMA_signal_13437, new_AGEMA_signal_13436, mcs1_mcs_mat1_7_n120}), .b ({new_AGEMA_signal_15731, new_AGEMA_signal_15730, mcs1_mcs_mat1_7_n119}), .c ({temp_next_s2[33], temp_next_s1[33], temp_next_s0[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U83 ( .a ({new_AGEMA_signal_15269, new_AGEMA_signal_15268, mcs1_mcs_mat1_7_mcs_out[25]}), .b ({new_AGEMA_signal_11377, new_AGEMA_signal_11376, mcs1_mcs_mat1_7_mcs_out[29]}), .c ({new_AGEMA_signal_15731, new_AGEMA_signal_15730, mcs1_mcs_mat1_7_n119}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U82 ( .a ({new_AGEMA_signal_12967, new_AGEMA_signal_12966, mcs1_mcs_mat1_7_mcs_out[17]}), .b ({new_AGEMA_signal_12965, new_AGEMA_signal_12964, mcs1_mcs_mat1_7_mcs_out[21]}), .c ({new_AGEMA_signal_13437, new_AGEMA_signal_13436, mcs1_mcs_mat1_7_n120}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U81 ( .a ({new_AGEMA_signal_12249, new_AGEMA_signal_12248, mcs1_mcs_mat1_7_n118}), .b ({new_AGEMA_signal_14755, new_AGEMA_signal_14754, mcs1_mcs_mat1_7_n117}), .c ({temp_next_s2[32], temp_next_s1[32], temp_next_s0[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U80 ( .a ({new_AGEMA_signal_14355, new_AGEMA_signal_14354, mcs1_mcs_mat1_7_mcs_out[24]}), .b ({new_AGEMA_signal_12963, new_AGEMA_signal_12962, mcs1_mcs_mat1_7_mcs_out[28]}), .c ({new_AGEMA_signal_14755, new_AGEMA_signal_14754, mcs1_mcs_mat1_7_n117}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U79 ( .a ({new_AGEMA_signal_11393, new_AGEMA_signal_11392, mcs1_mcs_mat1_7_mcs_out[16]}), .b ({new_AGEMA_signal_11387, new_AGEMA_signal_11386, mcs1_mcs_mat1_7_mcs_out[20]}), .c ({new_AGEMA_signal_12249, new_AGEMA_signal_12248, mcs1_mcs_mat1_7_n118}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U78 ( .a ({new_AGEMA_signal_13885, new_AGEMA_signal_13884, mcs1_mcs_mat1_7_n116}), .b ({new_AGEMA_signal_13439, new_AGEMA_signal_13438, mcs1_mcs_mat1_7_n115}), .c ({temp_next_s2[3], temp_next_s1[3], temp_next_s0[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U77 ( .a ({new_AGEMA_signal_11405, new_AGEMA_signal_11404, mcs1_mcs_mat1_7_mcs_out[3]}), .b ({new_AGEMA_signal_12975, new_AGEMA_signal_12974, mcs1_mcs_mat1_7_mcs_out[7]}), .c ({new_AGEMA_signal_13439, new_AGEMA_signal_13438, mcs1_mcs_mat1_7_n115}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U76 ( .a ({new_AGEMA_signal_13499, new_AGEMA_signal_13498, mcs1_mcs_mat1_7_mcs_out[11]}), .b ({new_AGEMA_signal_12969, new_AGEMA_signal_12968, mcs1_mcs_mat1_7_mcs_out[15]}), .c ({new_AGEMA_signal_13885, new_AGEMA_signal_13884, mcs1_mcs_mat1_7_n116}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U75 ( .a ({new_AGEMA_signal_13441, new_AGEMA_signal_13440, mcs1_mcs_mat1_7_n114}), .b ({new_AGEMA_signal_15733, new_AGEMA_signal_15732, mcs1_mcs_mat1_7_n113}), .c ({new_AGEMA_signal_16133, new_AGEMA_signal_16132, mcs_out[227]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U74 ( .a ({new_AGEMA_signal_15259, new_AGEMA_signal_15258, mcs1_mcs_mat1_7_mcs_out[123]}), .b ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_15733, new_AGEMA_signal_15732, mcs1_mcs_mat1_7_n113}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U73 ( .a ({new_AGEMA_signal_12271, new_AGEMA_signal_12270, mcs1_mcs_mat1_7_mcs_out[115]}), .b ({new_AGEMA_signal_12917, new_AGEMA_signal_12916, mcs1_mcs_mat1_7_mcs_out[119]}), .c ({new_AGEMA_signal_13441, new_AGEMA_signal_13440, mcs1_mcs_mat1_7_n114}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U72 ( .a ({new_AGEMA_signal_13443, new_AGEMA_signal_13442, mcs1_mcs_mat1_7_n112}), .b ({new_AGEMA_signal_14311, new_AGEMA_signal_14310, mcs1_mcs_mat1_7_n111}), .c ({new_AGEMA_signal_14757, new_AGEMA_signal_14756, mcs_out[226]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U71 ( .a ({new_AGEMA_signal_13899, new_AGEMA_signal_13898, mcs1_mcs_mat1_7_mcs_out[122]}), .b ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_14311, new_AGEMA_signal_14310, mcs1_mcs_mat1_7_n111}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U70 ( .a ({new_AGEMA_signal_11307, new_AGEMA_signal_11306, mcs1_mcs_mat1_7_mcs_out[114]}), .b ({new_AGEMA_signal_12919, new_AGEMA_signal_12918, mcs1_mcs_mat1_7_mcs_out[118]}), .c ({new_AGEMA_signal_13443, new_AGEMA_signal_13442, mcs1_mcs_mat1_7_n112}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U69 ( .a ({new_AGEMA_signal_15235, new_AGEMA_signal_15234, mcs1_mcs_mat1_7_n110}), .b ({new_AGEMA_signal_12251, new_AGEMA_signal_12250, mcs1_mcs_mat1_7_n109}), .c ({temp_next_s2[2], temp_next_s1[2], temp_next_s0[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U68 ( .a ({new_AGEMA_signal_11407, new_AGEMA_signal_11406, mcs1_mcs_mat1_7_mcs_out[2]}), .b ({new_AGEMA_signal_11403, new_AGEMA_signal_11402, mcs1_mcs_mat1_7_mcs_out[6]}), .c ({new_AGEMA_signal_12251, new_AGEMA_signal_12250, mcs1_mcs_mat1_7_n109}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U67 ( .a ({new_AGEMA_signal_14801, new_AGEMA_signal_14800, mcs1_mcs_mat1_7_mcs_out[10]}), .b ({new_AGEMA_signal_12351, new_AGEMA_signal_12350, mcs1_mcs_mat1_7_mcs_out[14]}), .c ({new_AGEMA_signal_15235, new_AGEMA_signal_15234, mcs1_mcs_mat1_7_n110}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U66 ( .a ({new_AGEMA_signal_12907, new_AGEMA_signal_12906, mcs1_mcs_mat1_7_n108}), .b ({new_AGEMA_signal_15737, new_AGEMA_signal_15736, mcs1_mcs_mat1_7_n107}), .c ({new_AGEMA_signal_16135, new_AGEMA_signal_16134, mcs_out[225]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U65 ( .a ({new_AGEMA_signal_15261, new_AGEMA_signal_15260, mcs1_mcs_mat1_7_mcs_out[121]}), .b ({new_AGEMA_signal_9409, new_AGEMA_signal_9408, mcs1_mcs_mat1_7_mcs_out[125]}), .c ({new_AGEMA_signal_15737, new_AGEMA_signal_15736, mcs1_mcs_mat1_7_n107}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U64 ( .a ({new_AGEMA_signal_10337, new_AGEMA_signal_10336, mcs1_mcs_mat1_7_mcs_out[113]}), .b ({new_AGEMA_signal_12269, new_AGEMA_signal_12268, mcs1_mcs_mat1_7_mcs_out[117]}), .c ({new_AGEMA_signal_12907, new_AGEMA_signal_12906, mcs1_mcs_mat1_7_n108}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U63 ( .a ({new_AGEMA_signal_13445, new_AGEMA_signal_13444, mcs1_mcs_mat1_7_n106}), .b ({new_AGEMA_signal_15237, new_AGEMA_signal_15236, mcs1_mcs_mat1_7_n105}), .c ({new_AGEMA_signal_15739, new_AGEMA_signal_15738, mcs_out[224]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U62 ( .a ({new_AGEMA_signal_14775, new_AGEMA_signal_14774, mcs1_mcs_mat1_7_mcs_out[120]}), .b ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_15237, new_AGEMA_signal_15236, mcs1_mcs_mat1_7_n105}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U61 ( .a ({new_AGEMA_signal_12921, new_AGEMA_signal_12920, mcs1_mcs_mat1_7_mcs_out[112]}), .b ({new_AGEMA_signal_11305, new_AGEMA_signal_11304, mcs1_mcs_mat1_7_mcs_out[116]}), .c ({new_AGEMA_signal_13445, new_AGEMA_signal_13444, mcs1_mcs_mat1_7_n106}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U60 ( .a ({new_AGEMA_signal_15239, new_AGEMA_signal_15238, mcs1_mcs_mat1_7_n104}), .b ({new_AGEMA_signal_13447, new_AGEMA_signal_13446, mcs1_mcs_mat1_7_n103}), .c ({new_AGEMA_signal_15741, new_AGEMA_signal_15740, mcs_out[195]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U59 ( .a ({new_AGEMA_signal_12923, new_AGEMA_signal_12922, mcs1_mcs_mat1_7_mcs_out[111]}), .b ({new_AGEMA_signal_12931, new_AGEMA_signal_12930, mcs1_mcs_mat1_7_mcs_out[99]}), .c ({new_AGEMA_signal_13447, new_AGEMA_signal_13446, mcs1_mcs_mat1_7_n103}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U58 ( .a ({new_AGEMA_signal_12281, new_AGEMA_signal_12280, mcs1_mcs_mat1_7_mcs_out[103]}), .b ({new_AGEMA_signal_14777, new_AGEMA_signal_14776, mcs1_mcs_mat1_7_mcs_out[107]}), .c ({new_AGEMA_signal_15239, new_AGEMA_signal_15238, mcs1_mcs_mat1_7_n104}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U57 ( .a ({new_AGEMA_signal_15241, new_AGEMA_signal_15240, mcs1_mcs_mat1_7_n102}), .b ({new_AGEMA_signal_13449, new_AGEMA_signal_13448, mcs1_mcs_mat1_7_n101}), .c ({new_AGEMA_signal_15743, new_AGEMA_signal_15742, mcs_out[194]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U56 ( .a ({new_AGEMA_signal_12925, new_AGEMA_signal_12924, mcs1_mcs_mat1_7_mcs_out[110]}), .b ({new_AGEMA_signal_11325, new_AGEMA_signal_11324, mcs1_mcs_mat1_7_mcs_out[98]}), .c ({new_AGEMA_signal_13449, new_AGEMA_signal_13448, mcs1_mcs_mat1_7_n101}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U55 ( .a ({new_AGEMA_signal_10347, new_AGEMA_signal_10346, mcs1_mcs_mat1_7_mcs_out[102]}), .b ({new_AGEMA_signal_14779, new_AGEMA_signal_14778, mcs1_mcs_mat1_7_mcs_out[106]}), .c ({new_AGEMA_signal_15241, new_AGEMA_signal_15240, mcs1_mcs_mat1_7_n102}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U54 ( .a ({new_AGEMA_signal_15243, new_AGEMA_signal_15242, mcs1_mcs_mat1_7_n100}), .b ({new_AGEMA_signal_13451, new_AGEMA_signal_13450, mcs1_mcs_mat1_7_n99}), .c ({new_AGEMA_signal_15745, new_AGEMA_signal_15744, mcs_out[193]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U53 ( .a ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, mcs1_mcs_mat1_7_mcs_out[109]}), .b ({new_AGEMA_signal_9427, new_AGEMA_signal_9426, mcs1_mcs_mat1_7_mcs_out[97]}), .c ({new_AGEMA_signal_13451, new_AGEMA_signal_13450, mcs1_mcs_mat1_7_n99}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U52 ( .a ({new_AGEMA_signal_11321, new_AGEMA_signal_11320, mcs1_mcs_mat1_7_mcs_out[101]}), .b ({new_AGEMA_signal_14781, new_AGEMA_signal_14780, mcs1_mcs_mat1_7_mcs_out[105]}), .c ({new_AGEMA_signal_15243, new_AGEMA_signal_15242, mcs1_mcs_mat1_7_n100}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U51 ( .a ({new_AGEMA_signal_15747, new_AGEMA_signal_15746, mcs1_mcs_mat1_7_n98}), .b ({new_AGEMA_signal_14313, new_AGEMA_signal_14312, mcs1_mcs_mat1_7_n97}), .c ({new_AGEMA_signal_16137, new_AGEMA_signal_16136, mcs_out[192]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U50 ( .a ({new_AGEMA_signal_12929, new_AGEMA_signal_12928, mcs1_mcs_mat1_7_mcs_out[108]}), .b ({new_AGEMA_signal_13907, new_AGEMA_signal_13906, mcs1_mcs_mat1_7_mcs_out[96]}), .c ({new_AGEMA_signal_14313, new_AGEMA_signal_14312, mcs1_mcs_mat1_7_n97}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U49 ( .a ({new_AGEMA_signal_12283, new_AGEMA_signal_12282, mcs1_mcs_mat1_7_mcs_out[100]}), .b ({new_AGEMA_signal_15263, new_AGEMA_signal_15262, mcs1_mcs_mat1_7_mcs_out[104]}), .c ({new_AGEMA_signal_15747, new_AGEMA_signal_15746, mcs1_mcs_mat1_7_n98}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U48 ( .a ({new_AGEMA_signal_12253, new_AGEMA_signal_12252, mcs1_mcs_mat1_7_n96}), .b ({new_AGEMA_signal_13887, new_AGEMA_signal_13886, mcs1_mcs_mat1_7_n95}), .c ({new_AGEMA_signal_14315, new_AGEMA_signal_14314, mcs_out[163]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U47 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_12287, new_AGEMA_signal_12286, mcs1_mcs_mat1_7_mcs_out[95]}), .c ({new_AGEMA_signal_13887, new_AGEMA_signal_13886, mcs1_mcs_mat1_7_n95}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U46 ( .a ({new_AGEMA_signal_11331, new_AGEMA_signal_11330, mcs1_mcs_mat1_7_mcs_out[83]}), .b ({new_AGEMA_signal_10363, new_AGEMA_signal_10362, mcs1_mcs_mat1_7_mcs_out[87]}), .c ({new_AGEMA_signal_12253, new_AGEMA_signal_12252, mcs1_mcs_mat1_7_n96}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U45 ( .a ({new_AGEMA_signal_12255, new_AGEMA_signal_12254, mcs1_mcs_mat1_7_n94}), .b ({new_AGEMA_signal_13889, new_AGEMA_signal_13888, mcs1_mcs_mat1_7_n93}), .c ({new_AGEMA_signal_14317, new_AGEMA_signal_14316, mcs_out[162]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U43 ( .a ({new_AGEMA_signal_11333, new_AGEMA_signal_11332, mcs1_mcs_mat1_7_mcs_out[82]}), .b ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_12255, new_AGEMA_signal_12254, mcs1_mcs_mat1_7_n94}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U42 ( .a ({new_AGEMA_signal_12257, new_AGEMA_signal_12256, mcs1_mcs_mat1_7_n92}), .b ({new_AGEMA_signal_13891, new_AGEMA_signal_13890, mcs1_mcs_mat1_7_n91}), .c ({new_AGEMA_signal_14319, new_AGEMA_signal_14318, mcs_out[161]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U41 ( .a ({new_AGEMA_signal_13479, new_AGEMA_signal_13478, mcs1_mcs_mat1_7_mcs_out[89]}), .b ({new_AGEMA_signal_10359, new_AGEMA_signal_10358, mcs1_mcs_mat1_7_mcs_out[93]}), .c ({new_AGEMA_signal_13891, new_AGEMA_signal_13890, mcs1_mcs_mat1_7_n91}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U40 ( .a ({new_AGEMA_signal_11335, new_AGEMA_signal_11334, mcs1_mcs_mat1_7_mcs_out[81]}), .b ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_12257, new_AGEMA_signal_12256, mcs1_mcs_mat1_7_n92}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U39 ( .a ({new_AGEMA_signal_12909, new_AGEMA_signal_12908, mcs1_mcs_mat1_7_n90}), .b ({new_AGEMA_signal_13453, new_AGEMA_signal_13452, mcs1_mcs_mat1_7_n89}), .c ({new_AGEMA_signal_13893, new_AGEMA_signal_13892, mcs_out[160]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U38 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_12933, new_AGEMA_signal_12932, mcs1_mcs_mat1_7_mcs_out[92]}), .c ({new_AGEMA_signal_13453, new_AGEMA_signal_13452, mcs1_mcs_mat1_7_n89}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U37 ( .a ({new_AGEMA_signal_12291, new_AGEMA_signal_12290, mcs1_mcs_mat1_7_mcs_out[80]}), .b ({new_AGEMA_signal_11329, new_AGEMA_signal_11328, mcs1_mcs_mat1_7_mcs_out[84]}), .c ({new_AGEMA_signal_12909, new_AGEMA_signal_12908, mcs1_mcs_mat1_7_n90}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U36 ( .a ({new_AGEMA_signal_12911, new_AGEMA_signal_12910, mcs1_mcs_mat1_7_n88}), .b ({new_AGEMA_signal_14759, new_AGEMA_signal_14758, mcs1_mcs_mat1_7_n87}), .c ({temp_next_s2[1], temp_next_s1[1], temp_next_s0[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U35 ( .a ({new_AGEMA_signal_9473, new_AGEMA_signal_9472, mcs1_mcs_mat1_7_mcs_out[5]}), .b ({new_AGEMA_signal_14357, new_AGEMA_signal_14356, mcs1_mcs_mat1_7_mcs_out[9]}), .c ({new_AGEMA_signal_14759, new_AGEMA_signal_14758, mcs1_mcs_mat1_7_n87}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U34 ( .a ({new_AGEMA_signal_12353, new_AGEMA_signal_12352, mcs1_mcs_mat1_7_mcs_out[13]}), .b ({new_AGEMA_signal_12361, new_AGEMA_signal_12360, mcs1_mcs_mat1_7_mcs_out[1]}), .c ({new_AGEMA_signal_12911, new_AGEMA_signal_12910, mcs1_mcs_mat1_7_n88}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U33 ( .a ({new_AGEMA_signal_13455, new_AGEMA_signal_13454, mcs1_mcs_mat1_7_n86}), .b ({new_AGEMA_signal_14321, new_AGEMA_signal_14320, mcs1_mcs_mat1_7_n85}), .c ({new_AGEMA_signal_14761, new_AGEMA_signal_14760, mcs_out[131]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U32 ( .a ({new_AGEMA_signal_13909, new_AGEMA_signal_13908, mcs1_mcs_mat1_7_mcs_out[75]}), .b ({new_AGEMA_signal_12293, new_AGEMA_signal_12292, mcs1_mcs_mat1_7_mcs_out[79]}), .c ({new_AGEMA_signal_14321, new_AGEMA_signal_14320, mcs1_mcs_mat1_7_n85}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U31 ( .a ({new_AGEMA_signal_12943, new_AGEMA_signal_12942, mcs1_mcs_mat1_7_mcs_out[67]}), .b ({new_AGEMA_signal_12301, new_AGEMA_signal_12300, mcs1_mcs_mat1_7_mcs_out[71]}), .c ({new_AGEMA_signal_13455, new_AGEMA_signal_13454, mcs1_mcs_mat1_7_n86}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U30 ( .a ({new_AGEMA_signal_13457, new_AGEMA_signal_13456, mcs1_mcs_mat1_7_n84}), .b ({new_AGEMA_signal_15749, new_AGEMA_signal_15748, mcs1_mcs_mat1_7_n83}), .c ({new_AGEMA_signal_16139, new_AGEMA_signal_16138, mcs_out[130]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U29 ( .a ({new_AGEMA_signal_15265, new_AGEMA_signal_15264, mcs1_mcs_mat1_7_mcs_out[74]}), .b ({new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_7_mcs_out[78]}), .c ({new_AGEMA_signal_15749, new_AGEMA_signal_15748, mcs1_mcs_mat1_7_n83}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U28 ( .a ({new_AGEMA_signal_12307, new_AGEMA_signal_12306, mcs1_mcs_mat1_7_mcs_out[66]}), .b ({new_AGEMA_signal_12939, new_AGEMA_signal_12938, mcs1_mcs_mat1_7_mcs_out[70]}), .c ({new_AGEMA_signal_13457, new_AGEMA_signal_13456, mcs1_mcs_mat1_7_n84}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U27 ( .a ({new_AGEMA_signal_13459, new_AGEMA_signal_13458, mcs1_mcs_mat1_7_n82}), .b ({new_AGEMA_signal_14763, new_AGEMA_signal_14762, mcs1_mcs_mat1_7_n81}), .c ({new_AGEMA_signal_15247, new_AGEMA_signal_15246, mcs_out[129]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U26 ( .a ({new_AGEMA_signal_14333, new_AGEMA_signal_14332, mcs1_mcs_mat1_7_mcs_out[73]}), .b ({new_AGEMA_signal_10373, new_AGEMA_signal_10372, mcs1_mcs_mat1_7_mcs_out[77]}), .c ({new_AGEMA_signal_14763, new_AGEMA_signal_14762, mcs1_mcs_mat1_7_n81}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U25 ( .a ({new_AGEMA_signal_10383, new_AGEMA_signal_10382, mcs1_mcs_mat1_7_mcs_out[65]}), .b ({new_AGEMA_signal_12941, new_AGEMA_signal_12940, mcs1_mcs_mat1_7_mcs_out[69]}), .c ({new_AGEMA_signal_13459, new_AGEMA_signal_13458, mcs1_mcs_mat1_7_n82}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U24 ( .a ({new_AGEMA_signal_13895, new_AGEMA_signal_13894, mcs1_mcs_mat1_7_n80}), .b ({new_AGEMA_signal_15751, new_AGEMA_signal_15750, mcs1_mcs_mat1_7_n79}), .c ({new_AGEMA_signal_16141, new_AGEMA_signal_16140, mcs_out[128]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U23 ( .a ({new_AGEMA_signal_15267, new_AGEMA_signal_15266, mcs1_mcs_mat1_7_mcs_out[72]}), .b ({new_AGEMA_signal_12935, new_AGEMA_signal_12934, mcs1_mcs_mat1_7_mcs_out[76]}), .c ({new_AGEMA_signal_15751, new_AGEMA_signal_15750, mcs1_mcs_mat1_7_n79}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U22 ( .a ({new_AGEMA_signal_13483, new_AGEMA_signal_13482, mcs1_mcs_mat1_7_mcs_out[64]}), .b ({new_AGEMA_signal_12305, new_AGEMA_signal_12304, mcs1_mcs_mat1_7_mcs_out[68]}), .c ({new_AGEMA_signal_13895, new_AGEMA_signal_13894, mcs1_mcs_mat1_7_n80}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U21 ( .a ({new_AGEMA_signal_12913, new_AGEMA_signal_12912, mcs1_mcs_mat1_7_n78}), .b ({new_AGEMA_signal_14765, new_AGEMA_signal_14764, mcs1_mcs_mat1_7_n77}), .c ({temp_next_s2[99], temp_next_s1[99], temp_next_s0[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U20 ( .a ({new_AGEMA_signal_14337, new_AGEMA_signal_14336, mcs1_mcs_mat1_7_mcs_out[59]}), .b ({new_AGEMA_signal_12311, new_AGEMA_signal_12310, mcs1_mcs_mat1_7_mcs_out[63]}), .c ({new_AGEMA_signal_14765, new_AGEMA_signal_14764, mcs1_mcs_mat1_7_n77}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U19 ( .a ({new_AGEMA_signal_10399, new_AGEMA_signal_10398, mcs1_mcs_mat1_7_mcs_out[51]}), .b ({new_AGEMA_signal_12321, new_AGEMA_signal_12320, mcs1_mcs_mat1_7_mcs_out[55]}), .c ({new_AGEMA_signal_12913, new_AGEMA_signal_12912, mcs1_mcs_mat1_7_n78}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U18 ( .a ({new_AGEMA_signal_13461, new_AGEMA_signal_13460, mcs1_mcs_mat1_7_n76}), .b ({new_AGEMA_signal_14323, new_AGEMA_signal_14322, mcs1_mcs_mat1_7_n75}), .c ({temp_next_s2[98], temp_next_s1[98], temp_next_s0[98]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U17 ( .a ({new_AGEMA_signal_13915, new_AGEMA_signal_13914, mcs1_mcs_mat1_7_mcs_out[58]}), .b ({new_AGEMA_signal_11349, new_AGEMA_signal_11348, mcs1_mcs_mat1_7_mcs_out[62]}), .c ({new_AGEMA_signal_14323, new_AGEMA_signal_14322, mcs1_mcs_mat1_7_n75}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U16 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_12949, new_AGEMA_signal_12948, mcs1_mcs_mat1_7_mcs_out[54]}), .c ({new_AGEMA_signal_13461, new_AGEMA_signal_13460, mcs1_mcs_mat1_7_n76}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U15 ( .a ({new_AGEMA_signal_13463, new_AGEMA_signal_13462, mcs1_mcs_mat1_7_n74}), .b ({new_AGEMA_signal_14769, new_AGEMA_signal_14768, mcs1_mcs_mat1_7_n73}), .c ({temp_next_s2[97], temp_next_s1[97], temp_next_s0[97]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U14 ( .a ({new_AGEMA_signal_14339, new_AGEMA_signal_14338, mcs1_mcs_mat1_7_mcs_out[57]}), .b ({new_AGEMA_signal_11351, new_AGEMA_signal_11350, mcs1_mcs_mat1_7_mcs_out[61]}), .c ({new_AGEMA_signal_14769, new_AGEMA_signal_14768, mcs1_mcs_mat1_7_n73}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U13 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_12951, new_AGEMA_signal_12950, mcs1_mcs_mat1_7_mcs_out[53]}), .c ({new_AGEMA_signal_13463, new_AGEMA_signal_13462, mcs1_mcs_mat1_7_n74}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U12 ( .a ({new_AGEMA_signal_12915, new_AGEMA_signal_12914, mcs1_mcs_mat1_7_n72}), .b ({new_AGEMA_signal_15253, new_AGEMA_signal_15252, mcs1_mcs_mat1_7_n71}), .c ({temp_next_s2[96], temp_next_s1[96], temp_next_s0[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U11 ( .a ({new_AGEMA_signal_14789, new_AGEMA_signal_14788, mcs1_mcs_mat1_7_mcs_out[56]}), .b ({new_AGEMA_signal_12947, new_AGEMA_signal_12946, mcs1_mcs_mat1_7_mcs_out[60]}), .c ({new_AGEMA_signal_15253, new_AGEMA_signal_15252, mcs1_mcs_mat1_7_n71}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U10 ( .a ({new_AGEMA_signal_11361, new_AGEMA_signal_11360, mcs1_mcs_mat1_7_mcs_out[48]}), .b ({new_AGEMA_signal_12325, new_AGEMA_signal_12324, mcs1_mcs_mat1_7_mcs_out[52]}), .c ({new_AGEMA_signal_12915, new_AGEMA_signal_12914, mcs1_mcs_mat1_7_n72}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U9 ( .a ({new_AGEMA_signal_13465, new_AGEMA_signal_13464, mcs1_mcs_mat1_7_n70}), .b ({new_AGEMA_signal_15255, new_AGEMA_signal_15254, mcs1_mcs_mat1_7_n69}), .c ({temp_next_s2[67], temp_next_s1[67], temp_next_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U8 ( .a ({new_AGEMA_signal_14791, new_AGEMA_signal_14790, mcs1_mcs_mat1_7_mcs_out[43]}), .b ({new_AGEMA_signal_12327, new_AGEMA_signal_12326, mcs1_mcs_mat1_7_mcs_out[47]}), .c ({new_AGEMA_signal_15255, new_AGEMA_signal_15254, mcs1_mcs_mat1_7_n69}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U7 ( .a ({new_AGEMA_signal_12333, new_AGEMA_signal_12332, mcs1_mcs_mat1_7_mcs_out[35]}), .b ({new_AGEMA_signal_12955, new_AGEMA_signal_12954, mcs1_mcs_mat1_7_mcs_out[39]}), .c ({new_AGEMA_signal_13465, new_AGEMA_signal_13464, mcs1_mcs_mat1_7_n70}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U6 ( .a ({new_AGEMA_signal_12259, new_AGEMA_signal_12258, mcs1_mcs_mat1_7_n68}), .b ({new_AGEMA_signal_15257, new_AGEMA_signal_15256, mcs1_mcs_mat1_7_n67}), .c ({temp_next_s2[66], temp_next_s1[66], temp_next_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U5 ( .a ({new_AGEMA_signal_14793, new_AGEMA_signal_14792, mcs1_mcs_mat1_7_mcs_out[42]}), .b ({new_AGEMA_signal_9451, new_AGEMA_signal_9450, mcs1_mcs_mat1_7_mcs_out[46]}), .c ({new_AGEMA_signal_15257, new_AGEMA_signal_15256, mcs1_mcs_mat1_7_n67}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U4 ( .a ({new_AGEMA_signal_11371, new_AGEMA_signal_11370, mcs1_mcs_mat1_7_mcs_out[34]}), .b ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, mcs1_mcs_mat1_7_mcs_out[38]}), .c ({new_AGEMA_signal_12259, new_AGEMA_signal_12258, mcs1_mcs_mat1_7_n68}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U3 ( .a ({new_AGEMA_signal_13897, new_AGEMA_signal_13896, mcs1_mcs_mat1_7_n66}), .b ({new_AGEMA_signal_15759, new_AGEMA_signal_15758, mcs1_mcs_mat1_7_n65}), .c ({temp_next_s2[0], temp_next_s1[0], temp_next_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U2 ( .a ({new_AGEMA_signal_13939, new_AGEMA_signal_13938, mcs1_mcs_mat1_7_mcs_out[4]}), .b ({new_AGEMA_signal_15271, new_AGEMA_signal_15270, mcs1_mcs_mat1_7_mcs_out[8]}), .c ({new_AGEMA_signal_15759, new_AGEMA_signal_15758, mcs1_mcs_mat1_7_n65}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_U1 ( .a ({new_AGEMA_signal_12363, new_AGEMA_signal_12362, mcs1_mcs_mat1_7_mcs_out[0]}), .b ({new_AGEMA_signal_13497, new_AGEMA_signal_13496, mcs1_mcs_mat1_7_mcs_out[12]}), .c ({new_AGEMA_signal_13897, new_AGEMA_signal_13896, mcs1_mcs_mat1_7_n66}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_14771, new_AGEMA_signal_14770, mcs1_mcs_mat1_7_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_15259, new_AGEMA_signal_15258, mcs1_mcs_mat1_7_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_14325, new_AGEMA_signal_14324, mcs1_mcs_mat1_7_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_11301, new_AGEMA_signal_11300, mcs1_mcs_mat1_7_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_14771, new_AGEMA_signal_14770, mcs1_mcs_mat1_7_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_12261, new_AGEMA_signal_12260, mcs1_mcs_mat1_7_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_13467, new_AGEMA_signal_13466, mcs1_mcs_mat1_7_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_13899, new_AGEMA_signal_13898, mcs1_mcs_mat1_7_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_12263, new_AGEMA_signal_12262, mcs1_mcs_mat1_7_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .c ({new_AGEMA_signal_13467, new_AGEMA_signal_13466, mcs1_mcs_mat1_7_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_14773, new_AGEMA_signal_14772, mcs1_mcs_mat1_7_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .c ({new_AGEMA_signal_15261, new_AGEMA_signal_15260, mcs1_mcs_mat1_7_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_14325, new_AGEMA_signal_14324, mcs1_mcs_mat1_7_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_14773, new_AGEMA_signal_14772, mcs1_mcs_mat1_7_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_13901, new_AGEMA_signal_13900, mcs1_mcs_mat1_7_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_13469, new_AGEMA_signal_13468, mcs1_mcs_mat1_7_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_14325, new_AGEMA_signal_14324, mcs1_mcs_mat1_7_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_14327, new_AGEMA_signal_14326, mcs1_mcs_mat1_7_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_14775, new_AGEMA_signal_14774, mcs1_mcs_mat1_7_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_13901, new_AGEMA_signal_13900, mcs1_mcs_mat1_7_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_12263, new_AGEMA_signal_12262, mcs1_mcs_mat1_7_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_14327, new_AGEMA_signal_14326, mcs1_mcs_mat1_7_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3110], Fresh[3109], Fresh[3108]}), .c ({new_AGEMA_signal_13901, new_AGEMA_signal_13900, mcs1_mcs_mat1_7_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3113], Fresh[3112], Fresh[3111]}), .c ({new_AGEMA_signal_12263, new_AGEMA_signal_12262, mcs1_mcs_mat1_7_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3116], Fresh[3115], Fresh[3114]}), .c ({new_AGEMA_signal_13469, new_AGEMA_signal_13468, mcs1_mcs_mat1_7_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_12265, new_AGEMA_signal_12264, mcs1_mcs_mat1_7_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .c ({new_AGEMA_signal_12917, new_AGEMA_signal_12916, mcs1_mcs_mat1_7_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_11303, new_AGEMA_signal_11302, mcs1_mcs_mat1_7_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_9415, new_AGEMA_signal_9414, mcs1_mcs_mat1_7_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_12265, new_AGEMA_signal_12264, mcs1_mcs_mat1_7_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_12267, new_AGEMA_signal_12266, mcs1_mcs_mat1_7_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_10333, new_AGEMA_signal_10332, mcs1_mcs_mat1_7_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_12919, new_AGEMA_signal_12918, mcs1_mcs_mat1_7_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_11303, new_AGEMA_signal_11302, mcs1_mcs_mat1_7_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .c ({new_AGEMA_signal_12267, new_AGEMA_signal_12266, mcs1_mcs_mat1_7_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_11303, new_AGEMA_signal_11302, mcs1_mcs_mat1_7_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10331, new_AGEMA_signal_10330, mcs1_mcs_mat1_7_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_12269, new_AGEMA_signal_12268, mcs1_mcs_mat1_7_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_10335, new_AGEMA_signal_10334, mcs1_mcs_mat1_7_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_11303, new_AGEMA_signal_11302, mcs1_mcs_mat1_7_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_9413, new_AGEMA_signal_9412, mcs1_mcs_mat1_7_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_10333, new_AGEMA_signal_10332, mcs1_mcs_mat1_7_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_11305, new_AGEMA_signal_11304, mcs1_mcs_mat1_7_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_7963, new_AGEMA_signal_7962, mcs1_mcs_mat1_7_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_9415, new_AGEMA_signal_9414, mcs1_mcs_mat1_7_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_10333, new_AGEMA_signal_10332, mcs1_mcs_mat1_7_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_9413, new_AGEMA_signal_9412, mcs1_mcs_mat1_7_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3119], Fresh[3118], Fresh[3117]}), .c ({new_AGEMA_signal_10335, new_AGEMA_signal_10334, mcs1_mcs_mat1_7_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3125], Fresh[3124], Fresh[3123]}), .c ({new_AGEMA_signal_9415, new_AGEMA_signal_9414, mcs1_mcs_mat1_7_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_11309, new_AGEMA_signal_11308, mcs1_mcs_mat1_7_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_8567, new_AGEMA_signal_8566, mcs1_mcs_mat1_7_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_12271, new_AGEMA_signal_12270, mcs1_mcs_mat1_7_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_9417, new_AGEMA_signal_9416, mcs1_mcs_mat1_7_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_9419, new_AGEMA_signal_9418, mcs1_mcs_mat1_7_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_10337, new_AGEMA_signal_10336, mcs1_mcs_mat1_7_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_11311, new_AGEMA_signal_11310, mcs1_mcs_mat1_7_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_12273, new_AGEMA_signal_12272, mcs1_mcs_mat1_7_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_12921, new_AGEMA_signal_12920, mcs1_mcs_mat1_7_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_11309, new_AGEMA_signal_11308, mcs1_mcs_mat1_7_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_12273, new_AGEMA_signal_12272, mcs1_mcs_mat1_7_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_7965, new_AGEMA_signal_7964, mcs1_mcs_mat1_7_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_10341, new_AGEMA_signal_10340, mcs1_mcs_mat1_7_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_11309, new_AGEMA_signal_11308, mcs1_mcs_mat1_7_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, mcs1_mcs_mat1_7_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_10339, new_AGEMA_signal_10338, mcs1_mcs_mat1_7_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_11311, new_AGEMA_signal_11310, mcs1_mcs_mat1_7_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3128], Fresh[3127], Fresh[3126]}), .c ({new_AGEMA_signal_10341, new_AGEMA_signal_10340, mcs1_mcs_mat1_7_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3131], Fresh[3130], Fresh[3129]}), .c ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, mcs1_mcs_mat1_7_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3134], Fresh[3133], Fresh[3132]}), .c ({new_AGEMA_signal_9419, new_AGEMA_signal_9418, mcs1_mcs_mat1_7_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({new_AGEMA_signal_12275, new_AGEMA_signal_12274, mcs1_mcs_mat1_7_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12923, new_AGEMA_signal_12922, mcs1_mcs_mat1_7_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({new_AGEMA_signal_12277, new_AGEMA_signal_12276, mcs1_mcs_mat1_7_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12925, new_AGEMA_signal_12924, mcs1_mcs_mat1_7_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_9421, new_AGEMA_signal_9420, mcs1_mcs_mat1_7_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_12275, new_AGEMA_signal_12274, mcs1_mcs_mat1_7_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, mcs1_mcs_mat1_7_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_7_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_11313, new_AGEMA_signal_11312, mcs1_mcs_mat1_7_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_12275, new_AGEMA_signal_12274, mcs1_mcs_mat1_7_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_10343, new_AGEMA_signal_10342, mcs1_mcs_mat1_7_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_12277, new_AGEMA_signal_12276, mcs1_mcs_mat1_7_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_12929, new_AGEMA_signal_12928, mcs1_mcs_mat1_7_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_11315, new_AGEMA_signal_11314, mcs1_mcs_mat1_7_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_12277, new_AGEMA_signal_12276, mcs1_mcs_mat1_7_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_9421, new_AGEMA_signal_9420, mcs1_mcs_mat1_7_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_10345, new_AGEMA_signal_10344, mcs1_mcs_mat1_7_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_11315, new_AGEMA_signal_11314, mcs1_mcs_mat1_7_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3137], Fresh[3136], Fresh[3135]}), .c ({new_AGEMA_signal_10345, new_AGEMA_signal_10344, mcs1_mcs_mat1_7_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3140], Fresh[3139], Fresh[3138]}), .c ({new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_7_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3143], Fresh[3142], Fresh[3141]}), .c ({new_AGEMA_signal_9421, new_AGEMA_signal_9420, mcs1_mcs_mat1_7_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_14331, new_AGEMA_signal_14330, mcs1_mcs_mat1_7_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_14329, new_AGEMA_signal_14328, mcs1_mcs_mat1_7_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_14777, new_AGEMA_signal_14776, mcs1_mcs_mat1_7_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_14329, new_AGEMA_signal_14328, mcs1_mcs_mat1_7_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_13471, new_AGEMA_signal_13470, mcs1_mcs_mat1_7_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_14779, new_AGEMA_signal_14778, mcs1_mcs_mat1_7_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, mcs1_mcs_mat1_7_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .c ({new_AGEMA_signal_13471, new_AGEMA_signal_13470, mcs1_mcs_mat1_7_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_14329, new_AGEMA_signal_14328, mcs1_mcs_mat1_7_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_14781, new_AGEMA_signal_14780, mcs1_mcs_mat1_7_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_13905, new_AGEMA_signal_13904, mcs1_mcs_mat1_7_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_11317, new_AGEMA_signal_11316, mcs1_mcs_mat1_7_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_14329, new_AGEMA_signal_14328, mcs1_mcs_mat1_7_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_14783, new_AGEMA_signal_14782, mcs1_mcs_mat1_7_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_15263, new_AGEMA_signal_15262, mcs1_mcs_mat1_7_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_14331, new_AGEMA_signal_14330, mcs1_mcs_mat1_7_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_13905, new_AGEMA_signal_13904, mcs1_mcs_mat1_7_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_14783, new_AGEMA_signal_14782, mcs1_mcs_mat1_7_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_13903, new_AGEMA_signal_13902, mcs1_mcs_mat1_7_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .c ({new_AGEMA_signal_14331, new_AGEMA_signal_14330, mcs1_mcs_mat1_7_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, mcs1_mcs_mat1_7_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_13473, new_AGEMA_signal_13472, mcs1_mcs_mat1_7_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_13903, new_AGEMA_signal_13902, mcs1_mcs_mat1_7_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3146], Fresh[3145], Fresh[3144]}), .c ({new_AGEMA_signal_13905, new_AGEMA_signal_13904, mcs1_mcs_mat1_7_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3149], Fresh[3148], Fresh[3147]}), .c ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, mcs1_mcs_mat1_7_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({new_AGEMA_signal_13473, new_AGEMA_signal_13472, mcs1_mcs_mat1_7_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_9423, new_AGEMA_signal_9422, mcs1_mcs_mat1_7_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_11319, new_AGEMA_signal_11318, mcs1_mcs_mat1_7_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_12281, new_AGEMA_signal_12280, mcs1_mcs_mat1_7_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_10353, new_AGEMA_signal_10352, mcs1_mcs_mat1_7_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_11319, new_AGEMA_signal_11318, mcs1_mcs_mat1_7_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_10349, new_AGEMA_signal_10348, mcs1_mcs_mat1_7_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_9425, new_AGEMA_signal_9424, mcs1_mcs_mat1_7_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_11321, new_AGEMA_signal_11320, mcs1_mcs_mat1_7_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_10351, new_AGEMA_signal_10350, mcs1_mcs_mat1_7_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_11323, new_AGEMA_signal_11322, mcs1_mcs_mat1_7_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_12283, new_AGEMA_signal_12282, mcs1_mcs_mat1_7_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_7969, new_AGEMA_signal_7968, mcs1_mcs_mat1_7_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_10353, new_AGEMA_signal_10352, mcs1_mcs_mat1_7_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_11323, new_AGEMA_signal_11322, mcs1_mcs_mat1_7_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_8573, new_AGEMA_signal_8572, mcs1_mcs_mat1_7_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .c ({new_AGEMA_signal_10351, new_AGEMA_signal_10350, mcs1_mcs_mat1_7_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3155], Fresh[3154], Fresh[3153]}), .c ({new_AGEMA_signal_10353, new_AGEMA_signal_10352, mcs1_mcs_mat1_7_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3158], Fresh[3157], Fresh[3156]}), .c ({new_AGEMA_signal_8573, new_AGEMA_signal_8572, mcs1_mcs_mat1_7_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3161], Fresh[3160], Fresh[3159]}), .c ({new_AGEMA_signal_9425, new_AGEMA_signal_9424, mcs1_mcs_mat1_7_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_13475, new_AGEMA_signal_13474, mcs1_mcs_mat1_7_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_9429, new_AGEMA_signal_9428, mcs1_mcs_mat1_7_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_13907, new_AGEMA_signal_13906, mcs1_mcs_mat1_7_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_12931, new_AGEMA_signal_12930, mcs1_mcs_mat1_7_mcs_out[99]}), .b ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .c ({new_AGEMA_signal_13475, new_AGEMA_signal_13474, mcs1_mcs_mat1_7_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_12285, new_AGEMA_signal_12284, mcs1_mcs_mat1_7_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .c ({new_AGEMA_signal_12931, new_AGEMA_signal_12930, mcs1_mcs_mat1_7_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_11325, new_AGEMA_signal_11324, mcs1_mcs_mat1_7_mcs_out[98]}), .b ({new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_7_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_12285, new_AGEMA_signal_12284, mcs1_mcs_mat1_7_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, mcs1_mcs_mat1_7_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_10355, new_AGEMA_signal_10354, mcs1_mcs_mat1_7_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_11325, new_AGEMA_signal_11324, mcs1_mcs_mat1_7_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3164], Fresh[3163], Fresh[3162]}), .c ({new_AGEMA_signal_10355, new_AGEMA_signal_10354, mcs1_mcs_mat1_7_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3167], Fresh[3166], Fresh[3165]}), .c ({new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_7_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3170], Fresh[3169], Fresh[3168]}), .c ({new_AGEMA_signal_9429, new_AGEMA_signal_9428, mcs1_mcs_mat1_7_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_11327, new_AGEMA_signal_11326, mcs1_mcs_mat1_7_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_12287, new_AGEMA_signal_12286, mcs1_mcs_mat1_7_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_9433, new_AGEMA_signal_9432, mcs1_mcs_mat1_7_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_9435, new_AGEMA_signal_9434, mcs1_mcs_mat1_7_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_10359, new_AGEMA_signal_10358, mcs1_mcs_mat1_7_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_12289, new_AGEMA_signal_12288, mcs1_mcs_mat1_7_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_8579, new_AGEMA_signal_8578, mcs1_mcs_mat1_7_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_12933, new_AGEMA_signal_12932, mcs1_mcs_mat1_7_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_11327, new_AGEMA_signal_11326, mcs1_mcs_mat1_7_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_12289, new_AGEMA_signal_12288, mcs1_mcs_mat1_7_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_7973, new_AGEMA_signal_7972, mcs1_mcs_mat1_7_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_10361, new_AGEMA_signal_10360, mcs1_mcs_mat1_7_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_11327, new_AGEMA_signal_11326, mcs1_mcs_mat1_7_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3173], Fresh[3172], Fresh[3171]}), .c ({new_AGEMA_signal_10361, new_AGEMA_signal_10360, mcs1_mcs_mat1_7_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3176], Fresh[3175], Fresh[3174]}), .c ({new_AGEMA_signal_8579, new_AGEMA_signal_8578, mcs1_mcs_mat1_7_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3179], Fresh[3178], Fresh[3177]}), .c ({new_AGEMA_signal_9435, new_AGEMA_signal_9434, mcs1_mcs_mat1_7_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_10369, new_AGEMA_signal_10368, mcs1_mcs_mat1_7_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_10371, new_AGEMA_signal_10370, mcs1_mcs_mat1_7_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_11331, new_AGEMA_signal_11330, mcs1_mcs_mat1_7_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_10365, new_AGEMA_signal_10364, mcs1_mcs_mat1_7_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_7975, new_AGEMA_signal_7974, mcs1_mcs_mat1_7_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_11333, new_AGEMA_signal_11332, mcs1_mcs_mat1_7_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_9437, new_AGEMA_signal_9436, mcs1_mcs_mat1_7_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_10365, new_AGEMA_signal_10364, mcs1_mcs_mat1_7_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_10367, new_AGEMA_signal_10366, mcs1_mcs_mat1_7_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_11335, new_AGEMA_signal_11334, mcs1_mcs_mat1_7_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, mcs1_mcs_mat1_7_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_9437, new_AGEMA_signal_9436, mcs1_mcs_mat1_7_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_10367, new_AGEMA_signal_10366, mcs1_mcs_mat1_7_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_11337, new_AGEMA_signal_11336, mcs1_mcs_mat1_7_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .c ({new_AGEMA_signal_12291, new_AGEMA_signal_12290, mcs1_mcs_mat1_7_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_10369, new_AGEMA_signal_10368, mcs1_mcs_mat1_7_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, mcs1_mcs_mat1_7_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_11337, new_AGEMA_signal_11336, mcs1_mcs_mat1_7_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({new_AGEMA_signal_10371, new_AGEMA_signal_10370, mcs1_mcs_mat1_7_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3185], Fresh[3184], Fresh[3183]}), .c ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, mcs1_mcs_mat1_7_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3188], Fresh[3187], Fresh[3186]}), .c ({new_AGEMA_signal_9437, new_AGEMA_signal_9436, mcs1_mcs_mat1_7_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_11339, new_AGEMA_signal_11338, mcs1_mcs_mat1_7_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_12293, new_AGEMA_signal_12292, mcs1_mcs_mat1_7_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_9439, new_AGEMA_signal_9438, mcs1_mcs_mat1_7_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_10373, new_AGEMA_signal_10372, mcs1_mcs_mat1_7_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_12295, new_AGEMA_signal_12294, mcs1_mcs_mat1_7_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_8585, new_AGEMA_signal_8584, mcs1_mcs_mat1_7_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_12935, new_AGEMA_signal_12934, mcs1_mcs_mat1_7_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_11339, new_AGEMA_signal_11338, mcs1_mcs_mat1_7_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .c ({new_AGEMA_signal_12295, new_AGEMA_signal_12294, mcs1_mcs_mat1_7_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_7977, new_AGEMA_signal_7976, mcs1_mcs_mat1_7_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_10375, new_AGEMA_signal_10374, mcs1_mcs_mat1_7_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_11339, new_AGEMA_signal_11338, mcs1_mcs_mat1_7_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3191], Fresh[3190], Fresh[3189]}), .c ({new_AGEMA_signal_10375, new_AGEMA_signal_10374, mcs1_mcs_mat1_7_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3194], Fresh[3193], Fresh[3192]}), .c ({new_AGEMA_signal_8585, new_AGEMA_signal_8584, mcs1_mcs_mat1_7_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3197], Fresh[3196], Fresh[3195]}), .c ({new_AGEMA_signal_9439, new_AGEMA_signal_9438, mcs1_mcs_mat1_7_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_14785, new_AGEMA_signal_14784, mcs1_mcs_mat1_7_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_15265, new_AGEMA_signal_15264, mcs1_mcs_mat1_7_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_14335, new_AGEMA_signal_14334, mcs1_mcs_mat1_7_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_13911, new_AGEMA_signal_13910, mcs1_mcs_mat1_7_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_14785, new_AGEMA_signal_14784, mcs1_mcs_mat1_7_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_12937, new_AGEMA_signal_12936, mcs1_mcs_mat1_7_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_13909, new_AGEMA_signal_13908, mcs1_mcs_mat1_7_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_13911, new_AGEMA_signal_13910, mcs1_mcs_mat1_7_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_12937, new_AGEMA_signal_12936, mcs1_mcs_mat1_7_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_14333, new_AGEMA_signal_14332, mcs1_mcs_mat1_7_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_12297, new_AGEMA_signal_12296, mcs1_mcs_mat1_7_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_12299, new_AGEMA_signal_12298, mcs1_mcs_mat1_7_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_12937, new_AGEMA_signal_12936, mcs1_mcs_mat1_7_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_13481, new_AGEMA_signal_13480, mcs1_mcs_mat1_7_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .c ({new_AGEMA_signal_13911, new_AGEMA_signal_13910, mcs1_mcs_mat1_7_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_14787, new_AGEMA_signal_14786, mcs1_mcs_mat1_7_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_12297, new_AGEMA_signal_12296, mcs1_mcs_mat1_7_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_15267, new_AGEMA_signal_15266, mcs1_mcs_mat1_7_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_14335, new_AGEMA_signal_14334, mcs1_mcs_mat1_7_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_13481, new_AGEMA_signal_13480, mcs1_mcs_mat1_7_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_14787, new_AGEMA_signal_14786, mcs1_mcs_mat1_7_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .b ({new_AGEMA_signal_13913, new_AGEMA_signal_13912, mcs1_mcs_mat1_7_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_14335, new_AGEMA_signal_14334, mcs1_mcs_mat1_7_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3200], Fresh[3199], Fresh[3198]}), .c ({new_AGEMA_signal_13913, new_AGEMA_signal_13912, mcs1_mcs_mat1_7_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3203], Fresh[3202], Fresh[3201]}), .c ({new_AGEMA_signal_12299, new_AGEMA_signal_12298, mcs1_mcs_mat1_7_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3206], Fresh[3205], Fresh[3204]}), .c ({new_AGEMA_signal_13481, new_AGEMA_signal_13480, mcs1_mcs_mat1_7_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_11343, new_AGEMA_signal_11342, mcs1_mcs_mat1_7_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_9441, new_AGEMA_signal_9440, mcs1_mcs_mat1_7_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_12301, new_AGEMA_signal_12300, mcs1_mcs_mat1_7_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_10379, new_AGEMA_signal_10378, mcs1_mcs_mat1_7_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_12303, new_AGEMA_signal_12302, mcs1_mcs_mat1_7_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12939, new_AGEMA_signal_12938, mcs1_mcs_mat1_7_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_11343, new_AGEMA_signal_11342, mcs1_mcs_mat1_7_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_12303, new_AGEMA_signal_12302, mcs1_mcs_mat1_7_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_12941, new_AGEMA_signal_12940, mcs1_mcs_mat1_7_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_9441, new_AGEMA_signal_9440, mcs1_mcs_mat1_7_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_11345, new_AGEMA_signal_11344, mcs1_mcs_mat1_7_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_12303, new_AGEMA_signal_12302, mcs1_mcs_mat1_7_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, mcs1_mcs_mat1_7_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_9441, new_AGEMA_signal_9440, mcs1_mcs_mat1_7_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_10377, new_AGEMA_signal_10376, mcs1_mcs_mat1_7_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .c ({new_AGEMA_signal_11343, new_AGEMA_signal_11342, mcs1_mcs_mat1_7_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_9443, new_AGEMA_signal_9442, mcs1_mcs_mat1_7_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7979, new_AGEMA_signal_7978, mcs1_mcs_mat1_7_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_10377, new_AGEMA_signal_10376, mcs1_mcs_mat1_7_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_11345, new_AGEMA_signal_11344, mcs1_mcs_mat1_7_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_10379, new_AGEMA_signal_10378, mcs1_mcs_mat1_7_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_12305, new_AGEMA_signal_12304, mcs1_mcs_mat1_7_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_9443, new_AGEMA_signal_9442, mcs1_mcs_mat1_7_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_10379, new_AGEMA_signal_10378, mcs1_mcs_mat1_7_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({new_AGEMA_signal_10381, new_AGEMA_signal_10380, mcs1_mcs_mat1_7_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_11345, new_AGEMA_signal_11344, mcs1_mcs_mat1_7_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3209], Fresh[3208], Fresh[3207]}), .c ({new_AGEMA_signal_10381, new_AGEMA_signal_10380, mcs1_mcs_mat1_7_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, mcs1_mcs_mat1_7_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3215], Fresh[3214], Fresh[3213]}), .c ({new_AGEMA_signal_9443, new_AGEMA_signal_9442, mcs1_mcs_mat1_7_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_12309, new_AGEMA_signal_12308, mcs1_mcs_mat1_7_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_12943, new_AGEMA_signal_12942, mcs1_mcs_mat1_7_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({new_AGEMA_signal_11347, new_AGEMA_signal_11346, mcs1_mcs_mat1_7_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_12307, new_AGEMA_signal_12306, mcs1_mcs_mat1_7_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_12945, new_AGEMA_signal_12944, mcs1_mcs_mat1_7_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_9445, new_AGEMA_signal_9444, mcs1_mcs_mat1_7_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_13483, new_AGEMA_signal_13482, mcs1_mcs_mat1_7_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_12309, new_AGEMA_signal_12308, mcs1_mcs_mat1_7_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .c ({new_AGEMA_signal_12945, new_AGEMA_signal_12944, mcs1_mcs_mat1_7_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_7_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_11347, new_AGEMA_signal_11346, mcs1_mcs_mat1_7_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_12309, new_AGEMA_signal_12308, mcs1_mcs_mat1_7_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_7981, new_AGEMA_signal_7980, mcs1_mcs_mat1_7_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_10385, new_AGEMA_signal_10384, mcs1_mcs_mat1_7_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_11347, new_AGEMA_signal_11346, mcs1_mcs_mat1_7_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3218], Fresh[3217], Fresh[3216]}), .c ({new_AGEMA_signal_10385, new_AGEMA_signal_10384, mcs1_mcs_mat1_7_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3221], Fresh[3220], Fresh[3219]}), .c ({new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_7_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3224], Fresh[3223], Fresh[3222]}), .c ({new_AGEMA_signal_9445, new_AGEMA_signal_9444, mcs1_mcs_mat1_7_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_11353, new_AGEMA_signal_11352, mcs1_mcs_mat1_7_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_9447, new_AGEMA_signal_9446, mcs1_mcs_mat1_7_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_12311, new_AGEMA_signal_12310, mcs1_mcs_mat1_7_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_8591, new_AGEMA_signal_8590, mcs1_mcs_mat1_7_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_10387, new_AGEMA_signal_10386, mcs1_mcs_mat1_7_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_11349, new_AGEMA_signal_11348, mcs1_mcs_mat1_7_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({new_AGEMA_signal_10389, new_AGEMA_signal_10388, mcs1_mcs_mat1_7_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_11351, new_AGEMA_signal_11350, mcs1_mcs_mat1_7_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3227], Fresh[3226], Fresh[3225]}), .c ({new_AGEMA_signal_10389, new_AGEMA_signal_10388, mcs1_mcs_mat1_7_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3230], Fresh[3229], Fresh[3228]}), .c ({new_AGEMA_signal_8591, new_AGEMA_signal_8590, mcs1_mcs_mat1_7_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3233], Fresh[3232], Fresh[3231]}), .c ({new_AGEMA_signal_9447, new_AGEMA_signal_9446, mcs1_mcs_mat1_7_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_12317, new_AGEMA_signal_12316, mcs1_mcs_mat1_7_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_13485, new_AGEMA_signal_13484, mcs1_mcs_mat1_7_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_13915, new_AGEMA_signal_13914, mcs1_mcs_mat1_7_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_12319, new_AGEMA_signal_12318, mcs1_mcs_mat1_7_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_13917, new_AGEMA_signal_13916, mcs1_mcs_mat1_7_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_14339, new_AGEMA_signal_14338, mcs1_mcs_mat1_7_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_14341, new_AGEMA_signal_14340, mcs1_mcs_mat1_7_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_13919, new_AGEMA_signal_13918, mcs1_mcs_mat1_7_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_14789, new_AGEMA_signal_14788, mcs1_mcs_mat1_7_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_13921, new_AGEMA_signal_13920, mcs1_mcs_mat1_7_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_14341, new_AGEMA_signal_14340, mcs1_mcs_mat1_7_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3236], Fresh[3235], Fresh[3234]}), .c ({new_AGEMA_signal_13921, new_AGEMA_signal_13920, mcs1_mcs_mat1_7_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3239], Fresh[3238], Fresh[3237]}), .c ({new_AGEMA_signal_12319, new_AGEMA_signal_12318, mcs1_mcs_mat1_7_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({new_AGEMA_signal_13485, new_AGEMA_signal_13484, mcs1_mcs_mat1_7_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_10393, new_AGEMA_signal_10392, mcs1_mcs_mat1_7_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_11357, new_AGEMA_signal_11356, mcs1_mcs_mat1_7_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_12321, new_AGEMA_signal_12320, mcs1_mcs_mat1_7_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_12323, new_AGEMA_signal_12322, mcs1_mcs_mat1_7_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_10391, new_AGEMA_signal_10390, mcs1_mcs_mat1_7_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_12949, new_AGEMA_signal_12948, mcs1_mcs_mat1_7_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_9449, new_AGEMA_signal_9448, mcs1_mcs_mat1_7_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_10391, new_AGEMA_signal_10390, mcs1_mcs_mat1_7_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({new_AGEMA_signal_12323, new_AGEMA_signal_12322, mcs1_mcs_mat1_7_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_12951, new_AGEMA_signal_12950, mcs1_mcs_mat1_7_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_7985, new_AGEMA_signal_7984, mcs1_mcs_mat1_7_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_11357, new_AGEMA_signal_11356, mcs1_mcs_mat1_7_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_12323, new_AGEMA_signal_12322, mcs1_mcs_mat1_7_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, mcs1_mcs_mat1_7_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_10397, new_AGEMA_signal_10396, mcs1_mcs_mat1_7_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_11357, new_AGEMA_signal_11356, mcs1_mcs_mat1_7_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_10395, new_AGEMA_signal_10394, mcs1_mcs_mat1_7_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_11359, new_AGEMA_signal_11358, mcs1_mcs_mat1_7_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_12325, new_AGEMA_signal_12324, mcs1_mcs_mat1_7_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_10393, new_AGEMA_signal_10392, mcs1_mcs_mat1_7_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, mcs1_mcs_mat1_7_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_11359, new_AGEMA_signal_11358, mcs1_mcs_mat1_7_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_9449, new_AGEMA_signal_9448, mcs1_mcs_mat1_7_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_10393, new_AGEMA_signal_10392, mcs1_mcs_mat1_7_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3245], Fresh[3244], Fresh[3243]}), .c ({new_AGEMA_signal_10397, new_AGEMA_signal_10396, mcs1_mcs_mat1_7_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3248], Fresh[3247], Fresh[3246]}), .c ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, mcs1_mcs_mat1_7_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3251], Fresh[3250], Fresh[3249]}), .c ({new_AGEMA_signal_9449, new_AGEMA_signal_9448, mcs1_mcs_mat1_7_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_9453, new_AGEMA_signal_9452, mcs1_mcs_mat1_7_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_12953, new_AGEMA_signal_12952, mcs1_mcs_mat1_7_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_7_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_13487, new_AGEMA_signal_13486, mcs1_mcs_mat1_7_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_12327, new_AGEMA_signal_12326, mcs1_mcs_mat1_7_mcs_out[47]}), .b ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_12953, new_AGEMA_signal_12952, mcs1_mcs_mat1_7_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_11363, new_AGEMA_signal_11362, mcs1_mcs_mat1_7_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .c ({new_AGEMA_signal_12327, new_AGEMA_signal_12326, mcs1_mcs_mat1_7_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_7987, new_AGEMA_signal_7986, mcs1_mcs_mat1_7_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_10403, new_AGEMA_signal_10402, mcs1_mcs_mat1_7_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_11363, new_AGEMA_signal_11362, mcs1_mcs_mat1_7_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3254], Fresh[3253], Fresh[3252]}), .c ({new_AGEMA_signal_10403, new_AGEMA_signal_10402, mcs1_mcs_mat1_7_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3257], Fresh[3256], Fresh[3255]}), .c ({new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_7_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3260], Fresh[3259], Fresh[3258]}), .c ({new_AGEMA_signal_9453, new_AGEMA_signal_9452, mcs1_mcs_mat1_7_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_14343, new_AGEMA_signal_14342, mcs1_mcs_mat1_7_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_13489, new_AGEMA_signal_13488, mcs1_mcs_mat1_7_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_14791, new_AGEMA_signal_14790, mcs1_mcs_mat1_7_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_13923, new_AGEMA_signal_13922, mcs1_mcs_mat1_7_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_12329, new_AGEMA_signal_12328, mcs1_mcs_mat1_7_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_14343, new_AGEMA_signal_14342, mcs1_mcs_mat1_7_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_14345, new_AGEMA_signal_14344, mcs1_mcs_mat1_7_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_13927, new_AGEMA_signal_13926, mcs1_mcs_mat1_7_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_14793, new_AGEMA_signal_14792, mcs1_mcs_mat1_7_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_14347, new_AGEMA_signal_14346, mcs1_mcs_mat1_7_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_11365, new_AGEMA_signal_11364, mcs1_mcs_mat1_7_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_14795, new_AGEMA_signal_14794, mcs1_mcs_mat1_7_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_13923, new_AGEMA_signal_13922, mcs1_mcs_mat1_7_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_13491, new_AGEMA_signal_13490, mcs1_mcs_mat1_7_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_14347, new_AGEMA_signal_14346, mcs1_mcs_mat1_7_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_13925, new_AGEMA_signal_13924, mcs1_mcs_mat1_7_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_13491, new_AGEMA_signal_13490, mcs1_mcs_mat1_7_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_14349, new_AGEMA_signal_14348, mcs1_mcs_mat1_7_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3263], Fresh[3262], Fresh[3261]}), .c ({new_AGEMA_signal_13927, new_AGEMA_signal_13926, mcs1_mcs_mat1_7_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3266], Fresh[3265], Fresh[3264]}), .c ({new_AGEMA_signal_12329, new_AGEMA_signal_12328, mcs1_mcs_mat1_7_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3269], Fresh[3268], Fresh[3267]}), .c ({new_AGEMA_signal_13491, new_AGEMA_signal_13490, mcs1_mcs_mat1_7_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_12331, new_AGEMA_signal_12330, mcs1_mcs_mat1_7_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_7989, new_AGEMA_signal_7988, mcs1_mcs_mat1_7_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_12955, new_AGEMA_signal_12954, mcs1_mcs_mat1_7_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_9457, new_AGEMA_signal_9456, mcs1_mcs_mat1_7_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_9455, new_AGEMA_signal_9454, mcs1_mcs_mat1_7_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, mcs1_mcs_mat1_7_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({new_AGEMA_signal_12331, new_AGEMA_signal_12330, mcs1_mcs_mat1_7_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_12957, new_AGEMA_signal_12956, mcs1_mcs_mat1_7_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_7_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_11367, new_AGEMA_signal_11366, mcs1_mcs_mat1_7_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_12331, new_AGEMA_signal_12330, mcs1_mcs_mat1_7_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_10409, new_AGEMA_signal_10408, mcs1_mcs_mat1_7_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9459, new_AGEMA_signal_9458, mcs1_mcs_mat1_7_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_11367, new_AGEMA_signal_11366, mcs1_mcs_mat1_7_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_10409, new_AGEMA_signal_10408, mcs1_mcs_mat1_7_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_9457, new_AGEMA_signal_9456, mcs1_mcs_mat1_7_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_11369, new_AGEMA_signal_11368, mcs1_mcs_mat1_7_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_8815, new_AGEMA_signal_8814, mcs1_mcs_mat1_7_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_9457, new_AGEMA_signal_9456, mcs1_mcs_mat1_7_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({new_AGEMA_signal_8597, new_AGEMA_signal_8596, mcs1_mcs_mat1_7_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_8815, new_AGEMA_signal_8814, mcs1_mcs_mat1_7_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({new_AGEMA_signal_10409, new_AGEMA_signal_10408, mcs1_mcs_mat1_7_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3275], Fresh[3274], Fresh[3273]}), .c ({new_AGEMA_signal_8597, new_AGEMA_signal_8596, mcs1_mcs_mat1_7_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3278], Fresh[3277], Fresh[3276]}), .c ({new_AGEMA_signal_9459, new_AGEMA_signal_9458, mcs1_mcs_mat1_7_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, mcs1_mcs_mat1_7_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_9461, new_AGEMA_signal_9460, mcs1_mcs_mat1_7_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_11371, new_AGEMA_signal_11370, mcs1_mcs_mat1_7_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, mcs1_mcs_mat1_7_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_8817, new_AGEMA_signal_8816, mcs1_mcs_mat1_7_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_12959, new_AGEMA_signal_12958, mcs1_mcs_mat1_7_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_7_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_13493, new_AGEMA_signal_13492, mcs1_mcs_mat1_7_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3281], Fresh[3280], Fresh[3279]}), .c ({new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_7_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3284], Fresh[3283], Fresh[3282]}), .c ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, mcs1_mcs_mat1_7_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3287], Fresh[3286], Fresh[3285]}), .c ({new_AGEMA_signal_9461, new_AGEMA_signal_9460, mcs1_mcs_mat1_7_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_12335, new_AGEMA_signal_12334, mcs1_mcs_mat1_7_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_11375, new_AGEMA_signal_11374, mcs1_mcs_mat1_7_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_12961, new_AGEMA_signal_12960, mcs1_mcs_mat1_7_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_8603, new_AGEMA_signal_8602, mcs1_mcs_mat1_7_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_11377, new_AGEMA_signal_11376, mcs1_mcs_mat1_7_mcs_out[29]}), .c ({new_AGEMA_signal_12335, new_AGEMA_signal_12334, mcs1_mcs_mat1_7_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_8601, new_AGEMA_signal_8600, mcs1_mcs_mat1_7_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_11375, new_AGEMA_signal_11374, mcs1_mcs_mat1_7_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_12337, new_AGEMA_signal_12336, mcs1_mcs_mat1_7_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_7_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .c ({new_AGEMA_signal_11375, new_AGEMA_signal_11374, mcs1_mcs_mat1_7_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_12339, new_AGEMA_signal_12338, mcs1_mcs_mat1_7_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_10415, new_AGEMA_signal_10414, mcs1_mcs_mat1_7_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_12963, new_AGEMA_signal_12962, mcs1_mcs_mat1_7_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_11379, new_AGEMA_signal_11378, mcs1_mcs_mat1_7_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, mcs1_mcs_mat1_7_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_12339, new_AGEMA_signal_12338, mcs1_mcs_mat1_7_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_9463, new_AGEMA_signal_9462, mcs1_mcs_mat1_7_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, mcs1_mcs_mat1_7_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_7_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8603, new_AGEMA_signal_8602, mcs1_mcs_mat1_7_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_11379, new_AGEMA_signal_11378, mcs1_mcs_mat1_7_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3290], Fresh[3289], Fresh[3288]}), .c ({new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_7_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3293], Fresh[3292], Fresh[3291]}), .c ({new_AGEMA_signal_8603, new_AGEMA_signal_8602, mcs1_mcs_mat1_7_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3296], Fresh[3295], Fresh[3294]}), .c ({new_AGEMA_signal_9463, new_AGEMA_signal_9462, mcs1_mcs_mat1_7_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_13929, new_AGEMA_signal_13928, mcs1_mcs_mat1_7_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_14351, new_AGEMA_signal_14350, mcs1_mcs_mat1_7_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_13495, new_AGEMA_signal_13494, mcs1_mcs_mat1_7_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_12341, new_AGEMA_signal_12340, mcs1_mcs_mat1_7_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_13929, new_AGEMA_signal_13928, mcs1_mcs_mat1_7_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_14353, new_AGEMA_signal_14352, mcs1_mcs_mat1_7_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_14797, new_AGEMA_signal_14796, mcs1_mcs_mat1_7_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_13933, new_AGEMA_signal_13932, mcs1_mcs_mat1_7_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_12341, new_AGEMA_signal_12340, mcs1_mcs_mat1_7_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_14353, new_AGEMA_signal_14352, mcs1_mcs_mat1_7_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_14799, new_AGEMA_signal_14798, mcs1_mcs_mat1_7_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .c ({new_AGEMA_signal_15269, new_AGEMA_signal_15268, mcs1_mcs_mat1_7_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_13933, new_AGEMA_signal_13932, mcs1_mcs_mat1_7_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_14355, new_AGEMA_signal_14354, mcs1_mcs_mat1_7_mcs_out[24]}), .c ({new_AGEMA_signal_14799, new_AGEMA_signal_14798, mcs1_mcs_mat1_7_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_13931, new_AGEMA_signal_13930, mcs1_mcs_mat1_7_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .c ({new_AGEMA_signal_14355, new_AGEMA_signal_14354, mcs1_mcs_mat1_7_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_13495, new_AGEMA_signal_13494, mcs1_mcs_mat1_7_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_11381, new_AGEMA_signal_11380, mcs1_mcs_mat1_7_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_13931, new_AGEMA_signal_13930, mcs1_mcs_mat1_7_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3299], Fresh[3298], Fresh[3297]}), .c ({new_AGEMA_signal_13933, new_AGEMA_signal_13932, mcs1_mcs_mat1_7_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({new_AGEMA_signal_12341, new_AGEMA_signal_12340, mcs1_mcs_mat1_7_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3305], Fresh[3304], Fresh[3303]}), .c ({new_AGEMA_signal_13495, new_AGEMA_signal_13494, mcs1_mcs_mat1_7_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_10421, new_AGEMA_signal_10420, mcs1_mcs_mat1_7_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .c ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, mcs1_mcs_mat1_7_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_9465, new_AGEMA_signal_9464, mcs1_mcs_mat1_7_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, mcs1_mcs_mat1_7_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_10421, new_AGEMA_signal_10420, mcs1_mcs_mat1_7_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_11385, new_AGEMA_signal_11384, mcs1_mcs_mat1_7_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .c ({new_AGEMA_signal_12343, new_AGEMA_signal_12342, mcs1_mcs_mat1_7_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_7_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, mcs1_mcs_mat1_7_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_11385, new_AGEMA_signal_11384, mcs1_mcs_mat1_7_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_12345, new_AGEMA_signal_12344, mcs1_mcs_mat1_7_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_12965, new_AGEMA_signal_12964, mcs1_mcs_mat1_7_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_7_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_11387, new_AGEMA_signal_11386, mcs1_mcs_mat1_7_mcs_out[20]}), .c ({new_AGEMA_signal_12345, new_AGEMA_signal_12344, mcs1_mcs_mat1_7_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, mcs1_mcs_mat1_7_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_11387, new_AGEMA_signal_11386, mcs1_mcs_mat1_7_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_9465, new_AGEMA_signal_9464, mcs1_mcs_mat1_7_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_7995, new_AGEMA_signal_7994, mcs1_mcs_mat1_7_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, mcs1_mcs_mat1_7_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3308], Fresh[3307], Fresh[3306]}), .c ({new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_7_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3311], Fresh[3310], Fresh[3309]}), .c ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, mcs1_mcs_mat1_7_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3314], Fresh[3313], Fresh[3312]}), .c ({new_AGEMA_signal_9465, new_AGEMA_signal_9464, mcs1_mcs_mat1_7_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_10427, new_AGEMA_signal_10426, mcs1_mcs_mat1_7_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_10433, new_AGEMA_signal_10432, mcs1_mcs_mat1_7_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, mcs1_mcs_mat1_7_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_7_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_7997, new_AGEMA_signal_7996, mcs1_mcs_mat1_7_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_12347, new_AGEMA_signal_12346, mcs1_mcs_mat1_7_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_12349, new_AGEMA_signal_12348, mcs1_mcs_mat1_7_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_8607, new_AGEMA_signal_8606, mcs1_mcs_mat1_7_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_12967, new_AGEMA_signal_12966, mcs1_mcs_mat1_7_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_7_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_12349, new_AGEMA_signal_12348, mcs1_mcs_mat1_7_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, mcs1_mcs_mat1_7_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .c ({new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_7_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_9467, new_AGEMA_signal_9466, mcs1_mcs_mat1_7_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_9469, new_AGEMA_signal_9468, mcs1_mcs_mat1_7_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, mcs1_mcs_mat1_7_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_7_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_8607, new_AGEMA_signal_8606, mcs1_mcs_mat1_7_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_11393, new_AGEMA_signal_11392, mcs1_mcs_mat1_7_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3317], Fresh[3316], Fresh[3315]}), .c ({new_AGEMA_signal_10433, new_AGEMA_signal_10432, mcs1_mcs_mat1_7_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3320], Fresh[3319], Fresh[3318]}), .c ({new_AGEMA_signal_8607, new_AGEMA_signal_8606, mcs1_mcs_mat1_7_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3323], Fresh[3322], Fresh[3321]}), .c ({new_AGEMA_signal_9469, new_AGEMA_signal_9468, mcs1_mcs_mat1_7_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_12355, new_AGEMA_signal_12354, mcs1_mcs_mat1_7_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_8819, new_AGEMA_signal_8818, mcs1_mcs_mat1_7_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_12969, new_AGEMA_signal_12968, mcs1_mcs_mat1_7_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_11399, new_AGEMA_signal_11398, mcs1_mcs_mat1_7_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, mcs1_mcs_mat1_7_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_12351, new_AGEMA_signal_12350, mcs1_mcs_mat1_7_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_10437, new_AGEMA_signal_10436, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_8609, new_AGEMA_signal_8608, mcs1_mcs_mat1_7_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, mcs1_mcs_mat1_7_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_8819, new_AGEMA_signal_8818, mcs1_mcs_mat1_7_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_7_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_12353, new_AGEMA_signal_12352, mcs1_mcs_mat1_7_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, mcs1_mcs_mat1_7_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_10437, new_AGEMA_signal_10436, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_7_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_7999, new_AGEMA_signal_7998, mcs1_mcs_mat1_7_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_8609, new_AGEMA_signal_8608, mcs1_mcs_mat1_7_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_8819, new_AGEMA_signal_8818, mcs1_mcs_mat1_7_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_12971, new_AGEMA_signal_12970, mcs1_mcs_mat1_7_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_13497, new_AGEMA_signal_13496, mcs1_mcs_mat1_7_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_12355, new_AGEMA_signal_12354, mcs1_mcs_mat1_7_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_10437, new_AGEMA_signal_10436, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_12971, new_AGEMA_signal_12970, mcs1_mcs_mat1_7_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_11399, new_AGEMA_signal_11398, mcs1_mcs_mat1_7_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_12355, new_AGEMA_signal_12354, mcs1_mcs_mat1_7_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, mcs1_mcs_mat1_7_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_11399, new_AGEMA_signal_11398, mcs1_mcs_mat1_7_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, shiftr_out[96]}), .b ({new_AGEMA_signal_9471, new_AGEMA_signal_9470, mcs1_mcs_mat1_7_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, mcs1_mcs_mat1_7_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3326], Fresh[3325], Fresh[3324]}), .c ({new_AGEMA_signal_10437, new_AGEMA_signal_10436, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3329], Fresh[3328], Fresh[3327]}), .c ({new_AGEMA_signal_8609, new_AGEMA_signal_8608, mcs1_mcs_mat1_7_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({new_AGEMA_signal_9471, new_AGEMA_signal_9470, mcs1_mcs_mat1_7_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_12973, new_AGEMA_signal_12972, mcs1_mcs_mat1_7_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .c ({new_AGEMA_signal_13499, new_AGEMA_signal_13498, mcs1_mcs_mat1_7_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_14359, new_AGEMA_signal_14358, mcs1_mcs_mat1_7_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_14801, new_AGEMA_signal_14800, mcs1_mcs_mat1_7_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_13935, new_AGEMA_signal_13934, mcs1_mcs_mat1_7_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_14357, new_AGEMA_signal_14356, mcs1_mcs_mat1_7_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_13501, new_AGEMA_signal_13500, mcs1_mcs_mat1_7_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_12973, new_AGEMA_signal_12972, mcs1_mcs_mat1_7_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_13935, new_AGEMA_signal_13934, mcs1_mcs_mat1_7_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, mcs1_mcs_mat1_7_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_12357, new_AGEMA_signal_12356, mcs1_mcs_mat1_7_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_12973, new_AGEMA_signal_12972, mcs1_mcs_mat1_7_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_14803, new_AGEMA_signal_14802, mcs1_mcs_mat1_7_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, shiftr_out[64]}), .c ({new_AGEMA_signal_15271, new_AGEMA_signal_15270, mcs1_mcs_mat1_7_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, mcs1_mcs_mat1_7_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_14359, new_AGEMA_signal_14358, mcs1_mcs_mat1_7_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_14803, new_AGEMA_signal_14802, mcs1_mcs_mat1_7_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_13937, new_AGEMA_signal_13936, mcs1_mcs_mat1_7_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_13501, new_AGEMA_signal_13500, mcs1_mcs_mat1_7_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_14359, new_AGEMA_signal_14358, mcs1_mcs_mat1_7_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3335], Fresh[3334], Fresh[3333]}), .c ({new_AGEMA_signal_13937, new_AGEMA_signal_13936, mcs1_mcs_mat1_7_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3338], Fresh[3337], Fresh[3336]}), .c ({new_AGEMA_signal_12357, new_AGEMA_signal_12356, mcs1_mcs_mat1_7_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12376, shiftr_out[67]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3341], Fresh[3340], Fresh[3339]}), .c ({new_AGEMA_signal_13501, new_AGEMA_signal_13500, mcs1_mcs_mat1_7_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_13503, new_AGEMA_signal_13502, mcs1_mcs_mat1_7_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_9475, new_AGEMA_signal_9474, mcs1_mcs_mat1_7_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_13939, new_AGEMA_signal_13938, mcs1_mcs_mat1_7_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_12975, new_AGEMA_signal_12974, mcs1_mcs_mat1_7_mcs_out[7]}), .b ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .c ({new_AGEMA_signal_13503, new_AGEMA_signal_13502, mcs1_mcs_mat1_7_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_12359, new_AGEMA_signal_12358, mcs1_mcs_mat1_7_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .c ({new_AGEMA_signal_12975, new_AGEMA_signal_12974, mcs1_mcs_mat1_7_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_11403, new_AGEMA_signal_11402, mcs1_mcs_mat1_7_mcs_out[6]}), .b ({new_AGEMA_signal_8613, new_AGEMA_signal_8612, mcs1_mcs_mat1_7_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_12359, new_AGEMA_signal_12358, mcs1_mcs_mat1_7_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, mcs1_mcs_mat1_7_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_10439, new_AGEMA_signal_10438, mcs1_mcs_mat1_7_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_11403, new_AGEMA_signal_11402, mcs1_mcs_mat1_7_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, shiftr_out[33]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3344], Fresh[3343], Fresh[3342]}), .c ({new_AGEMA_signal_10439, new_AGEMA_signal_10438, mcs1_mcs_mat1_7_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, shiftr_out[34]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3347], Fresh[3346], Fresh[3345]}), .c ({new_AGEMA_signal_8613, new_AGEMA_signal_8612, mcs1_mcs_mat1_7_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3350], Fresh[3349], Fresh[3348]}), .c ({new_AGEMA_signal_9475, new_AGEMA_signal_9474, mcs1_mcs_mat1_7_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_9477, new_AGEMA_signal_9476, mcs1_mcs_mat1_7_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, mcs1_mcs_mat1_7_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_11407, new_AGEMA_signal_11406, mcs1_mcs_mat1_7_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .b ({new_AGEMA_signal_9479, new_AGEMA_signal_9478, mcs1_mcs_mat1_7_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, mcs1_mcs_mat1_7_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_11409, new_AGEMA_signal_11408, mcs1_mcs_mat1_7_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_8615, new_AGEMA_signal_8614, mcs1_mcs_mat1_7_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_12361, new_AGEMA_signal_12360, mcs1_mcs_mat1_7_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_11411, new_AGEMA_signal_11410, mcs1_mcs_mat1_7_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_10445, new_AGEMA_signal_10444, mcs1_mcs_mat1_7_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_12363, new_AGEMA_signal_12362, mcs1_mcs_mat1_7_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, mcs1_mcs_mat1_7_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_8003, new_AGEMA_signal_8002, mcs1_mcs_mat1_7_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_11411, new_AGEMA_signal_11410, mcs1_mcs_mat1_7_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, shiftr_out[1]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3353], Fresh[3352], Fresh[3351]}), .c ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, mcs1_mcs_mat1_7_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, shiftr_out[2]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3356], Fresh[3355], Fresh[3354]}), .c ({new_AGEMA_signal_8615, new_AGEMA_signal_8614, mcs1_mcs_mat1_7_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3359], Fresh[3358], Fresh[3357]}), .c ({new_AGEMA_signal_9479, new_AGEMA_signal_9478, mcs1_mcs_mat1_7_mcs_rom0_31_x3x4}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16141, new_AGEMA_signal_16140, mcs_out[128]}), .a ({new_AGEMA_signal_16181, new_AGEMA_signal_16180, y0_1[0]}), .c ({y0_s2[0], y0_s1[0], y0_s0[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15247, new_AGEMA_signal_15246, mcs_out[129]}), .a ({new_AGEMA_signal_15307, new_AGEMA_signal_15306, y0_1[1]}), .c ({y0_s2[1], y0_s1[1], y0_s0[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16139, new_AGEMA_signal_16138, mcs_out[130]}), .a ({new_AGEMA_signal_16215, new_AGEMA_signal_16214, y0_1[2]}), .c ({y0_s2[2], y0_s1[2], y0_s0[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14761, new_AGEMA_signal_14760, mcs_out[131]}), .a ({new_AGEMA_signal_14841, new_AGEMA_signal_14840, y0_1[3]}), .c ({y0_s2[3], y0_s1[3], y0_s0[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15713, new_AGEMA_signal_15712, mcs_out[132]}), .a ({new_AGEMA_signal_15823, new_AGEMA_signal_15822, y0_1[4]}), .c ({y0_s2[4], y0_s1[4], y0_s0[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16121, new_AGEMA_signal_16120, mcs_out[133]}), .a ({new_AGEMA_signal_16219, new_AGEMA_signal_16218, y0_1[5]}), .c ({y0_s2[5], y0_s1[5], y0_s0[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16119, new_AGEMA_signal_16118, mcs_out[134]}), .a ({new_AGEMA_signal_16225, new_AGEMA_signal_16224, y0_1[6]}), .c ({y0_s2[6], y0_s1[6], y0_s0[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15707, new_AGEMA_signal_15706, mcs_out[135]}), .a ({new_AGEMA_signal_15839, new_AGEMA_signal_15838, y0_1[7]}), .c ({y0_s2[7], y0_s1[7], y0_s0[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16377, new_AGEMA_signal_16376, mcs_out[136]}), .a ({new_AGEMA_signal_16439, new_AGEMA_signal_16438, y0_1[8]}), .c ({y0_s2[8], y0_s1[8], y0_s0[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14671, new_AGEMA_signal_14670, mcs_out[137]}), .a ({new_AGEMA_signal_14859, new_AGEMA_signal_14858, y0_1[9]}), .c ({y0_s2[9], y0_s1[9], y0_s0[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15677, new_AGEMA_signal_15676, mcs_out[138]}), .a ({new_AGEMA_signal_15801, new_AGEMA_signal_15800, y0_1[10]}), .c ({y0_s2[10], y0_s1[10], y0_s0[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16103, new_AGEMA_signal_16102, mcs_out[139]}), .a ({new_AGEMA_signal_16197, new_AGEMA_signal_16196, y0_1[11]}), .c ({y0_s2[11], y0_s1[11], y0_s0[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16089, new_AGEMA_signal_16088, mcs_out[140]}), .a ({new_AGEMA_signal_16201, new_AGEMA_signal_16200, y0_1[12]}), .c ({y0_s2[12], y0_s1[12], y0_s0[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14615, new_AGEMA_signal_14614, mcs_out[141]}), .a ({new_AGEMA_signal_14831, new_AGEMA_signal_14830, y0_1[13]}), .c ({y0_s2[13], y0_s1[13], y0_s0[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13733, new_AGEMA_signal_13732, mcs_out[142]}), .a ({new_AGEMA_signal_13953, new_AGEMA_signal_13952, y0_1[14]}), .c ({y0_s2[14], y0_s1[14], y0_s0[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15647, new_AGEMA_signal_15646, mcs_out[143]}), .a ({new_AGEMA_signal_15809, new_AGEMA_signal_15808, y0_1[15]}), .c ({y0_s2[15], y0_s1[15], y0_s0[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16067, new_AGEMA_signal_16066, mcs_out[144]}), .a ({new_AGEMA_signal_16203, new_AGEMA_signal_16202, y0_1[16]}), .c ({y0_s2[16], y0_s1[16], y0_s0[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15057, new_AGEMA_signal_15056, mcs_out[145]}), .a ({new_AGEMA_signal_15305, new_AGEMA_signal_15304, y0_1[17]}), .c ({y0_s2[17], y0_s1[17], y0_s0[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16065, new_AGEMA_signal_16064, mcs_out[146]}), .a ({new_AGEMA_signal_16205, new_AGEMA_signal_16204, y0_1[18]}), .c ({y0_s2[18], y0_s1[18], y0_s0[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14563, new_AGEMA_signal_14562, mcs_out[147]}), .a ({new_AGEMA_signal_14833, new_AGEMA_signal_14832, y0_1[19]}), .c ({y0_s2[19], y0_s1[19], y0_s0[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15575, new_AGEMA_signal_15574, mcs_out[148]}), .a ({new_AGEMA_signal_15811, new_AGEMA_signal_15810, y0_1[20]}), .c ({y0_s2[20], y0_s1[20], y0_s0[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16047, new_AGEMA_signal_16046, mcs_out[149]}), .a ({new_AGEMA_signal_16207, new_AGEMA_signal_16206, y0_1[21]}), .c ({y0_s2[21], y0_s1[21], y0_s0[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16045, new_AGEMA_signal_16044, mcs_out[150]}), .a ({new_AGEMA_signal_16209, new_AGEMA_signal_16208, y0_1[22]}), .c ({y0_s2[22], y0_s1[22], y0_s0[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15569, new_AGEMA_signal_15568, mcs_out[151]}), .a ({new_AGEMA_signal_15813, new_AGEMA_signal_15812, y0_1[23]}), .c ({y0_s2[23], y0_s1[23], y0_s0[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16365, new_AGEMA_signal_16364, mcs_out[152]}), .a ({new_AGEMA_signal_16437, new_AGEMA_signal_16436, y0_1[24]}), .c ({y0_s2[24], y0_s1[24], y0_s0[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14473, new_AGEMA_signal_14472, mcs_out[153]}), .a ({new_AGEMA_signal_14835, new_AGEMA_signal_14834, y0_1[25]}), .c ({y0_s2[25], y0_s1[25], y0_s0[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15539, new_AGEMA_signal_15538, mcs_out[154]}), .a ({new_AGEMA_signal_15815, new_AGEMA_signal_15814, y0_1[26]}), .c ({y0_s2[26], y0_s1[26], y0_s0[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16029, new_AGEMA_signal_16028, mcs_out[155]}), .a ({new_AGEMA_signal_16211, new_AGEMA_signal_16210, y0_1[27]}), .c ({y0_s2[27], y0_s1[27], y0_s0[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16015, new_AGEMA_signal_16014, mcs_out[156]}), .a ({new_AGEMA_signal_16213, new_AGEMA_signal_16212, y0_1[28]}), .c ({y0_s2[28], y0_s1[28], y0_s0[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14417, new_AGEMA_signal_14416, mcs_out[157]}), .a ({new_AGEMA_signal_14837, new_AGEMA_signal_14836, y0_1[29]}), .c ({y0_s2[29], y0_s1[29], y0_s0[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13515, new_AGEMA_signal_13514, mcs_out[158]}), .a ({new_AGEMA_signal_13955, new_AGEMA_signal_13954, y0_1[30]}), .c ({y0_s2[30], y0_s1[30], y0_s0[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15509, new_AGEMA_signal_15508, mcs_out[159]}), .a ({new_AGEMA_signal_15817, new_AGEMA_signal_15816, y0_1[31]}), .c ({y0_s2[31], y0_s1[31], y0_s0[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_32_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13893, new_AGEMA_signal_13892, mcs_out[160]}), .a ({new_AGEMA_signal_13957, new_AGEMA_signal_13956, y0_1[32]}), .c ({y0_s2[32], y0_s1[32], y0_s0[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_33_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14319, new_AGEMA_signal_14318, mcs_out[161]}), .a ({new_AGEMA_signal_14369, new_AGEMA_signal_14368, y0_1[33]}), .c ({y0_s2[33], y0_s1[33], y0_s0[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_34_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14317, new_AGEMA_signal_14316, mcs_out[162]}), .a ({new_AGEMA_signal_14371, new_AGEMA_signal_14370, y0_1[34]}), .c ({y0_s2[34], y0_s1[34], y0_s0[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_35_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14315, new_AGEMA_signal_14314, mcs_out[163]}), .a ({new_AGEMA_signal_14373, new_AGEMA_signal_14372, y0_1[35]}), .c ({y0_s2[35], y0_s1[35], y0_s0[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_36_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15195, new_AGEMA_signal_15194, mcs_out[164]}), .a ({new_AGEMA_signal_15309, new_AGEMA_signal_15308, y0_1[36]}), .c ({y0_s2[36], y0_s1[36], y0_s0[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_37_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13831, new_AGEMA_signal_13830, mcs_out[165]}), .a ({new_AGEMA_signal_13959, new_AGEMA_signal_13958, y0_1[37]}), .c ({y0_s2[37], y0_s1[37], y0_s0[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_38_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, mcs_out[166]}), .a ({new_AGEMA_signal_12977, new_AGEMA_signal_12976, y0_1[38]}), .c ({y0_s2[38], y0_s1[38], y0_s0[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_39_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14715, new_AGEMA_signal_14714, mcs_out[167]}), .a ({new_AGEMA_signal_14839, new_AGEMA_signal_14838, y0_1[39]}), .c ({y0_s2[39], y0_s1[39], y0_s0[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_40_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15671, new_AGEMA_signal_15670, mcs_out[168]}), .a ({new_AGEMA_signal_15819, new_AGEMA_signal_15818, y0_1[40]}), .c ({y0_s2[40], y0_s1[40], y0_s0[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_41_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15147, new_AGEMA_signal_15146, mcs_out[169]}), .a ({new_AGEMA_signal_15311, new_AGEMA_signal_15310, y0_1[41]}), .c ({y0_s2[41], y0_s1[41], y0_s0[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_42_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15145, new_AGEMA_signal_15144, mcs_out[170]}), .a ({new_AGEMA_signal_15313, new_AGEMA_signal_15312, y0_1[42]}), .c ({y0_s2[42], y0_s1[42], y0_s0[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_43_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15143, new_AGEMA_signal_15142, mcs_out[171]}), .a ({new_AGEMA_signal_15315, new_AGEMA_signal_15314, y0_1[43]}), .c ({y0_s2[43], y0_s1[43], y0_s0[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_44_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16087, new_AGEMA_signal_16086, mcs_out[172]}), .a ({new_AGEMA_signal_16217, new_AGEMA_signal_16216, y0_1[44]}), .c ({y0_s2[44], y0_s1[44], y0_s0[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_45_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14613, new_AGEMA_signal_14612, mcs_out[173]}), .a ({new_AGEMA_signal_14843, new_AGEMA_signal_14842, y0_1[45]}), .c ({y0_s2[45], y0_s1[45], y0_s0[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_46_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14611, new_AGEMA_signal_14610, mcs_out[174]}), .a ({new_AGEMA_signal_14845, new_AGEMA_signal_14844, y0_1[46]}), .c ({y0_s2[46], y0_s1[46], y0_s0[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_47_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15641, new_AGEMA_signal_15640, mcs_out[175]}), .a ({new_AGEMA_signal_15821, new_AGEMA_signal_15820, y0_1[47]}), .c ({y0_s2[47], y0_s1[47], y0_s0[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_48_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13675, new_AGEMA_signal_13674, mcs_out[176]}), .a ({new_AGEMA_signal_13961, new_AGEMA_signal_13960, y0_1[48]}), .c ({y0_s2[48], y0_s1[48], y0_s0[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_49_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14133, new_AGEMA_signal_14132, mcs_out[177]}), .a ({new_AGEMA_signal_14375, new_AGEMA_signal_14374, y0_1[49]}), .c ({y0_s2[49], y0_s1[49], y0_s0[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_50_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14131, new_AGEMA_signal_14130, mcs_out[178]}), .a ({new_AGEMA_signal_14377, new_AGEMA_signal_14376, y0_1[50]}), .c ({y0_s2[50], y0_s1[50], y0_s0[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_51_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14129, new_AGEMA_signal_14128, mcs_out[179]}), .a ({new_AGEMA_signal_14379, new_AGEMA_signal_14378, y0_1[51]}), .c ({y0_s2[51], y0_s1[51], y0_s0[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_52_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15005, new_AGEMA_signal_15004, mcs_out[180]}), .a ({new_AGEMA_signal_15317, new_AGEMA_signal_15316, y0_1[52]}), .c ({y0_s2[52], y0_s1[52], y0_s0[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_53_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13613, new_AGEMA_signal_13612, mcs_out[181]}), .a ({new_AGEMA_signal_13963, new_AGEMA_signal_13962, y0_1[53]}), .c ({y0_s2[53], y0_s1[53], y0_s0[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_54_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_12547, new_AGEMA_signal_12546, mcs_out[182]}), .a ({new_AGEMA_signal_12979, new_AGEMA_signal_12978, y0_1[54]}), .c ({y0_s2[54], y0_s1[54], y0_s0[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_55_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14517, new_AGEMA_signal_14516, mcs_out[183]}), .a ({new_AGEMA_signal_14847, new_AGEMA_signal_14846, y0_1[55]}), .c ({y0_s2[55], y0_s1[55], y0_s0[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_56_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15533, new_AGEMA_signal_15532, mcs_out[184]}), .a ({new_AGEMA_signal_15825, new_AGEMA_signal_15824, y0_1[56]}), .c ({y0_s2[56], y0_s1[56], y0_s0[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_57_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14957, new_AGEMA_signal_14956, mcs_out[185]}), .a ({new_AGEMA_signal_15319, new_AGEMA_signal_15318, y0_1[57]}), .c ({y0_s2[57], y0_s1[57], y0_s0[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_58_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14955, new_AGEMA_signal_14954, mcs_out[186]}), .a ({new_AGEMA_signal_15321, new_AGEMA_signal_15320, y0_1[58]}), .c ({y0_s2[58], y0_s1[58], y0_s0[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_59_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14953, new_AGEMA_signal_14952, mcs_out[187]}), .a ({new_AGEMA_signal_15323, new_AGEMA_signal_15322, y0_1[59]}), .c ({y0_s2[59], y0_s1[59], y0_s0[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_60_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16013, new_AGEMA_signal_16012, mcs_out[188]}), .a ({new_AGEMA_signal_16221, new_AGEMA_signal_16220, y0_1[60]}), .c ({y0_s2[60], y0_s1[60], y0_s0[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_61_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14415, new_AGEMA_signal_14414, mcs_out[189]}), .a ({new_AGEMA_signal_14849, new_AGEMA_signal_14848, y0_1[61]}), .c ({y0_s2[61], y0_s1[61], y0_s0[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_62_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14413, new_AGEMA_signal_14412, mcs_out[190]}), .a ({new_AGEMA_signal_14851, new_AGEMA_signal_14850, y0_1[62]}), .c ({y0_s2[62], y0_s1[62], y0_s0[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_63_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15503, new_AGEMA_signal_15502, mcs_out[191]}), .a ({new_AGEMA_signal_15827, new_AGEMA_signal_15826, y0_1[63]}), .c ({y0_s2[63], y0_s1[63], y0_s0[63]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_64_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16137, new_AGEMA_signal_16136, mcs_out[192]}), .a ({new_AGEMA_signal_16223, new_AGEMA_signal_16222, y0_1[64]}), .c ({y0_s2[64], y0_s1[64], y0_s0[64]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_65_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15745, new_AGEMA_signal_15744, mcs_out[193]}), .a ({new_AGEMA_signal_15829, new_AGEMA_signal_15828, y0_1[65]}), .c ({y0_s2[65], y0_s1[65], y0_s0[65]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_66_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15743, new_AGEMA_signal_15742, mcs_out[194]}), .a ({new_AGEMA_signal_15831, new_AGEMA_signal_15830, y0_1[66]}), .c ({y0_s2[66], y0_s1[66], y0_s0[66]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_67_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15741, new_AGEMA_signal_15740, mcs_out[195]}), .a ({new_AGEMA_signal_15833, new_AGEMA_signal_15832, y0_1[67]}), .c ({y0_s2[67], y0_s1[67], y0_s0[67]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_68_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs_out[196]}), .a ({new_AGEMA_signal_15835, new_AGEMA_signal_15834, y0_1[68]}), .c ({y0_s2[68], y0_s1[68], y0_s0[68]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_69_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15191, new_AGEMA_signal_15190, mcs_out[197]}), .a ({new_AGEMA_signal_15325, new_AGEMA_signal_15324, y0_1[69]}), .c ({y0_s2[69], y0_s1[69], y0_s0[69]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_70_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14711, new_AGEMA_signal_14710, mcs_out[198]}), .a ({new_AGEMA_signal_14853, new_AGEMA_signal_14852, y0_1[70]}), .c ({y0_s2[70], y0_s1[70], y0_s0[70]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_71_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, mcs_out[199]}), .a ({new_AGEMA_signal_15837, new_AGEMA_signal_15836, y0_1[71]}), .c ({y0_s2[71], y0_s1[71], y0_s0[71]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_72_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16469, new_AGEMA_signal_16468, mcs_out[200]}), .a ({new_AGEMA_signal_16545, new_AGEMA_signal_16544, y0_1[72]}), .c ({y0_s2[72], y0_s1[72], y0_s0[72]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_73_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14221, new_AGEMA_signal_14220, mcs_out[201]}), .a ({new_AGEMA_signal_14381, new_AGEMA_signal_14380, y0_1[73]}), .c ({y0_s2[73], y0_s1[73], y0_s0[73]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_74_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15141, new_AGEMA_signal_15140, mcs_out[202]}), .a ({new_AGEMA_signal_15327, new_AGEMA_signal_15326, y0_1[74]}), .c ({y0_s2[74], y0_s1[74], y0_s0[74]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_75_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16101, new_AGEMA_signal_16100, mcs_out[203]}), .a ({new_AGEMA_signal_16227, new_AGEMA_signal_16226, y0_1[75]}), .c ({y0_s2[75], y0_s1[75], y0_s0[75]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_76_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16085, new_AGEMA_signal_16084, mcs_out[204]}), .a ({new_AGEMA_signal_16229, new_AGEMA_signal_16228, y0_1[76]}), .c ({y0_s2[76], y0_s1[76], y0_s0[76]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_77_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16083, new_AGEMA_signal_16082, mcs_out[205]}), .a ({new_AGEMA_signal_16231, new_AGEMA_signal_16230, y0_1[77]}), .c ({y0_s2[77], y0_s1[77], y0_s0[77]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_78_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16081, new_AGEMA_signal_16080, mcs_out[206]}), .a ({new_AGEMA_signal_16233, new_AGEMA_signal_16232, y0_1[78]}), .c ({y0_s2[78], y0_s1[78], y0_s0[78]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_79_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16079, new_AGEMA_signal_16078, mcs_out[207]}), .a ({new_AGEMA_signal_16235, new_AGEMA_signal_16234, y0_1[79]}), .c ({y0_s2[79], y0_s1[79], y0_s0[79]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_80_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16063, new_AGEMA_signal_16062, mcs_out[208]}), .a ({new_AGEMA_signal_16237, new_AGEMA_signal_16236, y0_1[80]}), .c ({y0_s2[80], y0_s1[80], y0_s0[80]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_81_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15607, new_AGEMA_signal_15606, mcs_out[209]}), .a ({new_AGEMA_signal_15841, new_AGEMA_signal_15840, y0_1[81]}), .c ({y0_s2[81], y0_s1[81], y0_s0[81]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_82_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15605, new_AGEMA_signal_15604, mcs_out[210]}), .a ({new_AGEMA_signal_15843, new_AGEMA_signal_15842, y0_1[82]}), .c ({y0_s2[82], y0_s1[82], y0_s0[82]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_83_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15603, new_AGEMA_signal_15602, mcs_out[211]}), .a ({new_AGEMA_signal_15845, new_AGEMA_signal_15844, y0_1[83]}), .c ({y0_s2[83], y0_s1[83], y0_s0[83]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_84_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15567, new_AGEMA_signal_15566, mcs_out[212]}), .a ({new_AGEMA_signal_15847, new_AGEMA_signal_15846, y0_1[84]}), .c ({y0_s2[84], y0_s1[84], y0_s0[84]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_85_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15001, new_AGEMA_signal_15000, mcs_out[213]}), .a ({new_AGEMA_signal_15329, new_AGEMA_signal_15328, y0_1[85]}), .c ({y0_s2[85], y0_s1[85], y0_s0[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_86_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14513, new_AGEMA_signal_14512, mcs_out[214]}), .a ({new_AGEMA_signal_14855, new_AGEMA_signal_14854, y0_1[86]}), .c ({y0_s2[86], y0_s1[86], y0_s0[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_87_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15565, new_AGEMA_signal_15564, mcs_out[215]}), .a ({new_AGEMA_signal_15849, new_AGEMA_signal_15848, y0_1[87]}), .c ({y0_s2[87], y0_s1[87], y0_s0[87]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_88_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16465, new_AGEMA_signal_16464, mcs_out[216]}), .a ({new_AGEMA_signal_16547, new_AGEMA_signal_16546, y0_1[88]}), .c ({y0_s2[88], y0_s1[88], y0_s0[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_89_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14035, new_AGEMA_signal_14034, mcs_out[217]}), .a ({new_AGEMA_signal_14383, new_AGEMA_signal_14382, y0_1[89]}), .c ({y0_s2[89], y0_s1[89], y0_s0[89]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_90_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14951, new_AGEMA_signal_14950, mcs_out[218]}), .a ({new_AGEMA_signal_15331, new_AGEMA_signal_15330, y0_1[90]}), .c ({y0_s2[90], y0_s1[90], y0_s0[90]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_91_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16027, new_AGEMA_signal_16026, mcs_out[219]}), .a ({new_AGEMA_signal_16239, new_AGEMA_signal_16238, y0_1[91]}), .c ({y0_s2[91], y0_s1[91], y0_s0[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_92_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16011, new_AGEMA_signal_16010, mcs_out[220]}), .a ({new_AGEMA_signal_16241, new_AGEMA_signal_16240, y0_1[92]}), .c ({y0_s2[92], y0_s1[92], y0_s0[92]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_93_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16009, new_AGEMA_signal_16008, mcs_out[221]}), .a ({new_AGEMA_signal_16243, new_AGEMA_signal_16242, y0_1[93]}), .c ({y0_s2[93], y0_s1[93], y0_s0[93]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_94_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16007, new_AGEMA_signal_16006, mcs_out[222]}), .a ({new_AGEMA_signal_16245, new_AGEMA_signal_16244, y0_1[94]}), .c ({y0_s2[94], y0_s1[94], y0_s0[94]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_95_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16005, new_AGEMA_signal_16004, mcs_out[223]}), .a ({new_AGEMA_signal_16247, new_AGEMA_signal_16246, y0_1[95]}), .c ({y0_s2[95], y0_s1[95], y0_s0[95]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_96_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15739, new_AGEMA_signal_15738, mcs_out[224]}), .a ({new_AGEMA_signal_15851, new_AGEMA_signal_15850, y0_1[96]}), .c ({y0_s2[96], y0_s1[96], y0_s0[96]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_97_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16135, new_AGEMA_signal_16134, mcs_out[225]}), .a ({new_AGEMA_signal_16249, new_AGEMA_signal_16248, y0_1[97]}), .c ({y0_s2[97], y0_s1[97], y0_s0[97]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_98_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14757, new_AGEMA_signal_14756, mcs_out[226]}), .a ({new_AGEMA_signal_14857, new_AGEMA_signal_14856, y0_1[98]}), .c ({y0_s2[98], y0_s1[98], y0_s0[98]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_99_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16133, new_AGEMA_signal_16132, mcs_out[227]}), .a ({new_AGEMA_signal_16251, new_AGEMA_signal_16250, y0_1[99]}), .c ({y0_s2[99], y0_s1[99], y0_s0[99]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_100_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15187, new_AGEMA_signal_15186, mcs_out[228]}), .a ({new_AGEMA_signal_15297, new_AGEMA_signal_15296, y0_1[100]}), .c ({y0_s2[100], y0_s1[100], y0_s0[100]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_101_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15701, new_AGEMA_signal_15700, mcs_out[229]}), .a ({new_AGEMA_signal_15797, new_AGEMA_signal_15796, y0_1[101]}), .c ({y0_s2[101], y0_s1[101], y0_s0[101]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_102_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16117, new_AGEMA_signal_16116, mcs_out[230]}), .a ({new_AGEMA_signal_16183, new_AGEMA_signal_16182, y0_1[102]}), .c ({y0_s2[102], y0_s1[102], y0_s0[102]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_103_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16115, new_AGEMA_signal_16114, mcs_out[231]}), .a ({new_AGEMA_signal_16185, new_AGEMA_signal_16184, y0_1[103]}), .c ({y0_s2[103], y0_s1[103], y0_s0[103]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_104_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16099, new_AGEMA_signal_16098, mcs_out[232]}), .a ({new_AGEMA_signal_16187, new_AGEMA_signal_16186, y0_1[104]}), .c ({y0_s2[104], y0_s1[104], y0_s0[104]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_105_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14661, new_AGEMA_signal_14660, mcs_out[233]}), .a ({new_AGEMA_signal_14825, new_AGEMA_signal_14824, y0_1[105]}), .c ({y0_s2[105], y0_s1[105], y0_s0[105]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_106_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15137, new_AGEMA_signal_15136, mcs_out[234]}), .a ({new_AGEMA_signal_15299, new_AGEMA_signal_15298, y0_1[106]}), .c ({y0_s2[106], y0_s1[106], y0_s0[106]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_107_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15665, new_AGEMA_signal_15664, mcs_out[235]}), .a ({new_AGEMA_signal_15799, new_AGEMA_signal_15798, y0_1[107]}), .c ({y0_s2[107], y0_s1[107], y0_s0[107]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_108_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13731, new_AGEMA_signal_13730, mcs_out[236]}), .a ({new_AGEMA_signal_13945, new_AGEMA_signal_13944, y0_1[108]}), .c ({y0_s2[108], y0_s1[108], y0_s0[108]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_109_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14179, new_AGEMA_signal_14178, mcs_out[237]}), .a ({new_AGEMA_signal_14361, new_AGEMA_signal_14360, y0_1[109]}), .c ({y0_s2[109], y0_s1[109], y0_s0[109]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_110_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14177, new_AGEMA_signal_14176, mcs_out[238]}), .a ({new_AGEMA_signal_14363, new_AGEMA_signal_14362, y0_1[110]}), .c ({y0_s2[110], y0_s1[110], y0_s0[110]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_111_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13725, new_AGEMA_signal_13724, mcs_out[239]}), .a ({new_AGEMA_signal_13947, new_AGEMA_signal_13946, y0_1[111]}), .c ({y0_s2[111], y0_s1[111], y0_s0[111]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_112_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15601, new_AGEMA_signal_15600, mcs_out[240]}), .a ({new_AGEMA_signal_15803, new_AGEMA_signal_15802, y0_1[112]}), .c ({y0_s2[112], y0_s1[112], y0_s0[112]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_113_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16061, new_AGEMA_signal_16060, mcs_out[241]}), .a ({new_AGEMA_signal_16189, new_AGEMA_signal_16188, y0_1[113]}), .c ({y0_s2[113], y0_s1[113], y0_s0[113]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_114_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14559, new_AGEMA_signal_14558, mcs_out[242]}), .a ({new_AGEMA_signal_14827, new_AGEMA_signal_14826, y0_1[114]}), .c ({y0_s2[114], y0_s1[114], y0_s0[114]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_115_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16059, new_AGEMA_signal_16058, mcs_out[243]}), .a ({new_AGEMA_signal_16191, new_AGEMA_signal_16190, y0_1[115]}), .c ({y0_s2[115], y0_s1[115], y0_s0[115]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_116_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14997, new_AGEMA_signal_14996, mcs_out[244]}), .a ({new_AGEMA_signal_15301, new_AGEMA_signal_15300, y0_1[116]}), .c ({y0_s2[116], y0_s1[116], y0_s0[116]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_117_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15563, new_AGEMA_signal_15562, mcs_out[245]}), .a ({new_AGEMA_signal_15805, new_AGEMA_signal_15804, y0_1[117]}), .c ({y0_s2[117], y0_s1[117], y0_s0[117]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_118_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16043, new_AGEMA_signal_16042, mcs_out[246]}), .a ({new_AGEMA_signal_16193, new_AGEMA_signal_16192, y0_1[118]}), .c ({y0_s2[118], y0_s1[118], y0_s0[118]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_119_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16041, new_AGEMA_signal_16040, mcs_out[247]}), .a ({new_AGEMA_signal_16195, new_AGEMA_signal_16194, y0_1[119]}), .c ({y0_s2[119], y0_s1[119], y0_s0[119]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_120_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16025, new_AGEMA_signal_16024, mcs_out[248]}), .a ({new_AGEMA_signal_16199, new_AGEMA_signal_16198, y0_1[120]}), .c ({y0_s2[120], y0_s1[120], y0_s0[120]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_121_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14463, new_AGEMA_signal_14462, mcs_out[249]}), .a ({new_AGEMA_signal_14829, new_AGEMA_signal_14828, y0_1[121]}), .c ({y0_s2[121], y0_s1[121], y0_s0[121]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_122_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14947, new_AGEMA_signal_14946, mcs_out[250]}), .a ({new_AGEMA_signal_15303, new_AGEMA_signal_15302, y0_1[122]}), .c ({y0_s2[122], y0_s1[122], y0_s0[122]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_123_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15527, new_AGEMA_signal_15526, mcs_out[251]}), .a ({new_AGEMA_signal_15807, new_AGEMA_signal_15806, y0_1[123]}), .c ({y0_s2[123], y0_s1[123], y0_s0[123]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_124_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13513, new_AGEMA_signal_13512, mcs_out[252]}), .a ({new_AGEMA_signal_13949, new_AGEMA_signal_13948, y0_1[124]}), .c ({y0_s2[124], y0_s1[124], y0_s0[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_125_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13993, new_AGEMA_signal_13992, mcs_out[253]}), .a ({new_AGEMA_signal_14365, new_AGEMA_signal_14364, y0_1[125]}), .c ({y0_s2[125], y0_s1[125], y0_s0[125]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_126_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13991, new_AGEMA_signal_13990, mcs_out[254]}), .a ({new_AGEMA_signal_14367, new_AGEMA_signal_14366, y0_1[126]}), .c ({y0_s2[126], y0_s1[126], y0_s0[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MUX_inst2_MUXInst_127_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_13507, new_AGEMA_signal_13506, mcs_out[255]}), .a ({new_AGEMA_signal_13951, new_AGEMA_signal_13950, y0_1[127]}), .c ({y0_s2[127], y0_s1[127], y0_s0[127]}) ) ;

endmodule
