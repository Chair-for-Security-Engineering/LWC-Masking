/* modified netlist. Source: module xoodoo_round in file ./test/xoodoo_round.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module xoodoo_round_HPC2_ClockGating_d2 (state_in_s0, rc, clk, state_in_s1, state_in_s2, Fresh, /*rst,*/ state_out_s0, state_out_s1, state_out_s2/*, Synch*/);
    input [383:0] state_in_s0 ;
    input [31:0] rc ;
    input clk ;
    input [383:0] state_in_s1 ;
    input [383:0] state_in_s2 ;
    //input rst ;
    input [1151:0] Fresh ;
    output [383:0] state_out_s0 ;
    output [383:0] state_out_s1 ;
    output [383:0] state_out_s2 ;
    //output Synch ;
    wire rd_I_n2624 ;
    wire rd_I_n2623 ;
    wire rd_I_n2622 ;
    wire rd_I_n2621 ;
    wire rd_I_n2620 ;
    wire rd_I_n2619 ;
    wire rd_I_n2618 ;
    wire rd_I_n2617 ;
    wire rd_I_n2616 ;
    wire rd_I_n2615 ;
    wire rd_I_n2614 ;
    wire rd_I_n2613 ;
    wire rd_I_n2612 ;
    wire rd_I_n2611 ;
    wire rd_I_n2610 ;
    wire rd_I_n2609 ;
    wire rd_I_n2608 ;
    wire rd_I_n2607 ;
    wire rd_I_n2606 ;
    wire rd_I_n2605 ;
    wire rd_I_n2604 ;
    wire rd_I_n2603 ;
    wire rd_I_n2602 ;
    wire rd_I_n2601 ;
    wire rd_I_n2600 ;
    wire rd_I_n2599 ;
    wire rd_I_n2598 ;
    wire rd_I_n2597 ;
    wire rd_I_n2596 ;
    wire rd_I_n2595 ;
    wire rd_I_n2594 ;
    wire rd_I_n2593 ;
    wire rd_I_n2592 ;
    wire rd_I_n2591 ;
    wire rd_I_n2590 ;
    wire rd_I_n2589 ;
    wire rd_I_n2588 ;
    wire rd_I_n2587 ;
    wire rd_I_n2586 ;
    wire rd_I_n2585 ;
    wire rd_I_n2584 ;
    wire rd_I_n2583 ;
    wire rd_I_n2582 ;
    wire rd_I_n2581 ;
    wire rd_I_n2580 ;
    wire rd_I_n2579 ;
    wire rd_I_n2578 ;
    wire rd_I_n2577 ;
    wire rd_I_n2576 ;
    wire rd_I_n2575 ;
    wire rd_I_n2574 ;
    wire rd_I_n2573 ;
    wire rd_I_n2572 ;
    wire rd_I_n2571 ;
    wire rd_I_n2570 ;
    wire rd_I_n2569 ;
    wire rd_I_n2568 ;
    wire rd_I_n2567 ;
    wire rd_I_n2566 ;
    wire rd_I_n2565 ;
    wire rd_I_n2564 ;
    wire rd_I_n2563 ;
    wire rd_I_n2562 ;
    wire rd_I_n2561 ;
    wire rd_I_n2560 ;
    wire rd_I_n2559 ;
    wire rd_I_n2558 ;
    wire rd_I_n2557 ;
    wire rd_I_n2556 ;
    wire rd_I_n2555 ;
    wire rd_I_n2554 ;
    wire rd_I_n2553 ;
    wire rd_I_n2552 ;
    wire rd_I_n2551 ;
    wire rd_I_n2550 ;
    wire rd_I_n2549 ;
    wire rd_I_n2548 ;
    wire rd_I_n2547 ;
    wire rd_I_n2546 ;
    wire rd_I_n2545 ;
    wire rd_I_n2544 ;
    wire rd_I_n2543 ;
    wire rd_I_n2542 ;
    wire rd_I_n2541 ;
    wire rd_I_n2540 ;
    wire rd_I_n2539 ;
    wire rd_I_n2538 ;
    wire rd_I_n2537 ;
    wire rd_I_n2536 ;
    wire rd_I_n2535 ;
    wire rd_I_n2534 ;
    wire rd_I_n2533 ;
    wire rd_I_n2532 ;
    wire rd_I_n2531 ;
    wire rd_I_n2530 ;
    wire rd_I_n2529 ;
    wire rd_I_n2528 ;
    wire rd_I_n2527 ;
    wire rd_I_n2526 ;
    wire rd_I_n2525 ;
    wire rd_I_n2524 ;
    wire rd_I_n2523 ;
    wire rd_I_n2522 ;
    wire rd_I_n2521 ;
    wire rd_I_n2520 ;
    wire rd_I_n2519 ;
    wire rd_I_n2518 ;
    wire rd_I_n2517 ;
    wire rd_I_n2516 ;
    wire rd_I_n2515 ;
    wire rd_I_n2514 ;
    wire rd_I_n2513 ;
    wire rd_I_n2512 ;
    wire rd_I_n2511 ;
    wire rd_I_n2510 ;
    wire rd_I_n2509 ;
    wire rd_I_n2508 ;
    wire rd_I_n2507 ;
    wire rd_I_n2506 ;
    wire rd_I_n2505 ;
    wire rd_I_n2504 ;
    wire rd_I_n2503 ;
    wire rd_I_n2502 ;
    wire rd_I_n2501 ;
    wire rd_I_n2500 ;
    wire rd_I_n2499 ;
    wire rd_I_n2498 ;
    wire rd_I_n2497 ;
    wire rd_I_n2496 ;
    wire rd_I_n2495 ;
    wire rd_I_n2494 ;
    wire rd_I_n2493 ;
    wire rd_I_n2492 ;
    wire rd_I_n2491 ;
    wire rd_I_n2490 ;
    wire rd_I_n2489 ;
    wire rd_I_n2488 ;
    wire rd_I_n2487 ;
    wire rd_I_n2486 ;
    wire rd_I_n2485 ;
    wire rd_I_n2484 ;
    wire rd_I_n2483 ;
    wire rd_I_n2482 ;
    wire rd_I_n2481 ;
    wire rd_I_n2480 ;
    wire rd_I_n2479 ;
    wire rd_I_n2478 ;
    wire rd_I_n2477 ;
    wire rd_I_n2476 ;
    wire rd_I_n2475 ;
    wire rd_I_n2474 ;
    wire rd_I_n2473 ;
    wire rd_I_n2472 ;
    wire rd_I_n2471 ;
    wire rd_I_n2470 ;
    wire rd_I_n2469 ;
    wire rd_I_n2468 ;
    wire rd_I_n2467 ;
    wire rd_I_n2466 ;
    wire rd_I_n2465 ;
    wire rd_I_n2464 ;
    wire rd_I_n2463 ;
    wire rd_I_n2462 ;
    wire rd_I_n2461 ;
    wire rd_I_n2460 ;
    wire rd_I_n2459 ;
    wire rd_I_n2458 ;
    wire rd_I_n2457 ;
    wire rd_I_n2456 ;
    wire rd_I_n2455 ;
    wire rd_I_n2454 ;
    wire rd_I_n2453 ;
    wire rd_I_n2452 ;
    wire rd_I_n2451 ;
    wire rd_I_n2450 ;
    wire rd_I_n2449 ;
    wire rd_I_n2448 ;
    wire rd_I_n2447 ;
    wire rd_I_n2446 ;
    wire rd_I_n2445 ;
    wire rd_I_n2444 ;
    wire rd_I_n2443 ;
    wire rd_I_n2442 ;
    wire rd_I_n2441 ;
    wire rd_I_n2440 ;
    wire rd_I_n2439 ;
    wire rd_I_n2438 ;
    wire rd_I_n2437 ;
    wire rd_I_n2436 ;
    wire rd_I_n2435 ;
    wire rd_I_n2434 ;
    wire rd_I_n2433 ;
    wire rd_I_n2432 ;
    wire rd_I_n2431 ;
    wire rd_I_n2430 ;
    wire rd_I_n2429 ;
    wire rd_I_n2428 ;
    wire rd_I_n2427 ;
    wire rd_I_n2426 ;
    wire rd_I_n2425 ;
    wire rd_I_n2424 ;
    wire rd_I_n2423 ;
    wire rd_I_n2422 ;
    wire rd_I_n2421 ;
    wire rd_I_n2420 ;
    wire rd_I_n2419 ;
    wire rd_I_n2418 ;
    wire rd_I_n2417 ;
    wire rd_I_n2416 ;
    wire rd_I_n2415 ;
    wire rd_I_n2414 ;
    wire rd_I_n2413 ;
    wire rd_I_n2412 ;
    wire rd_I_n2411 ;
    wire rd_I_n2410 ;
    wire rd_I_n2409 ;
    wire rd_I_n2408 ;
    wire rd_I_n2407 ;
    wire rd_I_n2406 ;
    wire rd_I_n2405 ;
    wire rd_I_n2404 ;
    wire rd_I_n2403 ;
    wire rd_I_n2402 ;
    wire rd_I_n2401 ;
    wire rd_I_n2400 ;
    wire rd_I_n2399 ;
    wire rd_I_n2398 ;
    wire rd_I_n2397 ;
    wire rd_I_n2396 ;
    wire rd_I_n2395 ;
    wire rd_I_n2394 ;
    wire rd_I_n2393 ;
    wire rd_I_n2392 ;
    wire rd_I_n2391 ;
    wire rd_I_n2390 ;
    wire rd_I_n2389 ;
    wire rd_I_n2388 ;
    wire rd_I_n2387 ;
    wire rd_I_n2386 ;
    wire rd_I_n2385 ;
    wire rd_I_n2384 ;
    wire rd_I_n2383 ;
    wire rd_I_n2382 ;
    wire rd_I_n2381 ;
    wire rd_I_n2380 ;
    wire rd_I_n2379 ;
    wire rd_I_n2378 ;
    wire rd_I_n2377 ;
    wire rd_I_n2376 ;
    wire rd_I_n2375 ;
    wire rd_I_n2374 ;
    wire rd_I_n2373 ;
    wire rd_I_n2372 ;
    wire rd_I_n2371 ;
    wire rd_I_n2370 ;
    wire rd_I_n2369 ;
    wire rd_I_n2368 ;
    wire rd_I_n2367 ;
    wire rd_I_n2366 ;
    wire rd_I_n2365 ;
    wire rd_I_n2364 ;
    wire rd_I_n2363 ;
    wire rd_I_n2362 ;
    wire rd_I_n2361 ;
    wire rd_I_n2360 ;
    wire rd_I_n2359 ;
    wire rd_I_n2358 ;
    wire rd_I_n2357 ;
    wire rd_I_n2356 ;
    wire rd_I_n2355 ;
    wire rd_I_n2354 ;
    wire rd_I_n2353 ;
    wire rd_I_n2352 ;
    wire rd_I_n2351 ;
    wire rd_I_n2350 ;
    wire rd_I_n2349 ;
    wire rd_I_n2348 ;
    wire rd_I_n2347 ;
    wire rd_I_n2346 ;
    wire rd_I_n2345 ;
    wire rd_I_n2344 ;
    wire rd_I_n2343 ;
    wire rd_I_n2342 ;
    wire rd_I_n2341 ;
    wire rd_I_n2340 ;
    wire rd_I_n2339 ;
    wire rd_I_n2338 ;
    wire rd_I_n2337 ;
    wire rd_I_n2336 ;
    wire rd_I_n2335 ;
    wire rd_I_n2334 ;
    wire rd_I_n2333 ;
    wire rd_I_n2332 ;
    wire rd_I_n2331 ;
    wire rd_I_n2330 ;
    wire rd_I_n2329 ;
    wire rd_I_n2328 ;
    wire rd_I_n2327 ;
    wire rd_I_n2326 ;
    wire rd_I_n2325 ;
    wire rd_I_n2324 ;
    wire rd_I_n2323 ;
    wire rd_I_n2322 ;
    wire rd_I_n2321 ;
    wire rd_I_n2320 ;
    wire rd_I_n2319 ;
    wire rd_I_n2318 ;
    wire rd_I_n2317 ;
    wire rd_I_n2316 ;
    wire rd_I_n2315 ;
    wire rd_I_n2314 ;
    wire rd_I_n2313 ;
    wire rd_I_n2312 ;
    wire rd_I_n2311 ;
    wire rd_I_n2310 ;
    wire rd_I_n2309 ;
    wire rd_I_n2308 ;
    wire rd_I_n2307 ;
    wire rd_I_n2306 ;
    wire rd_I_n2305 ;
    wire rd_I_n2304 ;
    wire rd_I_n2303 ;
    wire rd_I_n2302 ;
    wire rd_I_n2301 ;
    wire rd_I_n2300 ;
    wire rd_I_n2299 ;
    wire rd_I_n2298 ;
    wire rd_I_n2297 ;
    wire rd_I_n2296 ;
    wire rd_I_n2295 ;
    wire rd_I_n2294 ;
    wire rd_I_n2293 ;
    wire rd_I_n2292 ;
    wire rd_I_n2291 ;
    wire rd_I_n2290 ;
    wire rd_I_n2289 ;
    wire rd_I_n2288 ;
    wire rd_I_n2287 ;
    wire rd_I_n2286 ;
    wire rd_I_n2285 ;
    wire rd_I_n2284 ;
    wire rd_I_n2283 ;
    wire rd_I_n2282 ;
    wire rd_I_n2281 ;
    wire rd_I_n2280 ;
    wire rd_I_n2279 ;
    wire rd_I_n2278 ;
    wire rd_I_n2277 ;
    wire rd_I_n2276 ;
    wire rd_I_n2275 ;
    wire rd_I_n2274 ;
    wire rd_I_n2273 ;
    wire rd_I_n2272 ;
    wire rd_I_n2271 ;
    wire rd_I_n2270 ;
    wire rd_I_n2269 ;
    wire rd_I_n2268 ;
    wire rd_I_n2267 ;
    wire rd_I_n2266 ;
    wire rd_I_n2265 ;
    wire rd_I_n2264 ;
    wire rd_I_n2263 ;
    wire rd_I_n2262 ;
    wire rd_I_n2261 ;
    wire rd_I_n2260 ;
    wire rd_I_n2259 ;
    wire rd_I_n2258 ;
    wire rd_I_n2257 ;
    wire rd_I_n2256 ;
    wire rd_I_n2255 ;
    wire rd_I_n2254 ;
    wire rd_I_n2253 ;
    wire rd_I_n2252 ;
    wire rd_I_n2251 ;
    wire rd_I_n2250 ;
    wire rd_I_n2249 ;
    wire rd_I_n2248 ;
    wire rd_I_n2247 ;
    wire rd_I_n2246 ;
    wire rd_I_n2245 ;
    wire rd_I_n2244 ;
    wire rd_I_n2243 ;
    wire rd_I_n2242 ;
    wire rd_I_n2241 ;
    wire rd_I_n2240 ;
    wire rd_I_n2239 ;
    wire rd_I_n2238 ;
    wire rd_I_n2237 ;
    wire rd_I_n2236 ;
    wire rd_I_n2235 ;
    wire rd_I_n2234 ;
    wire rd_I_n2233 ;
    wire rd_I_n2232 ;
    wire rd_I_n2231 ;
    wire rd_I_n2230 ;
    wire rd_I_n2229 ;
    wire rd_I_n2228 ;
    wire rd_I_n2227 ;
    wire rd_I_n2226 ;
    wire rd_I_n2225 ;
    wire rd_I_n2224 ;
    wire rd_I_n2223 ;
    wire rd_I_n2222 ;
    wire rd_I_n2221 ;
    wire rd_I_n2220 ;
    wire rd_I_n2219 ;
    wire rd_I_n2218 ;
    wire rd_I_n2217 ;
    wire rd_I_n2216 ;
    wire rd_I_n2215 ;
    wire rd_I_n2214 ;
    wire rd_I_n2213 ;
    wire rd_I_n2212 ;
    wire rd_I_n2211 ;
    wire rd_I_n2210 ;
    wire rd_I_n2209 ;
    wire rd_I_n2208 ;
    wire rd_I_n2207 ;
    wire rd_I_n2206 ;
    wire rd_I_n2205 ;
    wire rd_I_n2204 ;
    wire rd_I_n2203 ;
    wire rd_I_n2202 ;
    wire rd_I_n2201 ;
    wire rd_I_n2200 ;
    wire rd_I_n2199 ;
    wire rd_I_n2198 ;
    wire rd_I_n2197 ;
    wire rd_I_n2196 ;
    wire rd_I_n2195 ;
    wire rd_I_n2194 ;
    wire rd_I_n2193 ;
    wire rd_I_n2192 ;
    wire rd_I_n2191 ;
    wire rd_I_n2190 ;
    wire rd_I_n2189 ;
    wire rd_I_n2188 ;
    wire rd_I_n2187 ;
    wire rd_I_n2186 ;
    wire rd_I_n2185 ;
    wire rd_I_n2184 ;
    wire rd_I_n2183 ;
    wire rd_I_n2182 ;
    wire rd_I_n2181 ;
    wire rd_I_n2180 ;
    wire rd_I_n2179 ;
    wire rd_I_n2178 ;
    wire rd_I_n2177 ;
    wire rd_I_n2176 ;
    wire rd_I_n2175 ;
    wire rd_I_n2174 ;
    wire rd_I_n2173 ;
    wire rd_I_n2172 ;
    wire rd_I_n2171 ;
    wire rd_I_n2170 ;
    wire rd_I_n2169 ;
    wire rd_I_n2168 ;
    wire rd_I_n2167 ;
    wire rd_I_n2166 ;
    wire rd_I_n2165 ;
    wire rd_I_n2164 ;
    wire rd_I_n2163 ;
    wire rd_I_n2162 ;
    wire rd_I_n2161 ;
    wire rd_I_n2160 ;
    wire rd_I_n2159 ;
    wire rd_I_n2158 ;
    wire rd_I_n2157 ;
    wire rd_I_n2156 ;
    wire rd_I_n2155 ;
    wire rd_I_n2154 ;
    wire rd_I_n2153 ;
    wire rd_I_n2152 ;
    wire rd_I_n2151 ;
    wire rd_I_n2150 ;
    wire rd_I_n2149 ;
    wire rd_I_n2148 ;
    wire rd_I_n2147 ;
    wire rd_I_n2146 ;
    wire rd_I_n2145 ;
    wire rd_I_n2144 ;
    wire rd_I_n2143 ;
    wire rd_I_n2142 ;
    wire rd_I_n2141 ;
    wire rd_I_n2140 ;
    wire rd_I_n2139 ;
    wire rd_I_n2138 ;
    wire rd_I_n2137 ;
    wire rd_I_n2136 ;
    wire rd_I_n2135 ;
    wire rd_I_n2134 ;
    wire rd_I_n2133 ;
    wire rd_I_n2132 ;
    wire rd_I_n2131 ;
    wire rd_I_n2130 ;
    wire rd_I_n2129 ;
    wire rd_I_n2128 ;
    wire rd_I_n2127 ;
    wire rd_I_n2126 ;
    wire rd_I_n2125 ;
    wire rd_I_n2124 ;
    wire rd_I_n2123 ;
    wire rd_I_n2122 ;
    wire rd_I_n2121 ;
    wire rd_I_n2120 ;
    wire rd_I_n2119 ;
    wire rd_I_n2118 ;
    wire rd_I_n2117 ;
    wire rd_I_n2116 ;
    wire rd_I_n2115 ;
    wire rd_I_n2114 ;
    wire rd_I_n2113 ;
    wire rd_I_n2112 ;
    wire rd_I_n2111 ;
    wire rd_I_n2110 ;
    wire rd_I_n2109 ;
    wire rd_I_n2108 ;
    wire rd_I_n2107 ;
    wire rd_I_n2106 ;
    wire rd_I_n2105 ;
    wire rd_I_n2104 ;
    wire rd_I_n2103 ;
    wire rd_I_n2102 ;
    wire rd_I_n2101 ;
    wire rd_I_n2100 ;
    wire rd_I_n2099 ;
    wire rd_I_n2098 ;
    wire rd_I_n2097 ;
    wire rd_I_n2096 ;
    wire rd_I_n2095 ;
    wire rd_I_n2094 ;
    wire rd_I_n2093 ;
    wire rd_I_n2092 ;
    wire rd_I_n2091 ;
    wire rd_I_n2090 ;
    wire rd_I_n2089 ;
    wire rd_I_n2088 ;
    wire rd_I_n2087 ;
    wire rd_I_n2086 ;
    wire rd_I_n2085 ;
    wire rd_I_n2084 ;
    wire rd_I_n2083 ;
    wire rd_I_n2082 ;
    wire rd_I_n2081 ;
    wire rd_I_n2080 ;
    wire rd_I_n2079 ;
    wire rd_I_n2078 ;
    wire rd_I_n2077 ;
    wire rd_I_n2076 ;
    wire rd_I_n2075 ;
    wire rd_I_n2074 ;
    wire rd_I_n2073 ;
    wire rd_I_n2072 ;
    wire rd_I_n2071 ;
    wire rd_I_n2070 ;
    wire rd_I_n2069 ;
    wire rd_I_n2068 ;
    wire rd_I_n2067 ;
    wire rd_I_n2066 ;
    wire rd_I_n2065 ;
    wire rd_I_n2064 ;
    wire rd_I_n2063 ;
    wire rd_I_n2062 ;
    wire rd_I_n2061 ;
    wire rd_I_n2060 ;
    wire rd_I_n2059 ;
    wire rd_I_n2058 ;
    wire rd_I_n2057 ;
    wire rd_I_n2056 ;
    wire rd_I_n2055 ;
    wire rd_I_n2054 ;
    wire rd_I_n2053 ;
    wire rd_I_n2052 ;
    wire rd_I_n2051 ;
    wire rd_I_n2050 ;
    wire rd_I_n2049 ;
    wire rd_I_n2048 ;
    wire rd_I_n2047 ;
    wire rd_I_n2046 ;
    wire rd_I_n2045 ;
    wire rd_I_n2044 ;
    wire rd_I_n2043 ;
    wire rd_I_n2042 ;
    wire rd_I_n2041 ;
    wire rd_I_n2040 ;
    wire rd_I_n2039 ;
    wire rd_I_n2038 ;
    wire rd_I_n2037 ;
    wire rd_I_n2036 ;
    wire rd_I_n2035 ;
    wire rd_I_n2034 ;
    wire rd_I_n2033 ;
    wire rd_I_n2032 ;
    wire rd_I_n2031 ;
    wire rd_I_n2030 ;
    wire rd_I_n2029 ;
    wire rd_I_n2028 ;
    wire rd_I_n2027 ;
    wire rd_I_n2026 ;
    wire rd_I_n2025 ;
    wire rd_I_n2024 ;
    wire rd_I_n2023 ;
    wire rd_I_n2022 ;
    wire rd_I_n2021 ;
    wire rd_I_n2020 ;
    wire rd_I_n2019 ;
    wire rd_I_n2018 ;
    wire rd_I_n2017 ;
    wire rd_I_n2016 ;
    wire rd_I_n2015 ;
    wire rd_I_n2014 ;
    wire rd_I_n2013 ;
    wire rd_I_n2012 ;
    wire rd_I_n2011 ;
    wire rd_I_n2010 ;
    wire rd_I_n2009 ;
    wire rd_I_n2008 ;
    wire rd_I_n2007 ;
    wire rd_I_n2006 ;
    wire rd_I_n2005 ;
    wire rd_I_n2004 ;
    wire rd_I_n2003 ;
    wire rd_I_n2002 ;
    wire rd_I_n2001 ;
    wire rd_I_n2000 ;
    wire rd_I_n1999 ;
    wire rd_I_n1998 ;
    wire rd_I_n1997 ;
    wire rd_I_n1996 ;
    wire rd_I_n1995 ;
    wire rd_I_n1994 ;
    wire rd_I_n1993 ;
    wire rd_I_n1992 ;
    wire rd_I_n1991 ;
    wire rd_I_n1990 ;
    wire rd_I_n1989 ;
    wire rd_I_n1988 ;
    wire rd_I_n1987 ;
    wire rd_I_n1986 ;
    wire rd_I_n1985 ;
    wire rd_I_n1984 ;
    wire rd_I_n1983 ;
    wire rd_I_n1982 ;
    wire rd_I_n1981 ;
    wire rd_I_n1980 ;
    wire rd_I_n1979 ;
    wire rd_I_n1978 ;
    wire rd_I_n1977 ;
    wire rd_I_n1976 ;
    wire rd_I_n1975 ;
    wire rd_I_n1974 ;
    wire rd_I_n1973 ;
    wire rd_I_n1972 ;
    wire rd_I_n1971 ;
    wire rd_I_n1970 ;
    wire rd_I_n1969 ;
    wire rd_I_n1968 ;
    wire rd_I_n1967 ;
    wire rd_I_n1966 ;
    wire rd_I_n1965 ;
    wire rd_I_n1964 ;
    wire rd_I_n1963 ;
    wire rd_I_n1962 ;
    wire rd_I_n1961 ;
    wire rd_I_n1960 ;
    wire rd_I_n1959 ;
    wire rd_I_n1958 ;
    wire rd_I_n1957 ;
    wire rd_I_n1956 ;
    wire rd_I_n1955 ;
    wire rd_I_n1954 ;
    wire rd_I_n1953 ;
    wire rd_I_n1952 ;
    wire rd_I_n1951 ;
    wire rd_I_n1950 ;
    wire rd_I_n1949 ;
    wire rd_I_n1948 ;
    wire rd_I_n1947 ;
    wire rd_I_n1946 ;
    wire rd_I_n1945 ;
    wire rd_I_n1944 ;
    wire rd_I_n1943 ;
    wire rd_I_n1942 ;
    wire rd_I_n1941 ;
    wire rd_I_n1940 ;
    wire rd_I_n1939 ;
    wire rd_I_n1938 ;
    wire rd_I_n1937 ;
    wire rd_I_n1936 ;
    wire rd_I_n1935 ;
    wire rd_I_n1934 ;
    wire rd_I_n1933 ;
    wire rd_I_n1932 ;
    wire rd_I_n1931 ;
    wire rd_I_n1930 ;
    wire rd_I_n1929 ;
    wire rd_I_n1928 ;
    wire rd_I_n1927 ;
    wire rd_I_n1926 ;
    wire rd_I_n1925 ;
    wire rd_I_n1924 ;
    wire rd_I_n1923 ;
    wire rd_I_n1922 ;
    wire rd_I_n1921 ;
    wire rd_I_n1920 ;
    wire rd_I_n1919 ;
    wire rd_I_n1918 ;
    wire rd_I_n1917 ;
    wire rd_I_n1916 ;
    wire rd_I_n1915 ;
    wire rd_I_n1914 ;
    wire rd_I_n1913 ;
    wire rd_I_n1912 ;
    wire rd_I_n1911 ;
    wire rd_I_n1910 ;
    wire rd_I_n1909 ;
    wire rd_I_n1908 ;
    wire rd_I_n1907 ;
    wire rd_I_n1906 ;
    wire rd_I_n1905 ;
    wire rd_I_n1904 ;
    wire rd_I_n1903 ;
    wire rd_I_n1902 ;
    wire rd_I_n1901 ;
    wire rd_I_n1900 ;
    wire rd_I_n1899 ;
    wire rd_I_n1898 ;
    wire rd_I_n1897 ;
    wire rd_I_n1896 ;
    wire rd_I_n1895 ;
    wire rd_I_n1894 ;
    wire rd_I_n1893 ;
    wire rd_I_n1892 ;
    wire rd_I_n1891 ;
    wire rd_I_n1890 ;
    wire rd_I_n1889 ;
    wire rd_I_n1888 ;
    wire rd_I_n1887 ;
    wire rd_I_n1886 ;
    wire rd_I_n1885 ;
    wire rd_I_n1884 ;
    wire rd_I_n1883 ;
    wire rd_I_n1882 ;
    wire rd_I_n1881 ;
    wire rd_I_n1880 ;
    wire rd_I_n1879 ;
    wire rd_I_n1878 ;
    wire rd_I_n1877 ;
    wire rd_I_n1876 ;
    wire rd_I_n1875 ;
    wire rd_I_n1874 ;
    wire rd_I_n1873 ;
    wire rd_I_n1872 ;
    wire rd_I_n1871 ;
    wire rd_I_n1870 ;
    wire rd_I_n1869 ;
    wire rd_I_n1868 ;
    wire rd_I_n1867 ;
    wire rd_I_n1866 ;
    wire rd_I_n1865 ;
    wire rd_I_n1864 ;
    wire rd_I_n1863 ;
    wire rd_I_n1862 ;
    wire rd_I_n1861 ;
    wire rd_I_n1860 ;
    wire rd_I_n1859 ;
    wire rd_I_n1858 ;
    wire rd_I_n1857 ;
    wire rd_I_n1856 ;
    wire rd_I_n1855 ;
    wire rd_I_n1854 ;
    wire rd_I_n1853 ;
    wire rd_I_n1852 ;
    wire rd_I_n1851 ;
    wire rd_I_n1850 ;
    wire rd_I_n1849 ;
    wire rd_I_n1848 ;
    wire rd_I_n1847 ;
    wire rd_I_n1846 ;
    wire rd_I_n1845 ;
    wire rd_I_n1844 ;
    wire rd_I_n1843 ;
    wire rd_I_n1842 ;
    wire rd_I_n1841 ;
    wire rd_I_n1840 ;
    wire rd_I_n1839 ;
    wire rd_I_n1838 ;
    wire rd_I_n1837 ;
    wire rd_I_n1836 ;
    wire rd_I_n1835 ;
    wire rd_I_n1834 ;
    wire rd_I_n1833 ;
    wire rd_I_n1832 ;
    wire rd_I_n1831 ;
    wire rd_I_n1830 ;
    wire rd_I_n1829 ;
    wire rd_I_n1828 ;
    wire rd_I_n1827 ;
    wire rd_I_n1826 ;
    wire rd_I_n1825 ;
    wire rd_I_n1824 ;
    wire rd_I_n1823 ;
    wire rd_I_n1822 ;
    wire rd_I_n1821 ;
    wire rd_I_n1820 ;
    wire rd_I_n1819 ;
    wire rd_I_n1818 ;
    wire rd_I_n1817 ;
    wire rd_I_n1816 ;
    wire rd_I_n1815 ;
    wire rd_I_n1814 ;
    wire rd_I_n1813 ;
    wire rd_I_n1812 ;
    wire rd_I_n1811 ;
    wire rd_I_n1810 ;
    wire rd_I_n1809 ;
    wire rd_I_n1808 ;
    wire rd_I_n1807 ;
    wire rd_I_n1806 ;
    wire rd_I_n1805 ;
    wire rd_I_n1804 ;
    wire rd_I_n1803 ;
    wire rd_I_n1802 ;
    wire rd_I_n1801 ;
    wire rd_I_n1800 ;
    wire rd_I_n1799 ;
    wire rd_I_n1798 ;
    wire rd_I_n1797 ;
    wire rd_I_n1796 ;
    wire rd_I_n1795 ;
    wire rd_I_n1794 ;
    wire rd_I_n1793 ;
    wire rd_I_n1792 ;
    wire rd_I_n1791 ;
    wire rd_I_n1790 ;
    wire rd_I_n1789 ;
    wire rd_I_n1788 ;
    wire rd_I_n1787 ;
    wire rd_I_n1786 ;
    wire rd_I_n1785 ;
    wire rd_I_n1784 ;
    wire rd_I_n1783 ;
    wire rd_I_n1782 ;
    wire rd_I_n1781 ;
    wire rd_I_n1780 ;
    wire rd_I_n1779 ;
    wire rd_I_n1778 ;
    wire rd_I_n1777 ;
    wire rd_I_n1776 ;
    wire rd_I_n1775 ;
    wire rd_I_n1774 ;
    wire rd_I_n1773 ;
    wire rd_I_n1772 ;
    wire rd_I_n1771 ;
    wire rd_I_n1770 ;
    wire rd_I_n1769 ;
    wire rd_I_n1768 ;
    wire rd_I_n1767 ;
    wire rd_I_n1766 ;
    wire rd_I_n1765 ;
    wire rd_I_n1764 ;
    wire rd_I_n1763 ;
    wire rd_I_n1762 ;
    wire rd_I_n1761 ;
    wire rd_I_n1760 ;
    wire rd_I_n1759 ;
    wire rd_I_n1758 ;
    wire rd_I_n1757 ;
    wire rd_I_n1756 ;
    wire rd_I_n1755 ;
    wire rd_I_n1754 ;
    wire rd_I_n1753 ;
    wire rd_I_n1752 ;
    wire rd_I_n1751 ;
    wire rd_I_n1750 ;
    wire rd_I_n1749 ;
    wire rd_I_n1748 ;
    wire rd_I_n1747 ;
    wire rd_I_n1746 ;
    wire rd_I_n1745 ;
    wire rd_I_n1744 ;
    wire rd_I_n1743 ;
    wire rd_I_n1742 ;
    wire rd_I_n1741 ;
    wire rd_I_n1740 ;
    wire rd_I_n1739 ;
    wire rd_I_n1738 ;
    wire rd_I_n1737 ;
    wire rd_I_n1736 ;
    wire rd_I_n1735 ;
    wire rd_I_n1734 ;
    wire rd_I_n1733 ;
    wire rd_I_n1732 ;
    wire rd_I_n1731 ;
    wire rd_I_n1730 ;
    wire rd_I_n1729 ;
    wire rd_I_n1728 ;
    wire rd_I_n1727 ;
    wire rd_I_n1726 ;
    wire rd_I_n1725 ;
    wire rd_I_n1724 ;
    wire rd_I_n1723 ;
    wire rd_I_n1722 ;
    wire rd_I_n1721 ;
    wire rd_I_n1720 ;
    wire rd_I_n1719 ;
    wire rd_I_n1718 ;
    wire rd_I_n1717 ;
    wire rd_I_n1716 ;
    wire rd_I_n1715 ;
    wire rd_I_n1714 ;
    wire rd_I_n1713 ;
    wire rd_I_n1712 ;
    wire rd_I_n1711 ;
    wire rd_I_n1710 ;
    wire rd_I_n1709 ;
    wire rd_I_n1708 ;
    wire rd_I_n1707 ;
    wire rd_I_n1706 ;
    wire rd_I_n1705 ;
    wire rd_I_n1704 ;
    wire rd_I_n1703 ;
    wire rd_I_n1702 ;
    wire rd_I_n1701 ;
    wire rd_I_n1700 ;
    wire rd_I_n1699 ;
    wire rd_I_n1698 ;
    wire rd_I_n1697 ;
    wire rd_I_n1696 ;
    wire rd_I_n1695 ;
    wire rd_I_n1694 ;
    wire rd_I_n1693 ;
    wire rd_I_n1692 ;
    wire rd_I_n1691 ;
    wire rd_I_n1690 ;
    wire rd_I_n1689 ;
    wire rd_I_n1688 ;
    wire rd_I_n1687 ;
    wire rd_I_n1686 ;
    wire rd_I_n1685 ;
    wire rd_I_n1684 ;
    wire rd_I_n1683 ;
    wire rd_I_n1682 ;
    wire rd_I_n1681 ;
    wire rd_I_n1680 ;
    wire rd_I_n1679 ;
    wire rd_I_n1678 ;
    wire rd_I_n1677 ;
    wire rd_I_n1676 ;
    wire rd_I_n1675 ;
    wire rd_I_n1674 ;
    wire rd_I_n1673 ;
    wire rd_I_n1672 ;
    wire rd_I_n1671 ;
    wire rd_I_n1670 ;
    wire rd_I_n1669 ;
    wire rd_I_n1668 ;
    wire rd_I_n1667 ;
    wire rd_I_n1666 ;
    wire rd_I_n1665 ;
    wire rd_I_n1664 ;
    wire rd_I_n1663 ;
    wire rd_I_n1662 ;
    wire rd_I_n1661 ;
    wire rd_I_n1660 ;
    wire rd_I_n1659 ;
    wire rd_I_n1658 ;
    wire rd_I_n1657 ;
    wire rd_I_n1656 ;
    wire rd_I_n1655 ;
    wire rd_I_n1654 ;
    wire rd_I_n1653 ;
    wire rd_I_n1652 ;
    wire rd_I_n1651 ;
    wire rd_I_n1650 ;
    wire rd_I_n1649 ;
    wire rd_I_n1648 ;
    wire rd_I_n1647 ;
    wire rd_I_n1646 ;
    wire rd_I_n1645 ;
    wire rd_I_n1644 ;
    wire rd_I_n1643 ;
    wire rd_I_n1642 ;
    wire rd_I_n1641 ;
    wire rd_I_n1640 ;
    wire rd_I_n1639 ;
    wire rd_I_n1638 ;
    wire rd_I_n1637 ;
    wire rd_I_n1636 ;
    wire rd_I_n1635 ;
    wire rd_I_n1634 ;
    wire rd_I_n1633 ;
    wire rd_I_n1632 ;
    wire rd_I_n1631 ;
    wire rd_I_n1630 ;
    wire rd_I_n1629 ;
    wire rd_I_n1628 ;
    wire rd_I_n1627 ;
    wire rd_I_n1626 ;
    wire rd_I_n1625 ;
    wire rd_I_n1624 ;
    wire rd_I_n1623 ;
    wire rd_I_n1622 ;
    wire rd_I_n1621 ;
    wire rd_I_n1620 ;
    wire rd_I_n1619 ;
    wire rd_I_n1618 ;
    wire rd_I_n1617 ;
    wire rd_I_n1616 ;
    wire rd_I_n1615 ;
    wire rd_I_n1614 ;
    wire rd_I_n1613 ;
    wire rd_I_n1612 ;
    wire rd_I_n1611 ;
    wire rd_I_n1610 ;
    wire rd_I_n1609 ;
    wire rd_I_n1608 ;
    wire rd_I_n1607 ;
    wire rd_I_n1606 ;
    wire rd_I_n1605 ;
    wire rd_I_n1604 ;
    wire rd_I_n1603 ;
    wire rd_I_n1602 ;
    wire rd_I_n1601 ;
    wire rd_I_n1600 ;
    wire rd_I_n1599 ;
    wire rd_I_n1598 ;
    wire rd_I_n1597 ;
    wire rd_I_n1596 ;
    wire rd_I_n1595 ;
    wire rd_I_n1594 ;
    wire rd_I_n1593 ;
    wire rd_I_n1592 ;
    wire rd_I_n1591 ;
    wire rd_I_n1590 ;
    wire rd_I_n1589 ;
    wire rd_I_n1588 ;
    wire rd_I_n1587 ;
    wire rd_I_n1586 ;
    wire rd_I_n1585 ;
    wire rd_I_n1584 ;
    wire rd_I_n1583 ;
    wire rd_I_n1582 ;
    wire rd_I_n1581 ;
    wire rd_I_n1580 ;
    wire rd_I_n1579 ;
    wire rd_I_n1578 ;
    wire rd_I_n1577 ;
    wire rd_I_n1576 ;
    wire rd_I_n1575 ;
    wire rd_I_n1574 ;
    wire rd_I_n1573 ;
    wire rd_I_n1572 ;
    wire rd_I_n1571 ;
    wire rd_I_n1570 ;
    wire rd_I_n1569 ;
    wire rd_I_n1568 ;
    wire rd_I_n1567 ;
    wire rd_I_n1566 ;
    wire rd_I_n1565 ;
    wire rd_I_n1564 ;
    wire rd_I_n1563 ;
    wire rd_I_n1562 ;
    wire rd_I_n1561 ;
    wire rd_I_n1560 ;
    wire rd_I_n1559 ;
    wire rd_I_n1558 ;
    wire rd_I_n1557 ;
    wire rd_I_n1556 ;
    wire rd_I_n1555 ;
    wire rd_I_n1554 ;
    wire rd_I_n1553 ;
    wire rd_I_n1552 ;
    wire rd_I_n1551 ;
    wire rd_I_n1550 ;
    wire rd_I_n1549 ;
    wire rd_I_n1548 ;
    wire rd_I_n1547 ;
    wire rd_I_n1546 ;
    wire rd_I_n1545 ;
    wire rd_I_n1544 ;
    wire rd_I_n1543 ;
    wire rd_I_n1542 ;
    wire rd_I_n1541 ;
    wire rd_I_n1540 ;
    wire rd_I_n1539 ;
    wire rd_I_n1538 ;
    wire rd_I_n1537 ;
    wire rd_I_n1536 ;
    wire rd_I_n1535 ;
    wire rd_I_n1534 ;
    wire rd_I_n1533 ;
    wire rd_I_n1532 ;
    wire rd_I_n1531 ;
    wire rd_I_n1530 ;
    wire rd_I_n1529 ;
    wire rd_I_n1528 ;
    wire rd_I_n1527 ;
    wire rd_I_n1526 ;
    wire rd_I_n1525 ;
    wire rd_I_n1524 ;
    wire rd_I_n1523 ;
    wire rd_I_n1522 ;
    wire rd_I_n1521 ;
    wire rd_I_n1520 ;
    wire rd_I_n1519 ;
    wire rd_I_n1518 ;
    wire rd_I_n1517 ;
    wire rd_I_n1516 ;
    wire rd_I_n1515 ;
    wire rd_I_n1514 ;
    wire rd_I_n1513 ;
    wire rd_I_n1512 ;
    wire rd_I_n1511 ;
    wire rd_I_n1510 ;
    wire rd_I_n1509 ;
    wire rd_I_n1508 ;
    wire rd_I_n1507 ;
    wire rd_I_n1506 ;
    wire rd_I_n1505 ;
    wire rd_I_n1504 ;
    wire rd_I_n1503 ;
    wire rd_I_n1502 ;
    wire rd_I_n1501 ;
    wire rd_I_n1500 ;
    wire rd_I_n1499 ;
    wire rd_I_n1498 ;
    wire rd_I_n1497 ;
    wire rd_I_n1496 ;
    wire rd_I_n1495 ;
    wire rd_I_n1494 ;
    wire rd_I_n1493 ;
    wire rd_I_n1492 ;
    wire rd_I_n1491 ;
    wire rd_I_n1490 ;
    wire rd_I_n1489 ;
    wire rd_I_n1488 ;
    wire rd_I_n1487 ;
    wire rd_I_n1486 ;
    wire rd_I_n1485 ;
    wire rd_I_n1484 ;
    wire rd_I_n1483 ;
    wire rd_I_n1482 ;
    wire rd_I_n1481 ;
    wire rd_I_n1480 ;
    wire rd_I_n1479 ;
    wire rd_I_n1478 ;
    wire rd_I_n1477 ;
    wire rd_I_n1476 ;
    wire rd_I_n1475 ;
    wire rd_I_n1474 ;
    wire rd_I_n1473 ;
    wire rd_I_n1472 ;
    wire rd_I_n1471 ;
    wire rd_I_n1470 ;
    wire rd_I_n1469 ;
    wire rd_I_n1468 ;
    wire rd_I_n1467 ;
    wire rd_I_n1466 ;
    wire rd_I_n1465 ;
    wire rd_I_n1464 ;
    wire rd_I_n1463 ;
    wire rd_I_n1462 ;
    wire rd_I_n1461 ;
    wire rd_I_n1460 ;
    wire rd_I_n1459 ;
    wire rd_I_n1458 ;
    wire rd_I_n1457 ;
    wire rd_I_n1456 ;
    wire rd_I_n1455 ;
    wire rd_I_n1454 ;
    wire rd_I_n1453 ;
    wire rd_I_n1452 ;
    wire rd_I_n1451 ;
    wire rd_I_n1450 ;
    wire rd_I_n1449 ;
    wire rd_I_n1448 ;
    wire rd_I_n1447 ;
    wire rd_I_n1446 ;
    wire rd_I_n1445 ;
    wire rd_I_n1444 ;
    wire rd_I_n1443 ;
    wire rd_I_n1442 ;
    wire rd_I_n1441 ;
    wire rd_I_n1440 ;
    wire rd_I_n1439 ;
    wire rd_I_n1438 ;
    wire rd_I_n1437 ;
    wire rd_I_n1436 ;
    wire rd_I_n1435 ;
    wire rd_I_n1434 ;
    wire rd_I_n1433 ;
    wire rd_I_n1432 ;
    wire rd_I_n1431 ;
    wire rd_I_n1430 ;
    wire rd_I_n1429 ;
    wire rd_I_n1428 ;
    wire rd_I_n1427 ;
    wire rd_I_n1426 ;
    wire rd_I_n1425 ;
    wire rd_I_n1424 ;
    wire rd_I_n1423 ;
    wire rd_I_n1422 ;
    wire rd_I_n1421 ;
    wire rd_I_n1420 ;
    wire rd_I_n1419 ;
    wire rd_I_n1418 ;
    wire rd_I_n1417 ;
    wire rd_I_n1416 ;
    wire rd_I_n1415 ;
    wire rd_I_n1414 ;
    wire rd_I_n1413 ;
    wire rd_I_n1412 ;
    wire rd_I_n1411 ;
    wire rd_I_n1410 ;
    wire rd_I_n1409 ;
    wire rd_I_n1408 ;
    wire rd_I_n1407 ;
    wire rd_I_n1406 ;
    wire rd_I_n1405 ;
    wire rd_I_n1404 ;
    wire rd_I_n1403 ;
    wire rd_I_n1402 ;
    wire rd_I_n1401 ;
    wire rd_I_n1400 ;
    wire rd_I_n1399 ;
    wire rd_I_n1398 ;
    wire rd_I_n1397 ;
    wire rd_I_n1396 ;
    wire rd_I_n1395 ;
    wire rd_I_n1394 ;
    wire rd_I_n1393 ;
    wire rd_I_n1392 ;
    wire rd_I_n1391 ;
    wire rd_I_n1390 ;
    wire rd_I_n1389 ;
    wire rd_I_n1388 ;
    wire rd_I_n1387 ;
    wire rd_I_n1386 ;
    wire rd_I_n1385 ;
    wire rd_I_n1384 ;
    wire rd_I_n1383 ;
    wire rd_I_n1382 ;
    wire rd_I_n1381 ;
    wire rd_I_n1380 ;
    wire rd_I_n1379 ;
    wire rd_I_n1378 ;
    wire rd_I_n1377 ;
    wire rd_I_n1376 ;
    wire rd_I_n1375 ;
    wire rd_I_n1374 ;
    wire rd_I_n1373 ;
    wire rd_I_n1372 ;
    wire rd_I_n1371 ;
    wire rd_I_n1370 ;
    wire rd_I_n1369 ;
    wire rd_I_n1368 ;
    wire rd_I_n1367 ;
    wire rd_I_n1366 ;
    wire rd_I_n1365 ;
    wire rd_I_n1364 ;
    wire rd_I_n1363 ;
    wire rd_I_n1362 ;
    wire rd_I_n1361 ;
    wire rd_I_n1360 ;
    wire rd_I_n1359 ;
    wire rd_I_n1358 ;
    wire rd_I_n1357 ;
    wire rd_I_n1356 ;
    wire rd_I_n1355 ;
    wire rd_I_n1354 ;
    wire rd_I_n1353 ;
    wire rd_I_n1352 ;
    wire rd_I_n1351 ;
    wire rd_I_n1350 ;
    wire rd_I_n1349 ;
    wire rd_I_n1348 ;
    wire rd_I_n1347 ;
    wire rd_I_n1346 ;
    wire rd_I_n1345 ;
    wire rd_I_n1344 ;
    wire rd_I_n1343 ;
    wire rd_I_n1342 ;
    wire rd_I_n1341 ;
    wire rd_I_n1340 ;
    wire rd_I_n1339 ;
    wire rd_I_n1338 ;
    wire rd_I_n1337 ;
    wire rd_I_n1336 ;
    wire rd_I_n1335 ;
    wire rd_I_n1334 ;
    wire rd_I_n1333 ;
    wire rd_I_n1332 ;
    wire rd_I_n1331 ;
    wire rd_I_n1330 ;
    wire rd_I_n1329 ;
    wire rd_I_n1328 ;
    wire rd_I_n1327 ;
    wire rd_I_n1326 ;
    wire rd_I_n1325 ;
    wire rd_I_n1324 ;
    wire rd_I_n1323 ;
    wire rd_I_n1322 ;
    wire rd_I_n1321 ;
    wire rd_I_n1320 ;
    wire rd_I_n1319 ;
    wire rd_I_n1318 ;
    wire rd_I_n1317 ;
    wire rd_I_n1316 ;
    wire rd_I_n1315 ;
    wire rd_I_n1314 ;
    wire rd_I_n1313 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire clk_gated ;

    /* cells in depth 0 */
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1684 ( .a ({new_AGEMA_signal_4120, new_AGEMA_signal_4119, rd_I_n2600}), .b ({new_AGEMA_signal_4462, new_AGEMA_signal_4461, rd_I_n2602}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1677 ( .a ({new_AGEMA_signal_3690, new_AGEMA_signal_3689, rd_I_n2587}), .b ({new_AGEMA_signal_4468, new_AGEMA_signal_4467, rd_I_n2589}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1670 ( .a ({new_AGEMA_signal_3730, new_AGEMA_signal_3729, rd_I_n2574}), .b ({new_AGEMA_signal_4474, new_AGEMA_signal_4473, rd_I_n2576}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1667 ( .a ({new_AGEMA_signal_3736, new_AGEMA_signal_3735, rd_I_n2569}), .b ({new_AGEMA_signal_4476, new_AGEMA_signal_4475, rd_I_n2571}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1664 ( .a ({new_AGEMA_signal_3874, new_AGEMA_signal_3873, rd_I_n2597}), .b ({new_AGEMA_signal_4478, new_AGEMA_signal_4477, rd_I_n2567}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1661 ( .a ({new_AGEMA_signal_3876, new_AGEMA_signal_3875, rd_I_n2622}), .b ({new_AGEMA_signal_4480, new_AGEMA_signal_4479, rd_I_n2565}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1656 ( .a ({new_AGEMA_signal_4122, new_AGEMA_signal_4121, rd_I_n2556}), .b ({new_AGEMA_signal_4484, new_AGEMA_signal_4483, rd_I_n2558}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1653 ( .a ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, rd_I_n2551}), .b ({new_AGEMA_signal_5240, new_AGEMA_signal_5239, rd_I_n2553}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1650 ( .a ({new_AGEMA_signal_3856, new_AGEMA_signal_3855, rd_I_n2546}), .b ({new_AGEMA_signal_4486, new_AGEMA_signal_4485, rd_I_n2548}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1647 ( .a ({new_AGEMA_signal_4228, new_AGEMA_signal_4227, rd_I_n2541}), .b ({new_AGEMA_signal_4488, new_AGEMA_signal_4487, rd_I_n2543}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1638 ( .a ({new_AGEMA_signal_3778, new_AGEMA_signal_3777, rd_I_n2530}), .b ({new_AGEMA_signal_4496, new_AGEMA_signal_4495, rd_I_n2532}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1631 ( .a ({new_AGEMA_signal_3942, new_AGEMA_signal_3941, rd_I_n2520}), .b ({new_AGEMA_signal_4502, new_AGEMA_signal_4501, rd_I_n2522}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1628 ( .a ({new_AGEMA_signal_3834, new_AGEMA_signal_3833, rd_I_n2515}), .b ({new_AGEMA_signal_4504, new_AGEMA_signal_4503, rd_I_n2517}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1625 ( .a ({new_AGEMA_signal_3840, new_AGEMA_signal_3839, rd_I_n2510}), .b ({new_AGEMA_signal_4506, new_AGEMA_signal_4505, rd_I_n2512}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1622 ( .a ({new_AGEMA_signal_3976, new_AGEMA_signal_3975, rd_I_n2505}), .b ({new_AGEMA_signal_4508, new_AGEMA_signal_4507, rd_I_n2507}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1619 ( .a ({new_AGEMA_signal_3970, new_AGEMA_signal_3969, rd_I_n2500}), .b ({new_AGEMA_signal_4510, new_AGEMA_signal_4509, rd_I_n2502}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1616 ( .a ({new_AGEMA_signal_4408, new_AGEMA_signal_4407, rd_I_n2495}), .b ({new_AGEMA_signal_4512, new_AGEMA_signal_4511, rd_I_n2497}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1613 ( .a ({new_AGEMA_signal_4426, new_AGEMA_signal_4425, rd_I_n2490}), .b ({new_AGEMA_signal_4514, new_AGEMA_signal_4513, rd_I_n2492}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1606 ( .a ({new_AGEMA_signal_4218, new_AGEMA_signal_4217, rd_I_n2477}), .b ({new_AGEMA_signal_4520, new_AGEMA_signal_4519, rd_I_n2479}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1597 ( .a ({new_AGEMA_signal_3706, new_AGEMA_signal_3705, rd_I_n2466}), .b ({new_AGEMA_signal_4528, new_AGEMA_signal_4527, rd_I_n2468}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1594 ( .a ({new_AGEMA_signal_3700, new_AGEMA_signal_3699, rd_I_n2461}), .b ({new_AGEMA_signal_4530, new_AGEMA_signal_4529, rd_I_n2463}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1583 ( .a ({new_AGEMA_signal_3748, new_AGEMA_signal_3747, rd_I_n2610}), .b ({new_AGEMA_signal_4540, new_AGEMA_signal_4539, rd_I_n2443}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1580 ( .a ({new_AGEMA_signal_3688, new_AGEMA_signal_3687, rd_I_n2614}), .b ({new_AGEMA_signal_4542, new_AGEMA_signal_4541, rd_I_n2441}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1577 ( .a ({new_AGEMA_signal_4014, new_AGEMA_signal_4013, rd_I_n2436}), .b ({new_AGEMA_signal_4544, new_AGEMA_signal_4543, rd_I_n2438}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1562 ( .a ({new_AGEMA_signal_4132, new_AGEMA_signal_4131, rd_I_n2410}), .b ({new_AGEMA_signal_4558, new_AGEMA_signal_4557, rd_I_n2412}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1559 ( .a ({new_AGEMA_signal_4390, new_AGEMA_signal_4389, rd_I_n2405}), .b ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, rd_I_n2407}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1556 ( .a ({new_AGEMA_signal_3916, new_AGEMA_signal_3915, rd_I_n2487}), .b ({new_AGEMA_signal_4562, new_AGEMA_signal_4561, rd_I_n2403}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1551 ( .a ({new_AGEMA_signal_4108, new_AGEMA_signal_4107, rd_I_n2394}), .b ({new_AGEMA_signal_4566, new_AGEMA_signal_4565, rd_I_n2396}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1548 ( .a ({new_AGEMA_signal_3988, new_AGEMA_signal_3987, rd_I_n2389}), .b ({new_AGEMA_signal_4568, new_AGEMA_signal_4567, rd_I_n2391}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1545 ( .a ({new_AGEMA_signal_3708, new_AGEMA_signal_3707, rd_I_n2384}), .b ({new_AGEMA_signal_4570, new_AGEMA_signal_4569, rd_I_n2386}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1540 ( .a ({new_AGEMA_signal_4354, new_AGEMA_signal_4353, rd_I_n2375}), .b ({new_AGEMA_signal_4574, new_AGEMA_signal_4573, rd_I_n2377}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1531 ( .a ({new_AGEMA_signal_3754, new_AGEMA_signal_3753, rd_I_n2446}), .b ({new_AGEMA_signal_4582, new_AGEMA_signal_4581, rd_I_n2361}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1526 ( .a ({state_in_s2[40], state_in_s1[40], state_in_s0[40]}), .b ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, rd_I_n2355}), .c ({new_AGEMA_signal_3684, new_AGEMA_signal_3683, rd_I_n2613}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1525 ( .a ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, rd_I_n2354}), .b ({state_in_s2[136], state_in_s1[136], state_in_s0[136]}), .c ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, rd_I_n2616}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1524 ( .a ({state_in_s2[317], state_in_s1[317], state_in_s0[317]}), .b ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, rd_I_n2353}), .c ({new_AGEMA_signal_3688, new_AGEMA_signal_3687, rd_I_n2614}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1521 ( .a ({new_AGEMA_signal_4296, new_AGEMA_signal_4295, rd_I_n2348}), .b ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, rd_I_n2350}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1518 ( .a ({new_AGEMA_signal_4290, new_AGEMA_signal_4289, rd_I_n2343}), .b ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, rd_I_n2345}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1515 ( .a ({new_AGEMA_signal_3808, new_AGEMA_signal_3807, rd_I_n2338}), .b ({new_AGEMA_signal_4592, new_AGEMA_signal_4591, rd_I_n2340}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1512 ( .a ({new_AGEMA_signal_3760, new_AGEMA_signal_3759, rd_I_n2606}), .b ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, rd_I_n2336}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1509 ( .a ({new_AGEMA_signal_4134, new_AGEMA_signal_4133, rd_I_n2400}), .b ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, rd_I_n2334}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1506 ( .a ({new_AGEMA_signal_3892, new_AGEMA_signal_3891, rd_I_n2562}), .b ({new_AGEMA_signal_4598, new_AGEMA_signal_4597, rd_I_n2332}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1503 ( .a ({new_AGEMA_signal_3820, new_AGEMA_signal_3819, rd_I_n2327}), .b ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, rd_I_n2329}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1496 ( .a ({new_AGEMA_signal_4264, new_AGEMA_signal_4263, rd_I_n2314}), .b ({new_AGEMA_signal_4606, new_AGEMA_signal_4605, rd_I_n2316}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1493 ( .a ({new_AGEMA_signal_4084, new_AGEMA_signal_4083, rd_I_n2309}), .b ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, rd_I_n2311}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1490 ( .a ({new_AGEMA_signal_4110, new_AGEMA_signal_4109, rd_I_n2420}), .b ({new_AGEMA_signal_4610, new_AGEMA_signal_4609, rd_I_n2307}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1487 ( .a ({new_AGEMA_signal_3922, new_AGEMA_signal_3921, rd_I_n2302}), .b ({new_AGEMA_signal_4612, new_AGEMA_signal_4611, rd_I_n2304}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1484 ( .a ({new_AGEMA_signal_4000, new_AGEMA_signal_3999, rd_I_n2297}), .b ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, rd_I_n2299}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1479 ( .a ({new_AGEMA_signal_4366, new_AGEMA_signal_4365, rd_I_n2291}), .b ({new_AGEMA_signal_4616, new_AGEMA_signal_4615, rd_I_n2293}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1472 ( .a ({new_AGEMA_signal_3910, new_AGEMA_signal_3909, rd_I_n2278}), .b ({new_AGEMA_signal_4622, new_AGEMA_signal_4621, rd_I_n2280}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1469 ( .a ({new_AGEMA_signal_3904, new_AGEMA_signal_3903, rd_I_n2273}), .b ({new_AGEMA_signal_4624, new_AGEMA_signal_4623, rd_I_n2275}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1462 ( .a ({new_AGEMA_signal_4372, new_AGEMA_signal_4371, rd_I_n2266}), .b ({new_AGEMA_signal_4630, new_AGEMA_signal_4629, rd_I_n2268}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1459 ( .a ({new_AGEMA_signal_4026, new_AGEMA_signal_4025, rd_I_n2368}), .b ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, rd_I_n2264}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1456 ( .a ({new_AGEMA_signal_4338, new_AGEMA_signal_4337, rd_I_n2259}), .b ({new_AGEMA_signal_4634, new_AGEMA_signal_4633, rd_I_n2261}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1453 ( .a ({new_AGEMA_signal_4438, new_AGEMA_signal_4437, rd_I_n2254}), .b ({new_AGEMA_signal_4636, new_AGEMA_signal_4635, rd_I_n2256}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1448 ( .a ({new_AGEMA_signal_3886, new_AGEMA_signal_3885, rd_I_n2245}), .b ({new_AGEMA_signal_4640, new_AGEMA_signal_4639, rd_I_n2247}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1446 ( .a ({state_in_s2[225], state_in_s1[225], state_in_s0[225]}), .b ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, rd_I_n2243}), .c ({new_AGEMA_signal_3690, new_AGEMA_signal_3689, rd_I_n2587}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1444 ( .a ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, rd_I_n2242}), .b ({1'b0, 1'b0, rc[1]}), .c ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, rd_I_n2588}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1443 ( .a ({state_in_s2[1], state_in_s1[1], state_in_s0[1]}), .b ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, rd_I_n2241}), .c ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, rd_I_n2242}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1442 ( .a ({state_in_s2[278], state_in_s1[278], state_in_s0[278]}), .b ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, rd_I_n2240}), .c ({new_AGEMA_signal_3694, new_AGEMA_signal_3693, rd_I_n2590}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1439 ( .a ({new_AGEMA_signal_4152, new_AGEMA_signal_4151, rd_I_n2235}), .b ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, rd_I_n2237}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1436 ( .a ({new_AGEMA_signal_4098, new_AGEMA_signal_4097, rd_I_n2230}), .b ({new_AGEMA_signal_4646, new_AGEMA_signal_4645, rd_I_n2232}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1433 ( .a ({new_AGEMA_signal_4266, new_AGEMA_signal_4265, rd_I_n2225}), .b ({new_AGEMA_signal_4648, new_AGEMA_signal_4647, rd_I_n2227}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1430 ( .a ({new_AGEMA_signal_4416, new_AGEMA_signal_4415, rd_I_n2220}), .b ({new_AGEMA_signal_4650, new_AGEMA_signal_4649, rd_I_n2222}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1427 ( .a ({new_AGEMA_signal_4302, new_AGEMA_signal_4301, rd_I_n2251}), .b ({new_AGEMA_signal_4652, new_AGEMA_signal_4651, rd_I_n2218}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1424 ( .a ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, rd_I_n2216}), .b ({state_in_s2[68], state_in_s1[68], state_in_s0[68]}), .c ({new_AGEMA_signal_3696, new_AGEMA_signal_3695, rd_I_n2464}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1423 ( .a ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, rd_I_n2215}), .b ({state_in_s2[164], state_in_s1[164], state_in_s0[164]}), .c ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, rd_I_n2462}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1422 ( .a ({new_AGEMA_signal_3658, new_AGEMA_signal_3657, rd_I_n2214}), .b ({state_in_s2[345], state_in_s1[345], state_in_s0[345]}), .c ({new_AGEMA_signal_3700, new_AGEMA_signal_3699, rd_I_n2461}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1419 ( .a ({state_in_s2[91], state_in_s1[91], state_in_s0[91]}), .b ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, rd_I_n2212}), .c ({new_AGEMA_signal_3702, new_AGEMA_signal_3701, rd_I_n2469}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1418 ( .a ({state_in_s2[187], state_in_s1[187], state_in_s0[187]}), .b ({new_AGEMA_signal_3456, new_AGEMA_signal_3455, rd_I_n2211}), .c ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, rd_I_n2467}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1417 ( .a ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, rd_I_n2210}), .b ({state_in_s2[336], state_in_s1[336], state_in_s0[336]}), .c ({new_AGEMA_signal_3706, new_AGEMA_signal_3705, rd_I_n2466}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1414 ( .a ({new_AGEMA_signal_3934, new_AGEMA_signal_3933, rd_I_n2205}), .b ({new_AGEMA_signal_4658, new_AGEMA_signal_4657, rd_I_n2207}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1409 ( .a ({new_AGEMA_signal_4032, new_AGEMA_signal_4031, rd_I_n2196}), .b ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, rd_I_n2198}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1406 ( .a ({new_AGEMA_signal_4164, new_AGEMA_signal_4163, rd_I_n2191}), .b ({new_AGEMA_signal_4664, new_AGEMA_signal_4663, rd_I_n2193}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1401 ( .a ({new_AGEMA_signal_4444, new_AGEMA_signal_4443, rd_I_n2324}), .b ({new_AGEMA_signal_4668, new_AGEMA_signal_4667, rd_I_n2188}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1398 ( .a ({new_AGEMA_signal_3724, new_AGEMA_signal_3723, rd_I_n2381}), .b ({new_AGEMA_signal_4670, new_AGEMA_signal_4669, rd_I_n2186}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1395 ( .a ({new_AGEMA_signal_3718, new_AGEMA_signal_3717, rd_I_n2527}), .b ({new_AGEMA_signal_4672, new_AGEMA_signal_4671, rd_I_n2184}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1388 ( .a ({new_AGEMA_signal_3826, new_AGEMA_signal_3825, rd_I_n2171}), .b ({new_AGEMA_signal_4678, new_AGEMA_signal_4677, rd_I_n2173}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1385 ( .a ({new_AGEMA_signal_3832, new_AGEMA_signal_3831, rd_I_n2202}), .b ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, rd_I_n2169}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1378 ( .a ({new_AGEMA_signal_3784, new_AGEMA_signal_3783, rd_I_n2372}), .b ({new_AGEMA_signal_4686, new_AGEMA_signal_4685, rd_I_n2162}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1375 ( .a ({new_AGEMA_signal_3940, new_AGEMA_signal_3939, rd_I_n2157}), .b ({new_AGEMA_signal_4688, new_AGEMA_signal_4687, rd_I_n2159}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1372 ( .a ({new_AGEMA_signal_4086, new_AGEMA_signal_4085, rd_I_n2152}), .b ({new_AGEMA_signal_4690, new_AGEMA_signal_4689, rd_I_n2154}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1364 ( .a ({state_in_s2[269], state_in_s1[269], state_in_s0[269]}), .b ({new_AGEMA_signal_3438, new_AGEMA_signal_3437, rd_I_n2144}), .c ({new_AGEMA_signal_3708, new_AGEMA_signal_3707, rd_I_n2384}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1362 ( .a ({state_in_s2[248], state_in_s1[248], state_in_s0[248]}), .b ({new_AGEMA_signal_3604, new_AGEMA_signal_3603, rd_I_n2143}), .c ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, rd_I_n2385}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1361 ( .a ({1'b0, 1'b0, rc[24]}), .b ({new_AGEMA_signal_3712, new_AGEMA_signal_3711, rd_I_n2142}), .c ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, rd_I_n2387}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1360 ( .a ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, rd_I_n2141}), .b ({state_in_s2[24], state_in_s1[24], state_in_s0[24]}), .c ({new_AGEMA_signal_3712, new_AGEMA_signal_3711, rd_I_n2142}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1357 ( .a ({new_AGEMA_signal_3742, new_AGEMA_signal_3741, rd_I_n2593}), .b ({new_AGEMA_signal_4700, new_AGEMA_signal_4699, rd_I_n2139}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1352 ( .a ({state_in_s2[33], state_in_s1[33], state_in_s0[33]}), .b ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, rd_I_n2133}), .c ({new_AGEMA_signal_3714, new_AGEMA_signal_3713, rd_I_n2526}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1351 ( .a ({state_in_s2[129], state_in_s1[129], state_in_s0[129]}), .b ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, rd_I_n2241}), .c ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, rd_I_n2529}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1350 ( .a ({state_in_s2[310], state_in_s1[310], state_in_s0[310]}), .b ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, rd_I_n2132}), .c ({new_AGEMA_signal_3718, new_AGEMA_signal_3717, rd_I_n2527}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1347 ( .a ({new_AGEMA_signal_3790, new_AGEMA_signal_3789, rd_I_n2149}), .b ({new_AGEMA_signal_4706, new_AGEMA_signal_4705, rd_I_n2130}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1344 ( .a ({new_AGEMA_signal_4002, new_AGEMA_signal_4001, rd_I_n2125}), .b ({new_AGEMA_signal_4708, new_AGEMA_signal_4707, rd_I_n2127}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1341 ( .a ({state_in_s2[56], state_in_s1[56], state_in_s0[56]}), .b ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, rd_I_n2123}), .c ({new_AGEMA_signal_3720, new_AGEMA_signal_3719, rd_I_n2380}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1340 ( .a ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, rd_I_n2141}), .b ({state_in_s2[152], state_in_s1[152], state_in_s0[152]}), .c ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, rd_I_n2383}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1339 ( .a ({state_in_s2[301], state_in_s1[301], state_in_s0[301]}), .b ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, rd_I_n2122}), .c ({new_AGEMA_signal_3724, new_AGEMA_signal_3723, rd_I_n2381}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1336 ( .a ({new_AGEMA_signal_3796, new_AGEMA_signal_3795, rd_I_n2117}), .b ({new_AGEMA_signal_4712, new_AGEMA_signal_4711, rd_I_n2119}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1333 ( .a ({new_AGEMA_signal_4398, new_AGEMA_signal_4397, rd_I_n2112}), .b ({new_AGEMA_signal_4714, new_AGEMA_signal_4713, rd_I_n2114}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1326 ( .a ({new_AGEMA_signal_3814, new_AGEMA_signal_3813, rd_I_n2358}), .b ({new_AGEMA_signal_4720, new_AGEMA_signal_4719, rd_I_n2105}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1321 ( .a ({state_in_s2[148], state_in_s1[148], state_in_s0[148]}), .b ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, rd_I_n2102}), .c ({new_AGEMA_signal_3726, new_AGEMA_signal_3725, rd_I_n2577}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1320 ( .a ({state_in_s2[297], state_in_s1[297], state_in_s0[297]}), .b ({new_AGEMA_signal_3538, new_AGEMA_signal_3537, rd_I_n2101}), .c ({new_AGEMA_signal_3728, new_AGEMA_signal_3727, rd_I_n2575}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1319 ( .a ({state_in_s2[52], state_in_s1[52], state_in_s0[52]}), .b ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, rd_I_n2100}), .c ({new_AGEMA_signal_3730, new_AGEMA_signal_3729, rd_I_n2574}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1316 ( .a ({state_in_s2[139], state_in_s1[139], state_in_s0[139]}), .b ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, rd_I_n2098}), .c ({new_AGEMA_signal_3732, new_AGEMA_signal_3731, rd_I_n2572}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1315 ( .a ({state_in_s2[288], state_in_s1[288], state_in_s0[288]}), .b ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, rd_I_n2097}), .c ({new_AGEMA_signal_3734, new_AGEMA_signal_3733, rd_I_n2570}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1314 ( .a ({state_in_s2[43], state_in_s1[43], state_in_s0[43]}), .b ({new_AGEMA_signal_3510, new_AGEMA_signal_3509, rd_I_n2096}), .c ({new_AGEMA_signal_3736, new_AGEMA_signal_3735, rd_I_n2569}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1309 ( .a ({new_AGEMA_signal_4176, new_AGEMA_signal_4175, rd_I_n2087}), .b ({new_AGEMA_signal_4730, new_AGEMA_signal_4729, rd_I_n2089}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1306 ( .a ({state_in_s2[54], state_in_s1[54], state_in_s0[54]}), .b ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, rd_I_n2132}), .c ({new_AGEMA_signal_3738, new_AGEMA_signal_3737, rd_I_n2592}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1305 ( .a ({state_in_s2[150], state_in_s1[150], state_in_s0[150]}), .b ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, rd_I_n2240}), .c ({new_AGEMA_signal_3740, new_AGEMA_signal_3739, rd_I_n2595}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1304 ( .a ({state_in_s2[299], state_in_s1[299], state_in_s0[299]}), .b ({new_AGEMA_signal_3510, new_AGEMA_signal_3509, rd_I_n2096}), .c ({new_AGEMA_signal_3742, new_AGEMA_signal_3741, rd_I_n2593}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1301 ( .a ({state_in_s2[63], state_in_s1[63], state_in_s0[63]}), .b ({new_AGEMA_signal_3436, new_AGEMA_signal_3435, rd_I_n2084}), .c ({new_AGEMA_signal_3744, new_AGEMA_signal_3743, rd_I_n2609}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1300 ( .a ({state_in_s2[159], state_in_s1[159], state_in_s0[159]}), .b ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, rd_I_n2083}), .c ({new_AGEMA_signal_3746, new_AGEMA_signal_3745, rd_I_n2612}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1299 ( .a ({state_in_s2[308], state_in_s1[308], state_in_s0[308]}), .b ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, rd_I_n2100}), .c ({new_AGEMA_signal_3748, new_AGEMA_signal_3747, rd_I_n2610}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1296 ( .a ({new_AGEMA_signal_3990, new_AGEMA_signal_3989, rd_I_n2364}), .b ({new_AGEMA_signal_4736, new_AGEMA_signal_4735, rd_I_n2081}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1293 ( .a ({state_in_s2[166], state_in_s1[166], state_in_s0[166]}), .b ({new_AGEMA_signal_3454, new_AGEMA_signal_3453, rd_I_n2079}), .c ({new_AGEMA_signal_3750, new_AGEMA_signal_3749, rd_I_n2445}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1292 ( .a ({state_in_s2[347], state_in_s1[347], state_in_s0[347]}), .b ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, rd_I_n2212}), .c ({new_AGEMA_signal_3752, new_AGEMA_signal_3751, rd_I_n2448}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1291 ( .a ({new_AGEMA_signal_3586, new_AGEMA_signal_3585, rd_I_n2078}), .b ({state_in_s2[70], state_in_s1[70], state_in_s0[70]}), .c ({new_AGEMA_signal_3754, new_AGEMA_signal_3753, rd_I_n2446}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1288 ( .a ({new_AGEMA_signal_4254, new_AGEMA_signal_4253, rd_I_n2073}), .b ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, rd_I_n2075}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1285 ( .a ({new_AGEMA_signal_4318, new_AGEMA_signal_4317, rd_I_n2068}), .b ({new_AGEMA_signal_4742, new_AGEMA_signal_4741, rd_I_n2070}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1274 ( .a ({new_AGEMA_signal_3772, new_AGEMA_signal_3771, rd_I_n2483}), .b ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, rd_I_n2053}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1269 ( .a ({new_AGEMA_signal_4150, new_AGEMA_signal_4149, rd_I_n2047}), .b ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, rd_I_n2049}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1264 ( .a ({state_in_s2[243], state_in_s1[243], state_in_s0[243]}), .b ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, rd_I_n2044}), .c ({new_AGEMA_signal_3756, new_AGEMA_signal_3755, rd_I_n2605}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1263 ( .a ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, rd_I_n2354}), .b ({state_in_s2[264], state_in_s1[264], state_in_s0[264]}), .c ({new_AGEMA_signal_3758, new_AGEMA_signal_3757, rd_I_n2608}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1262 ( .a ({new_AGEMA_signal_3550, new_AGEMA_signal_3549, rd_I_n2043}), .b ({new_AGEMA_signal_2122, new_AGEMA_signal_2121, rd_I_n2042}), .c ({new_AGEMA_signal_3760, new_AGEMA_signal_3759, rd_I_n2606}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1261 ( .a ({state_in_s2[19], state_in_s1[19], state_in_s0[19]}), .b ({1'b0, 1'b0, rc[19]}), .c ({new_AGEMA_signal_2122, new_AGEMA_signal_2121, rd_I_n2042}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1258 ( .a ({new_AGEMA_signal_3766, new_AGEMA_signal_3765, rd_I_n2429}), .b ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, rd_I_n2040}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1253 ( .a ({new_AGEMA_signal_4008, new_AGEMA_signal_4007, rd_I_n2181}), .b ({new_AGEMA_signal_4764, new_AGEMA_signal_4763, rd_I_n2037}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1250 ( .a ({new_AGEMA_signal_3846, new_AGEMA_signal_3845, rd_I_n2177}), .b ({new_AGEMA_signal_4766, new_AGEMA_signal_4765, rd_I_n2035}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1239 ( .a ({state_in_s2[147], state_in_s1[147], state_in_s0[147]}), .b ({new_AGEMA_signal_3550, new_AGEMA_signal_3549, rd_I_n2043}), .c ({new_AGEMA_signal_3762, new_AGEMA_signal_3761, rd_I_n2428}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1238 ( .a ({state_in_s2[296], state_in_s1[296], state_in_s0[296]}), .b ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, rd_I_n2355}), .c ({new_AGEMA_signal_3764, new_AGEMA_signal_3763, rd_I_n2431}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1237 ( .a ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, rd_I_n2029}), .b ({state_in_s2[51], state_in_s1[51], state_in_s0[51]}), .c ({new_AGEMA_signal_3766, new_AGEMA_signal_3765, rd_I_n2429}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1232 ( .a ({new_AGEMA_signal_4242, new_AGEMA_signal_4241, rd_I_n2424}), .b ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, rd_I_n2023}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1229 ( .a ({new_AGEMA_signal_3868, new_AGEMA_signal_3867, rd_I_n2018}), .b ({new_AGEMA_signal_4782, new_AGEMA_signal_4781, rd_I_n2020}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1226 ( .a ({state_in_s2[309], state_in_s1[309], state_in_s0[309]}), .b ({new_AGEMA_signal_3532, new_AGEMA_signal_3531, rd_I_n2016}), .c ({new_AGEMA_signal_3768, new_AGEMA_signal_3767, rd_I_n2482}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1225 ( .a ({state_in_s2[32], state_in_s1[32], state_in_s0[32]}), .b ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, rd_I_n2097}), .c ({new_AGEMA_signal_3770, new_AGEMA_signal_3769, rd_I_n2485}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1224 ( .a ({state_in_s2[128], state_in_s1[128], state_in_s0[128]}), .b ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, rd_I_n2015}), .c ({new_AGEMA_signal_3772, new_AGEMA_signal_3771, rd_I_n2483}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1221 ( .a ({new_AGEMA_signal_4056, new_AGEMA_signal_4055, rd_I_n2580}), .b ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, rd_I_n2013}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1218 ( .a ({state_in_s2[138], state_in_s1[138], state_in_s0[138]}), .b ({new_AGEMA_signal_3478, new_AGEMA_signal_3477, rd_I_n2011}), .c ({new_AGEMA_signal_3774, new_AGEMA_signal_3773, rd_I_n2533}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1217 ( .a ({state_in_s2[319], state_in_s1[319], state_in_s0[319]}), .b ({new_AGEMA_signal_3436, new_AGEMA_signal_3435, rd_I_n2084}), .c ({new_AGEMA_signal_3776, new_AGEMA_signal_3775, rd_I_n2531}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1216 ( .a ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, rd_I_n2010}), .b ({state_in_s2[42], state_in_s1[42], state_in_s0[42]}), .c ({new_AGEMA_signal_3778, new_AGEMA_signal_3777, rd_I_n2530}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1213 ( .a ({new_AGEMA_signal_4194, new_AGEMA_signal_4193, rd_I_n2005}), .b ({new_AGEMA_signal_4790, new_AGEMA_signal_4789, rd_I_n2007}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1210 ( .a ({new_AGEMA_signal_3862, new_AGEMA_signal_3861, rd_I_n2060}), .b ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, rd_I_n2003}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1207 ( .a ({new_AGEMA_signal_4378, new_AGEMA_signal_4377, rd_I_n1998}), .b ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, rd_I_n2000}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1200 ( .a ({new_AGEMA_signal_4396, new_AGEMA_signal_4395, rd_I_n1991}), .b ({new_AGEMA_signal_4800, new_AGEMA_signal_4799, rd_I_n1993}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1197 ( .a ({state_in_s2[306], state_in_s1[306], state_in_s0[306]}), .b ({new_AGEMA_signal_3634, new_AGEMA_signal_3633, rd_I_n1989}), .c ({new_AGEMA_signal_3780, new_AGEMA_signal_3779, rd_I_n2371}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1196 ( .a ({state_in_s2[61], state_in_s1[61], state_in_s0[61]}), .b ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, rd_I_n2353}), .c ({new_AGEMA_signal_3782, new_AGEMA_signal_3781, rd_I_n2374}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1195 ( .a ({state_in_s2[157], state_in_s1[157], state_in_s0[157]}), .b ({new_AGEMA_signal_3636, new_AGEMA_signal_3635, rd_I_n1988}), .c ({new_AGEMA_signal_3784, new_AGEMA_signal_3783, rd_I_n2372}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1192 ( .a ({new_AGEMA_signal_4288, new_AGEMA_signal_4287, rd_I_n2618}), .b ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, rd_I_n1986}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1189 ( .a ({new_AGEMA_signal_3952, new_AGEMA_signal_3951, rd_I_n1981}), .b ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, rd_I_n1983}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1186 ( .a ({new_AGEMA_signal_4356, new_AGEMA_signal_4355, rd_I_n1976}), .b ({new_AGEMA_signal_4808, new_AGEMA_signal_4807, rd_I_n1977}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1175 ( .a ({new_AGEMA_signal_3978, new_AGEMA_signal_3977, rd_I_n1967}), .b ({new_AGEMA_signal_4814, new_AGEMA_signal_4813, rd_I_n1969}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1170 ( .a ({state_in_s2[45], state_in_s1[45], state_in_s0[45]}), .b ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, rd_I_n2122}), .c ({new_AGEMA_signal_3786, new_AGEMA_signal_3785, rd_I_n2148}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1169 ( .a ({state_in_s2[141], state_in_s1[141], state_in_s0[141]}), .b ({new_AGEMA_signal_3438, new_AGEMA_signal_3437, rd_I_n2144}), .c ({new_AGEMA_signal_3788, new_AGEMA_signal_3787, rd_I_n2151}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1168 ( .a ({state_in_s2[290], state_in_s1[290], state_in_s0[290]}), .b ({new_AGEMA_signal_3444, new_AGEMA_signal_3443, rd_I_n1964}), .c ({new_AGEMA_signal_3790, new_AGEMA_signal_3789, rd_I_n2149}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1165 ( .a ({new_AGEMA_signal_4158, new_AGEMA_signal_4157, rd_I_n1959}), .b ({new_AGEMA_signal_4820, new_AGEMA_signal_4819, rd_I_n1961}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1162 ( .a ({new_AGEMA_signal_3894, new_AGEMA_signal_3893, rd_I_n2474}), .b ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, rd_I_n1957}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1157 ( .a ({new_AGEMA_signal_3802, new_AGEMA_signal_3801, rd_I_n2538}), .b ({new_AGEMA_signal_4826, new_AGEMA_signal_4825, rd_I_n1954}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1152 ( .a ({state_in_s2[66], state_in_s1[66], state_in_s0[66]}), .b ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, rd_I_n1951}), .c ({new_AGEMA_signal_3792, new_AGEMA_signal_3791, rd_I_n2120}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1151 ( .a ({state_in_s2[162], state_in_s1[162], state_in_s0[162]}), .b ({new_AGEMA_signal_3444, new_AGEMA_signal_3443, rd_I_n1964}), .c ({new_AGEMA_signal_3794, new_AGEMA_signal_3793, rd_I_n2118}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1150 ( .a ({state_in_s2[343], state_in_s1[343], state_in_s0[343]}), .b ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, rd_I_n1950}), .c ({new_AGEMA_signal_3796, new_AGEMA_signal_3795, rd_I_n2117}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1147 ( .a ({state_in_s2[192], state_in_s1[192], state_in_s0[192]}), .b ({new_AGEMA_signal_3508, new_AGEMA_signal_3507, rd_I_n1948}), .c ({new_AGEMA_signal_3798, new_AGEMA_signal_3797, rd_I_n2537}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1146 ( .a ({state_in_s2[373], state_in_s1[373], state_in_s0[373]}), .b ({new_AGEMA_signal_3480, new_AGEMA_signal_3479, rd_I_n1947}), .c ({new_AGEMA_signal_3800, new_AGEMA_signal_3799, rd_I_n2540}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1145 ( .a ({state_in_s2[96], state_in_s1[96], state_in_s0[96]}), .b ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, rd_I_n1946}), .c ({new_AGEMA_signal_3802, new_AGEMA_signal_3801, rd_I_n2538}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1140 ( .a ({new_AGEMA_signal_4186, new_AGEMA_signal_4185, rd_I_n1940}), .b ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, rd_I_n1942}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1137 ( .a ({new_AGEMA_signal_3580, new_AGEMA_signal_3579, rd_I_n1938}), .b ({state_in_s2[252], state_in_s1[252], state_in_s0[252]}), .c ({new_AGEMA_signal_3804, new_AGEMA_signal_3803, rd_I_n2341}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1136 ( .a ({new_AGEMA_signal_3568, new_AGEMA_signal_3567, rd_I_n1937}), .b ({state_in_s2[273], state_in_s1[273], state_in_s0[273]}), .c ({new_AGEMA_signal_3806, new_AGEMA_signal_3805, rd_I_n2339}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1135 ( .a ({new_AGEMA_signal_3472, new_AGEMA_signal_3471, rd_I_n1936}), .b ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, rd_I_n1935}), .c ({new_AGEMA_signal_3808, new_AGEMA_signal_3807, rd_I_n2338}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1134 ( .a ({state_in_s2[28], state_in_s1[28], state_in_s0[28]}), .b ({1'b0, 1'b0, rc[28]}), .c ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, rd_I_n1935}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1127 ( .a ({new_AGEMA_signal_3568, new_AGEMA_signal_3567, rd_I_n1937}), .b ({state_in_s2[145], state_in_s1[145], state_in_s0[145]}), .c ({new_AGEMA_signal_3810, new_AGEMA_signal_3809, rd_I_n2357}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1126 ( .a ({state_in_s2[294], state_in_s1[294], state_in_s0[294]}), .b ({new_AGEMA_signal_3454, new_AGEMA_signal_3453, rd_I_n2079}), .c ({new_AGEMA_signal_3812, new_AGEMA_signal_3811, rd_I_n2360}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1125 ( .a ({state_in_s2[49], state_in_s1[49], state_in_s0[49]}), .b ({new_AGEMA_signal_3460, new_AGEMA_signal_3459, rd_I_n1931}), .c ({new_AGEMA_signal_3814, new_AGEMA_signal_3813, rd_I_n2358}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1122 ( .a ({new_AGEMA_signal_4038, new_AGEMA_signal_4037, rd_I_n2065}), .b ({new_AGEMA_signal_4844, new_AGEMA_signal_4843, rd_I_n1929}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1119 ( .a ({state_in_s2[60], state_in_s1[60], state_in_s0[60]}), .b ({new_AGEMA_signal_3474, new_AGEMA_signal_3473, rd_I_n1927}), .c ({new_AGEMA_signal_3816, new_AGEMA_signal_3815, rd_I_n2330}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1118 ( .a ({state_in_s2[156], state_in_s1[156], state_in_s0[156]}), .b ({new_AGEMA_signal_3472, new_AGEMA_signal_3471, rd_I_n1936}), .c ({new_AGEMA_signal_3818, new_AGEMA_signal_3817, rd_I_n2328}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1117 ( .a ({state_in_s2[305], state_in_s1[305], state_in_s0[305]}), .b ({new_AGEMA_signal_3460, new_AGEMA_signal_3459, rd_I_n1931}), .c ({new_AGEMA_signal_3820, new_AGEMA_signal_3819, rd_I_n2327}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1110 ( .a ({state_in_s2[289], state_in_s1[289], state_in_s0[289]}), .b ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, rd_I_n2133}), .c ({new_AGEMA_signal_3822, new_AGEMA_signal_3821, rd_I_n2174}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1109 ( .a ({state_in_s2[44], state_in_s1[44], state_in_s0[44]}), .b ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, rd_I_n1923}), .c ({new_AGEMA_signal_3824, new_AGEMA_signal_3823, rd_I_n2172}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1108 ( .a ({state_in_s2[140], state_in_s1[140], state_in_s0[140]}), .b ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, rd_I_n1922}), .c ({new_AGEMA_signal_3826, new_AGEMA_signal_3825, rd_I_n2171}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1105 ( .a ({state_in_s2[312], state_in_s1[312], state_in_s0[312]}), .b ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, rd_I_n2123}), .c ({new_AGEMA_signal_3828, new_AGEMA_signal_3827, rd_I_n2201}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1104 ( .a ({state_in_s2[35], state_in_s1[35], state_in_s0[35]}), .b ({new_AGEMA_signal_3502, new_AGEMA_signal_3501, rd_I_n1920}), .c ({new_AGEMA_signal_3830, new_AGEMA_signal_3829, rd_I_n2204}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1103 ( .a ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, rd_I_n1919}), .b ({state_in_s2[131], state_in_s1[131], state_in_s0[131]}), .c ({new_AGEMA_signal_3832, new_AGEMA_signal_3831, rd_I_n2202}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1101 ( .a ({state_in_s2[268], state_in_s1[268], state_in_s0[268]}), .b ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, rd_I_n1922}), .c ({new_AGEMA_signal_3834, new_AGEMA_signal_3833, rd_I_n2515}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1099 ( .a ({state_in_s2[247], state_in_s1[247], state_in_s0[247]}), .b ({new_AGEMA_signal_3642, new_AGEMA_signal_3641, rd_I_n1917}), .c ({new_AGEMA_signal_3836, new_AGEMA_signal_3835, rd_I_n2516}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1098 ( .a ({1'b0, 1'b0, rc[23]}), .b ({new_AGEMA_signal_3838, new_AGEMA_signal_3837, rd_I_n1916}), .c ({new_AGEMA_signal_4856, new_AGEMA_signal_4855, rd_I_n2518}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1097 ( .a ({state_in_s2[23], state_in_s1[23], state_in_s0[23]}), .b ({new_AGEMA_signal_3646, new_AGEMA_signal_3645, rd_I_n1915}), .c ({new_AGEMA_signal_3838, new_AGEMA_signal_3837, rd_I_n1916}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1095 ( .a ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, rd_I_n1919}), .b ({state_in_s2[259], state_in_s1[259], state_in_s0[259]}), .c ({new_AGEMA_signal_3840, new_AGEMA_signal_3839, rd_I_n2510}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1093 ( .a ({state_in_s2[238], state_in_s1[238], state_in_s0[238]}), .b ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, rd_I_n1913}), .c ({new_AGEMA_signal_3842, new_AGEMA_signal_3841, rd_I_n2511}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1092 ( .a ({1'b0, 1'b0, rc[14]}), .b ({new_AGEMA_signal_3844, new_AGEMA_signal_3843, rd_I_n1912}), .c ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, rd_I_n2513}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1091 ( .a ({new_AGEMA_signal_3660, new_AGEMA_signal_3659, rd_I_n1911}), .b ({state_in_s2[14], state_in_s1[14], state_in_s0[14]}), .c ({new_AGEMA_signal_3844, new_AGEMA_signal_3843, rd_I_n1912}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1088 ( .a ({new_AGEMA_signal_3924, new_AGEMA_signal_3923, rd_I_n2433}), .b ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, rd_I_n1909}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1085 ( .a ({new_AGEMA_signal_4188, new_AGEMA_signal_4187, rd_I_n2136}), .b ({new_AGEMA_signal_4862, new_AGEMA_signal_4861, rd_I_n1907}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1077 ( .a ({state_in_s2[342], state_in_s1[342], state_in_s0[342]}), .b ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, rd_I_n1896}), .c ({new_AGEMA_signal_3846, new_AGEMA_signal_3845, rd_I_n2177}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1075 ( .a ({state_in_s2[161], state_in_s1[161], state_in_s0[161]}), .b ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, rd_I_n2133}), .c ({new_AGEMA_signal_3848, new_AGEMA_signal_3847, rd_I_n2179}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1074 ( .a ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, rd_I_n1895}), .b ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, rd_I_n1894}), .c ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, rd_I_n2133}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1073 ( .a ({state_in_s2[65], state_in_s1[65], state_in_s0[65]}), .b ({new_AGEMA_signal_3490, new_AGEMA_signal_3489, rd_I_n1893}), .c ({new_AGEMA_signal_3850, new_AGEMA_signal_3849, rd_I_n2176}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1070 ( .a ({state_in_s2[245], state_in_s1[245], state_in_s0[245]}), .b ({new_AGEMA_signal_3480, new_AGEMA_signal_3479, rd_I_n1947}), .c ({new_AGEMA_signal_3852, new_AGEMA_signal_3851, rd_I_n2549}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1069 ( .a ({state_in_s2[266], state_in_s1[266], state_in_s0[266]}), .b ({new_AGEMA_signal_3478, new_AGEMA_signal_3477, rd_I_n2011}), .c ({new_AGEMA_signal_3854, new_AGEMA_signal_3853, rd_I_n2547}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1068 ( .a ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, rd_I_n1891}), .b ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, rd_I_n1890}), .c ({new_AGEMA_signal_3856, new_AGEMA_signal_3855, rd_I_n2546}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1067 ( .a ({state_in_s2[21], state_in_s1[21], state_in_s0[21]}), .b ({1'b0, 1'b0, rc[21]}), .c ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, rd_I_n1890}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1064 ( .a ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, rd_I_n2010}), .b ({state_in_s2[298], state_in_s1[298], state_in_s0[298]}), .c ({new_AGEMA_signal_3858, new_AGEMA_signal_3857, rd_I_n2059}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1063 ( .a ({state_in_s2[53], state_in_s1[53], state_in_s0[53]}), .b ({new_AGEMA_signal_3532, new_AGEMA_signal_3531, rd_I_n2016}), .c ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, rd_I_n2062}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1062 ( .a ({state_in_s2[149], state_in_s1[149], state_in_s0[149]}), .b ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, rd_I_n1891}), .c ({new_AGEMA_signal_3862, new_AGEMA_signal_3861, rd_I_n2060}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1059 ( .a ({1'b0, 1'b0, rc[0]}), .b ({new_AGEMA_signal_3864, new_AGEMA_signal_3863, rd_I_n1887}), .c ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, rd_I_n2021}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1058 ( .a ({state_in_s2[0], state_in_s1[0], state_in_s0[0]}), .b ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, rd_I_n2015}), .c ({new_AGEMA_signal_3864, new_AGEMA_signal_3863, rd_I_n1887}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1057 ( .a ({state_in_s2[224], state_in_s1[224], state_in_s0[224]}), .b ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, rd_I_n1946}), .c ({new_AGEMA_signal_3866, new_AGEMA_signal_3865, rd_I_n2019}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1056 ( .a ({state_in_s2[277], state_in_s1[277], state_in_s0[277]}), .b ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, rd_I_n1891}), .c ({new_AGEMA_signal_3868, new_AGEMA_signal_3867, rd_I_n2018}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1055 ( .a ({new_AGEMA_signal_2932, new_AGEMA_signal_2931, rd_I_n1886}), .b ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, rd_I_n1885}), .c ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, rd_I_n1891}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1052 ( .a ({new_AGEMA_signal_4072, new_AGEMA_signal_4071, rd_I_n1900}), .b ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, rd_I_n1883}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1049 ( .a ({new_AGEMA_signal_4062, new_AGEMA_signal_4061, rd_I_n1904}), .b ({new_AGEMA_signal_4880, new_AGEMA_signal_4879, rd_I_n1881}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1046 ( .a ({state_in_s2[267], state_in_s1[267], state_in_s0[267]}), .b ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, rd_I_n2098}), .c ({new_AGEMA_signal_3870, new_AGEMA_signal_3869, rd_I_n2596}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1045 ( .a ({new_AGEMA_signal_3872, new_AGEMA_signal_3871, rd_I_n1879}), .b ({1'b0, 1'b0, rc[22]}), .c ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, rd_I_n2599}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1044 ( .a ({state_in_s2[22], state_in_s1[22], state_in_s0[22]}), .b ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, rd_I_n2240}), .c ({new_AGEMA_signal_3872, new_AGEMA_signal_3871, rd_I_n1879}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1043 ( .a ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, rd_I_n1878}), .b ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, rd_I_n1877}), .c ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, rd_I_n2240}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1042 ( .a ({state_in_s2[246], state_in_s1[246], state_in_s0[246]}), .b ({new_AGEMA_signal_3468, new_AGEMA_signal_3467, rd_I_n1876}), .c ({new_AGEMA_signal_3874, new_AGEMA_signal_3873, rd_I_n2597}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1040 ( .a ({state_in_s2[255], state_in_s1[255], state_in_s0[255]}), .b ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, rd_I_n1874}), .c ({new_AGEMA_signal_3876, new_AGEMA_signal_3875, rd_I_n2622}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1038 ( .a ({new_AGEMA_signal_3878, new_AGEMA_signal_3877, rd_I_n1873}), .b ({1'b0, 1'b0, rc[31]}), .c ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, rd_I_n2624}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1037 ( .a ({state_in_s2[31], state_in_s1[31], state_in_s0[31]}), .b ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, rd_I_n2083}), .c ({new_AGEMA_signal_3878, new_AGEMA_signal_3877, rd_I_n1873}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1036 ( .a ({state_in_s2[276], state_in_s1[276], state_in_s0[276]}), .b ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, rd_I_n2102}), .c ({new_AGEMA_signal_3880, new_AGEMA_signal_3879, rd_I_n2621}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1033 ( .a ({new_AGEMA_signal_4200, new_AGEMA_signal_4199, rd_I_n1868}), .b ({new_AGEMA_signal_4886, new_AGEMA_signal_4885, rd_I_n1870}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1030 ( .a ({state_in_s2[97], state_in_s1[97], state_in_s0[97]}), .b ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, rd_I_n2243}), .c ({new_AGEMA_signal_3882, new_AGEMA_signal_3881, rd_I_n2248}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1029 ( .a ({state_in_s2[193], state_in_s1[193], state_in_s0[193]}), .b ({new_AGEMA_signal_3490, new_AGEMA_signal_3489, rd_I_n1893}), .c ({new_AGEMA_signal_3884, new_AGEMA_signal_3883, rd_I_n2246}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1028 ( .a ({state_in_s2[374], state_in_s1[374], state_in_s0[374]}), .b ({new_AGEMA_signal_3468, new_AGEMA_signal_3467, rd_I_n1876}), .c ({new_AGEMA_signal_3886, new_AGEMA_signal_3885, rd_I_n2245}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1025 ( .a ({new_AGEMA_signal_4092, new_AGEMA_signal_4091, rd_I_n1862}), .b ({new_AGEMA_signal_4890, new_AGEMA_signal_4889, rd_I_n1864}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1020 ( .a ({new_AGEMA_signal_4320, new_AGEMA_signal_4319, rd_I_n1856}), .b ({new_AGEMA_signal_4894, new_AGEMA_signal_4893, rd_I_n1858}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1017 ( .a ({new_AGEMA_signal_3964, new_AGEMA_signal_3963, rd_I_n2416}), .b ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, rd_I_n1854}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U1014 ( .a ({new_AGEMA_signal_4206, new_AGEMA_signal_4205, rd_I_n2056}), .b ({new_AGEMA_signal_4898, new_AGEMA_signal_4897, rd_I_n1852}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1011 ( .a ({state_in_s2[371], state_in_s1[371], state_in_s0[371]}), .b ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, rd_I_n2044}), .c ({new_AGEMA_signal_3888, new_AGEMA_signal_3887, rd_I_n2561}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1010 ( .a ({state_in_s2[126], state_in_s1[126], state_in_s0[126]}), .b ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, rd_I_n1850}), .c ({new_AGEMA_signal_3890, new_AGEMA_signal_3889, rd_I_n2564}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1009 ( .a ({state_in_s2[222], state_in_s1[222], state_in_s0[222]}), .b ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, rd_I_n1849}), .c ({new_AGEMA_signal_3892, new_AGEMA_signal_3891, rd_I_n2562}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1003 ( .a ({state_in_s2[341], state_in_s1[341], state_in_s0[341]}), .b ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, rd_I_n1845}), .c ({new_AGEMA_signal_3894, new_AGEMA_signal_3893, rd_I_n2474}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1001 ( .a ({state_in_s2[160], state_in_s1[160], state_in_s0[160]}), .b ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, rd_I_n2097}), .c ({new_AGEMA_signal_3896, new_AGEMA_signal_3895, rd_I_n2476}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1000 ( .a ({new_AGEMA_signal_2970, new_AGEMA_signal_2969, rd_I_n1844}), .b ({new_AGEMA_signal_3034, new_AGEMA_signal_3033, rd_I_n1843}), .c ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, rd_I_n2097}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U999 ( .a ({state_in_s2[64], state_in_s1[64], state_in_s0[64]}), .b ({new_AGEMA_signal_3508, new_AGEMA_signal_3507, rd_I_n1948}), .c ({new_AGEMA_signal_3898, new_AGEMA_signal_3897, rd_I_n2473}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U988 ( .a ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, rd_I_n2215}), .b ({state_in_s2[36], state_in_s1[36], state_in_s0[36]}), .c ({new_AGEMA_signal_3900, new_AGEMA_signal_3899, rd_I_n2276}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U987 ( .a ({state_in_s2[132], state_in_s1[132], state_in_s0[132]}), .b ({new_AGEMA_signal_3618, new_AGEMA_signal_3617, rd_I_n1834}), .c ({new_AGEMA_signal_3902, new_AGEMA_signal_3901, rd_I_n2274}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U986 ( .a ({state_in_s2[313], state_in_s1[313], state_in_s0[313]}), .b ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, rd_I_n1833}), .c ({new_AGEMA_signal_3904, new_AGEMA_signal_3903, rd_I_n2273}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U983 ( .a ({state_in_s2[59], state_in_s1[59], state_in_s0[59]}), .b ({new_AGEMA_signal_3456, new_AGEMA_signal_3455, rd_I_n2211}), .c ({new_AGEMA_signal_3906, new_AGEMA_signal_3905, rd_I_n2281}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U982 ( .a ({new_AGEMA_signal_3592, new_AGEMA_signal_3591, rd_I_n1831}), .b ({state_in_s2[155], state_in_s1[155], state_in_s0[155]}), .c ({new_AGEMA_signal_3908, new_AGEMA_signal_3907, rd_I_n2279}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U981 ( .a ({state_in_s2[304], state_in_s1[304], state_in_s0[304]}), .b ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, rd_I_n1830}), .c ({new_AGEMA_signal_3910, new_AGEMA_signal_3909, rd_I_n2278}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U978 ( .a ({new_AGEMA_signal_4248, new_AGEMA_signal_4247, rd_I_n1825}), .b ({new_AGEMA_signal_4920, new_AGEMA_signal_4919, rd_I_n1826}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U975 ( .a ({state_in_s2[318], state_in_s1[318], state_in_s0[318]}), .b ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, rd_I_n1823}), .c ({new_AGEMA_signal_3912, new_AGEMA_signal_3911, rd_I_n2486}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U974 ( .a ({state_in_s2[41], state_in_s1[41], state_in_s0[41]}), .b ({new_AGEMA_signal_3538, new_AGEMA_signal_3537, rd_I_n2101}), .c ({new_AGEMA_signal_3914, new_AGEMA_signal_3913, rd_I_n2489}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U973 ( .a ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, rd_I_n1822}), .b ({state_in_s2[137], state_in_s1[137], state_in_s0[137]}), .c ({new_AGEMA_signal_3916, new_AGEMA_signal_3915, rd_I_n2487}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U970 ( .a ({new_AGEMA_signal_4054, new_AGEMA_signal_4053, rd_I_n2584}), .b ({new_AGEMA_signal_4924, new_AGEMA_signal_4923, rd_I_n1820}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U967 ( .a ({new_AGEMA_signal_4410, new_AGEMA_signal_4409, rd_I_n1815}), .b ({new_AGEMA_signal_4926, new_AGEMA_signal_4925, rd_I_n1817}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U962 ( .a ({state_in_s2[120], state_in_s1[120], state_in_s0[120]}), .b ({new_AGEMA_signal_3604, new_AGEMA_signal_3603, rd_I_n2143}), .c ({new_AGEMA_signal_3918, new_AGEMA_signal_3917, rd_I_n2305}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U961 ( .a ({state_in_s2[216], state_in_s1[216], state_in_s0[216]}), .b ({new_AGEMA_signal_3504, new_AGEMA_signal_3503, rd_I_n1812}), .c ({new_AGEMA_signal_3920, new_AGEMA_signal_3919, rd_I_n2303}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U960 ( .a ({new_AGEMA_signal_3654, new_AGEMA_signal_3653, rd_I_n1811}), .b ({state_in_s2[365], state_in_s1[365], state_in_s0[365]}), .c ({new_AGEMA_signal_3922, new_AGEMA_signal_3921, rd_I_n2302}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U957 ( .a ({new_AGEMA_signal_4230, new_AGEMA_signal_4229, rd_I_n2093}), .b ({new_AGEMA_signal_4930, new_AGEMA_signal_4929, rd_I_n1809}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U953 ( .a ({state_in_s2[340], state_in_s1[340], state_in_s0[340]}), .b ({new_AGEMA_signal_3544, new_AGEMA_signal_3543, rd_I_n1803}), .c ({new_AGEMA_signal_3924, new_AGEMA_signal_3923, rd_I_n2433}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U951 ( .a ({state_in_s2[191], state_in_s1[191], state_in_s0[191]}), .b ({new_AGEMA_signal_3436, new_AGEMA_signal_3435, rd_I_n2084}), .c ({new_AGEMA_signal_3926, new_AGEMA_signal_3925, rd_I_n2435}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U950 ( .a ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, rd_I_n1802}), .b ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, rd_I_n1801}), .c ({new_AGEMA_signal_3436, new_AGEMA_signal_3435, rd_I_n2084}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U949 ( .a ({state_in_s2[95], state_in_s1[95], state_in_s0[95]}), .b ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, rd_I_n1800}), .c ({new_AGEMA_signal_3928, new_AGEMA_signal_3927, rd_I_n2432}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U944 ( .a ({new_AGEMA_signal_3958, new_AGEMA_signal_3957, rd_I_n2450}), .b ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, rd_I_n1797}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U941 ( .a ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, rd_I_n1795}), .b ({state_in_s2[58], state_in_s1[58], state_in_s0[58]}), .c ({new_AGEMA_signal_3930, new_AGEMA_signal_3929, rd_I_n2208}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U940 ( .a ({state_in_s2[154], state_in_s1[154], state_in_s0[154]}), .b ({new_AGEMA_signal_3672, new_AGEMA_signal_3671, rd_I_n1794}), .c ({new_AGEMA_signal_3932, new_AGEMA_signal_3931, rd_I_n2206}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U939 ( .a ({state_in_s2[303], state_in_s1[303], state_in_s0[303]}), .b ({new_AGEMA_signal_3622, new_AGEMA_signal_3621, rd_I_n1793}), .c ({new_AGEMA_signal_3934, new_AGEMA_signal_3933, rd_I_n2205}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U932 ( .a ({state_in_s2[13], state_in_s1[13], state_in_s0[13]}), .b ({new_AGEMA_signal_3936, new_AGEMA_signal_3935, rd_I_n1789}), .c ({new_AGEMA_signal_4946, new_AGEMA_signal_4945, rd_I_n2160}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U931 ( .a ({1'b0, 1'b0, rc[13]}), .b ({new_AGEMA_signal_3438, new_AGEMA_signal_3437, rd_I_n2144}), .c ({new_AGEMA_signal_3936, new_AGEMA_signal_3935, rd_I_n1789}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U930 ( .a ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, rd_I_n1788}), .b ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, rd_I_n1878}), .c ({new_AGEMA_signal_3438, new_AGEMA_signal_3437, rd_I_n2144}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U929 ( .a ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, rd_I_n1787}), .b ({state_in_s2[104], state_in_s1[104], state_in_s0[104]}), .c ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, rd_I_n1878}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U928 ( .a ({state_in_s2[360], state_in_s1[360], state_in_s0[360]}), .b ({state_in_s2[232], state_in_s1[232], state_in_s0[232]}), .c ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, rd_I_n1787}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U927 ( .a ({new_AGEMA_signal_3654, new_AGEMA_signal_3653, rd_I_n1811}), .b ({state_in_s2[237], state_in_s1[237], state_in_s0[237]}), .c ({new_AGEMA_signal_3938, new_AGEMA_signal_3937, rd_I_n2158}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U926 ( .a ({new_AGEMA_signal_3648, new_AGEMA_signal_3647, rd_I_n1786}), .b ({state_in_s2[258], state_in_s1[258], state_in_s0[258]}), .c ({new_AGEMA_signal_3940, new_AGEMA_signal_3939, rd_I_n2157}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U923 ( .a ({new_AGEMA_signal_4308, new_AGEMA_signal_4307, rd_I_n2458}), .b ({new_AGEMA_signal_4948, new_AGEMA_signal_4947, rd_I_n1784}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U916 ( .a ({new_AGEMA_signal_4380, new_AGEMA_signal_4379, rd_I_n1777}), .b ({new_AGEMA_signal_4952, new_AGEMA_signal_4951, rd_I_n1779}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U908 ( .a ({state_in_s2[236], state_in_s1[236], state_in_s0[236]}), .b ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, rd_I_n1772}), .c ({new_AGEMA_signal_3942, new_AGEMA_signal_3941, rd_I_n2520}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U906 ( .a ({state_in_s2[12], state_in_s1[12], state_in_s0[12]}), .b ({new_AGEMA_signal_3944, new_AGEMA_signal_3943, rd_I_n1771}), .c ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, rd_I_n2521}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U905 ( .a ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, rd_I_n1922}), .b ({1'b0, 1'b0, rc[12]}), .c ({new_AGEMA_signal_3944, new_AGEMA_signal_3943, rd_I_n1771}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U904 ( .a ({new_AGEMA_signal_2932, new_AGEMA_signal_2931, rd_I_n1886}), .b ({new_AGEMA_signal_3190, new_AGEMA_signal_3189, rd_I_n1770}), .c ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, rd_I_n1922}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U903 ( .a ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, rd_I_n1769}), .b ({state_in_s2[359], state_in_s1[359], state_in_s0[359]}), .c ({new_AGEMA_signal_2932, new_AGEMA_signal_2931, rd_I_n1886}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U902 ( .a ({state_in_s2[103], state_in_s1[103], state_in_s0[103]}), .b ({state_in_s2[231], state_in_s1[231], state_in_s0[231]}), .c ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, rd_I_n1769}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U901 ( .a ({state_in_s2[257], state_in_s1[257], state_in_s0[257]}), .b ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, rd_I_n2241}), .c ({new_AGEMA_signal_3946, new_AGEMA_signal_3945, rd_I_n2523}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U900 ( .a ({new_AGEMA_signal_3186, new_AGEMA_signal_3185, rd_I_n1768}), .b ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, rd_I_n1767}), .c ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, rd_I_n2241}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U897 ( .a ({state_in_s2[119], state_in_s1[119], state_in_s0[119]}), .b ({new_AGEMA_signal_3642, new_AGEMA_signal_3641, rd_I_n1917}), .c ({new_AGEMA_signal_3948, new_AGEMA_signal_3947, rd_I_n1984}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U896 ( .a ({state_in_s2[215], state_in_s1[215], state_in_s0[215]}), .b ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, rd_I_n1950}), .c ({new_AGEMA_signal_3950, new_AGEMA_signal_3949, rd_I_n1982}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U895 ( .a ({state_in_s2[364], state_in_s1[364], state_in_s0[364]}), .b ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, rd_I_n1772}), .c ({new_AGEMA_signal_3952, new_AGEMA_signal_3951, rd_I_n1981}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U892 ( .a ({state_in_s2[175], state_in_s1[175], state_in_s0[175]}), .b ({new_AGEMA_signal_3622, new_AGEMA_signal_3621, rd_I_n1793}), .c ({new_AGEMA_signal_3954, new_AGEMA_signal_3953, rd_I_n2449}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U891 ( .a ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, rd_I_n2216}), .b ({state_in_s2[324], state_in_s1[324], state_in_s0[324]}), .c ({new_AGEMA_signal_3956, new_AGEMA_signal_3955, rd_I_n2452}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U890 ( .a ({state_in_s2[79], state_in_s1[79], state_in_s0[79]}), .b ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, rd_I_n1764}), .c ({new_AGEMA_signal_3958, new_AGEMA_signal_3957, rd_I_n2450}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U883 ( .a ({new_AGEMA_signal_4048, new_AGEMA_signal_4047, rd_I_n2320}), .b ({new_AGEMA_signal_4970, new_AGEMA_signal_4969, rd_I_n1760}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U880 ( .a ({new_AGEMA_signal_4024, new_AGEMA_signal_4023, rd_I_n2026}), .b ({new_AGEMA_signal_4972, new_AGEMA_signal_4971, rd_I_n1758}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U871 ( .a ({state_in_s2[94], state_in_s1[94], state_in_s0[94]}), .b ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, rd_I_n1849}), .c ({new_AGEMA_signal_3960, new_AGEMA_signal_3959, rd_I_n2415}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U870 ( .a ({state_in_s2[190], state_in_s1[190], state_in_s0[190]}), .b ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, rd_I_n1823}), .c ({new_AGEMA_signal_3962, new_AGEMA_signal_3961, rd_I_n2418}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U869 ( .a ({state_in_s2[339], state_in_s1[339], state_in_s0[339]}), .b ({new_AGEMA_signal_3574, new_AGEMA_signal_3573, rd_I_n1753}), .c ({new_AGEMA_signal_3964, new_AGEMA_signal_3963, rd_I_n2416}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U866 ( .a ({new_AGEMA_signal_3660, new_AGEMA_signal_3659, rd_I_n1911}), .b ({state_in_s2[142], state_in_s1[142], state_in_s0[142]}), .c ({new_AGEMA_signal_3966, new_AGEMA_signal_3965, rd_I_n2503}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U865 ( .a ({state_in_s2[291], state_in_s1[291], state_in_s0[291]}), .b ({new_AGEMA_signal_3502, new_AGEMA_signal_3501, rd_I_n1920}), .c ({new_AGEMA_signal_3968, new_AGEMA_signal_3967, rd_I_n2501}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U864 ( .a ({state_in_s2[46], state_in_s1[46], state_in_s0[46]}), .b ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, rd_I_n1751}), .c ({new_AGEMA_signal_3970, new_AGEMA_signal_3969, rd_I_n2500}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U859 ( .a ({new_AGEMA_signal_4078, new_AGEMA_signal_4077, rd_I_n1840}), .b ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, rd_I_n1745}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U856 ( .a ({state_in_s2[151], state_in_s1[151], state_in_s0[151]}), .b ({new_AGEMA_signal_3646, new_AGEMA_signal_3645, rd_I_n1915}), .c ({new_AGEMA_signal_3972, new_AGEMA_signal_3971, rd_I_n2508}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U855 ( .a ({state_in_s2[300], state_in_s1[300], state_in_s0[300]}), .b ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, rd_I_n1923}), .c ({new_AGEMA_signal_3974, new_AGEMA_signal_3973, rd_I_n2506}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U854 ( .a ({state_in_s2[55], state_in_s1[55], state_in_s0[55]}), .b ({new_AGEMA_signal_3498, new_AGEMA_signal_3497, rd_I_n1743}), .c ({new_AGEMA_signal_3976, new_AGEMA_signal_3975, rd_I_n2505}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U850 ( .a ({state_in_s2[311], state_in_s1[311], state_in_s0[311]}), .b ({new_AGEMA_signal_3498, new_AGEMA_signal_3497, rd_I_n1743}), .c ({new_AGEMA_signal_3978, new_AGEMA_signal_3977, rd_I_n1967}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U848 ( .a ({new_AGEMA_signal_3648, new_AGEMA_signal_3647, rd_I_n1786}), .b ({state_in_s2[130], state_in_s1[130], state_in_s0[130]}), .c ({new_AGEMA_signal_3980, new_AGEMA_signal_3979, rd_I_n1968}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U847 ( .a ({state_in_s2[34], state_in_s1[34], state_in_s0[34]}), .b ({new_AGEMA_signal_3444, new_AGEMA_signal_3443, rd_I_n1964}), .c ({new_AGEMA_signal_3982, new_AGEMA_signal_3981, rd_I_n1970}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U846 ( .a ({new_AGEMA_signal_2994, new_AGEMA_signal_2993, rd_I_n1740}), .b ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, rd_I_n1739}), .c ({new_AGEMA_signal_3444, new_AGEMA_signal_3443, rd_I_n1964}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U843 ( .a ({new_AGEMA_signal_4144, new_AGEMA_signal_4143, rd_I_n2165}), .b ({new_AGEMA_signal_4994, new_AGEMA_signal_4993, rd_I_n1737}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U840 ( .a ({state_in_s2[359], state_in_s1[359], state_in_s0[359]}), .b ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, rd_I_n1735}), .c ({new_AGEMA_signal_3984, new_AGEMA_signal_3983, rd_I_n2392}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U839 ( .a ({state_in_s2[114], state_in_s1[114], state_in_s0[114]}), .b ({new_AGEMA_signal_3630, new_AGEMA_signal_3629, rd_I_n1734}), .c ({new_AGEMA_signal_3986, new_AGEMA_signal_3985, rd_I_n2390}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U838 ( .a ({state_in_s2[210], state_in_s1[210], state_in_s0[210]}), .b ({new_AGEMA_signal_3484, new_AGEMA_signal_3483, rd_I_n1733}), .c ({new_AGEMA_signal_3988, new_AGEMA_signal_3987, rd_I_n2389}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U836 ( .a ({state_in_s2[338], state_in_s1[338], state_in_s0[338]}), .b ({new_AGEMA_signal_3484, new_AGEMA_signal_3483, rd_I_n1733}), .c ({new_AGEMA_signal_3990, new_AGEMA_signal_3989, rd_I_n2364}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U834 ( .a ({state_in_s2[189], state_in_s1[189], state_in_s0[189]}), .b ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, rd_I_n2353}), .c ({new_AGEMA_signal_3992, new_AGEMA_signal_3991, rd_I_n2366}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U833 ( .a ({new_AGEMA_signal_3060, new_AGEMA_signal_3059, rd_I_n1731}), .b ({new_AGEMA_signal_2944, new_AGEMA_signal_2943, rd_I_n1730}), .c ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, rd_I_n2353}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U832 ( .a ({state_in_s2[93], state_in_s1[93], state_in_s0[93]}), .b ({new_AGEMA_signal_3562, new_AGEMA_signal_3561, rd_I_n1729}), .c ({new_AGEMA_signal_3994, new_AGEMA_signal_3993, rd_I_n2363}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U829 ( .a ({new_AGEMA_signal_4428, new_AGEMA_signal_4427, rd_I_n2454}), .b ({new_AGEMA_signal_5000, new_AGEMA_signal_4999, rd_I_n1727}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U824 ( .a ({state_in_s2[111], state_in_s1[111], state_in_s0[111]}), .b ({new_AGEMA_signal_3616, new_AGEMA_signal_3615, rd_I_n1724}), .c ({new_AGEMA_signal_3996, new_AGEMA_signal_3995, rd_I_n2300}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U823 ( .a ({state_in_s2[207], state_in_s1[207], state_in_s0[207]}), .b ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, rd_I_n1764}), .c ({new_AGEMA_signal_3998, new_AGEMA_signal_3997, rd_I_n2298}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U822 ( .a ({state_in_s2[356], state_in_s1[356], state_in_s0[356]}), .b ({new_AGEMA_signal_3666, new_AGEMA_signal_3665, rd_I_n1723}), .c ({new_AGEMA_signal_4000, new_AGEMA_signal_3999, rd_I_n2297}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U820 ( .a ({state_in_s2[77], state_in_s1[77], state_in_s0[77]}), .b ({new_AGEMA_signal_3652, new_AGEMA_signal_3651, rd_I_n1721}), .c ({new_AGEMA_signal_4002, new_AGEMA_signal_4001, rd_I_n2125}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U818 ( .a ({state_in_s2[322], state_in_s1[322], state_in_s0[322]}), .b ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, rd_I_n1951}), .c ({new_AGEMA_signal_4004, new_AGEMA_signal_4003, rd_I_n2126}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U817 ( .a ({state_in_s2[173], state_in_s1[173], state_in_s0[173]}), .b ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, rd_I_n2122}), .c ({new_AGEMA_signal_4006, new_AGEMA_signal_4005, rd_I_n2128}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U816 ( .a ({new_AGEMA_signal_2998, new_AGEMA_signal_2997, rd_I_n1720}), .b ({new_AGEMA_signal_3222, new_AGEMA_signal_3221, rd_I_n1719}), .c ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, rd_I_n2122}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U812 ( .a ({state_in_s2[333], state_in_s1[333], state_in_s0[333]}), .b ({new_AGEMA_signal_3652, new_AGEMA_signal_3651, rd_I_n1721}), .c ({new_AGEMA_signal_4008, new_AGEMA_signal_4007, rd_I_n2181}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U810 ( .a ({state_in_s2[184], state_in_s1[184], state_in_s0[184]}), .b ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, rd_I_n2123}), .c ({new_AGEMA_signal_4010, new_AGEMA_signal_4009, rd_I_n2183}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U809 ( .a ({new_AGEMA_signal_3234, new_AGEMA_signal_3233, rd_I_n1716}), .b ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, rd_I_n1895}), .c ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, rd_I_n2123}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U808 ( .a ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, rd_I_n1715}), .b ({state_in_s2[147], state_in_s1[147], state_in_s0[147]}), .c ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, rd_I_n1895}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U807 ( .a ({state_in_s2[275], state_in_s1[275], state_in_s0[275]}), .b ({state_in_s2[19], state_in_s1[19], state_in_s0[19]}), .c ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, rd_I_n1715}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U806 ( .a ({state_in_s2[88], state_in_s1[88], state_in_s0[88]}), .b ({new_AGEMA_signal_3504, new_AGEMA_signal_3503, rd_I_n1812}), .c ({new_AGEMA_signal_4012, new_AGEMA_signal_4011, rd_I_n2180}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U804 ( .a ({state_in_s2[72], state_in_s1[72], state_in_s0[72]}), .b ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, rd_I_n1713}), .c ({new_AGEMA_signal_4014, new_AGEMA_signal_4013, rd_I_n2436}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U802 ( .a ({state_in_s2[349], state_in_s1[349], state_in_s0[349]}), .b ({new_AGEMA_signal_3562, new_AGEMA_signal_3561, rd_I_n1729}), .c ({new_AGEMA_signal_4016, new_AGEMA_signal_4015, rd_I_n2437}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U801 ( .a ({state_in_s2[168], state_in_s1[168], state_in_s0[168]}), .b ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, rd_I_n2355}), .c ({new_AGEMA_signal_4018, new_AGEMA_signal_4017, rd_I_n2439}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U800 ( .a ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, rd_I_n1712}), .b ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, rd_I_n1801}), .c ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, rd_I_n2355}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U799 ( .a ({state_in_s2[154], state_in_s1[154], state_in_s0[154]}), .b ({new_AGEMA_signal_2152, new_AGEMA_signal_2151, rd_I_n1711}), .c ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, rd_I_n1801}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U798 ( .a ({state_in_s2[282], state_in_s1[282], state_in_s0[282]}), .b ({state_in_s2[26], state_in_s1[26], state_in_s0[26]}), .c ({new_AGEMA_signal_2152, new_AGEMA_signal_2151, rd_I_n1711}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U795 ( .a ({new_AGEMA_signal_4272, new_AGEMA_signal_4271, rd_I_n1706}), .b ({new_AGEMA_signal_5014, new_AGEMA_signal_5013, rd_I_n1708}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U792 ( .a ({state_in_s2[83], state_in_s1[83], state_in_s0[83]}), .b ({new_AGEMA_signal_3574, new_AGEMA_signal_3573, rd_I_n1753}), .c ({new_AGEMA_signal_4020, new_AGEMA_signal_4019, rd_I_n2025}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U791 ( .a ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, rd_I_n2029}), .b ({state_in_s2[179], state_in_s1[179], state_in_s0[179]}), .c ({new_AGEMA_signal_4022, new_AGEMA_signal_4021, rd_I_n2028}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U790 ( .a ({state_in_s2[328], state_in_s1[328], state_in_s0[328]}), .b ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, rd_I_n1713}), .c ({new_AGEMA_signal_4024, new_AGEMA_signal_4023, rd_I_n2026}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U786 ( .a ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, rd_I_n1702}), .b ({state_in_s2[134], state_in_s1[134], state_in_s0[134]}), .c ({new_AGEMA_signal_4026, new_AGEMA_signal_4025, rd_I_n2368}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U784 ( .a ({state_in_s2[38], state_in_s1[38], state_in_s0[38]}), .b ({new_AGEMA_signal_3454, new_AGEMA_signal_3453, rd_I_n2079}), .c ({new_AGEMA_signal_4028, new_AGEMA_signal_4027, rd_I_n2370}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U783 ( .a ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, rd_I_n1701}), .b ({new_AGEMA_signal_2944, new_AGEMA_signal_2943, rd_I_n1730}), .c ({new_AGEMA_signal_3454, new_AGEMA_signal_3453, rd_I_n2079}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U782 ( .a ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, rd_I_n1700}), .b ({state_in_s2[152], state_in_s1[152], state_in_s0[152]}), .c ({new_AGEMA_signal_2944, new_AGEMA_signal_2943, rd_I_n1730}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U781 ( .a ({state_in_s2[280], state_in_s1[280], state_in_s0[280]}), .b ({state_in_s2[24], state_in_s1[24], state_in_s0[24]}), .c ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, rd_I_n1700}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U780 ( .a ({state_in_s2[315], state_in_s1[315], state_in_s0[315]}), .b ({new_AGEMA_signal_3456, new_AGEMA_signal_3455, rd_I_n2211}), .c ({new_AGEMA_signal_4030, new_AGEMA_signal_4029, rd_I_n2367}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U779 ( .a ({new_AGEMA_signal_3274, new_AGEMA_signal_3273, rd_I_n1699}), .b ({new_AGEMA_signal_3226, new_AGEMA_signal_3225, rd_I_n1698}), .c ({new_AGEMA_signal_3456, new_AGEMA_signal_3455, rd_I_n2211}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U776 ( .a ({new_AGEMA_signal_4282, new_AGEMA_signal_4281, rd_I_n2108}), .b ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, rd_I_n1696}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U774 ( .a ({new_AGEMA_signal_3600, new_AGEMA_signal_3599, rd_I_n1694}), .b ({state_in_s2[90], state_in_s1[90], state_in_s0[90]}), .c ({new_AGEMA_signal_4032, new_AGEMA_signal_4031, rd_I_n2196}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U772 ( .a ({state_in_s2[335], state_in_s1[335], state_in_s0[335]}), .b ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, rd_I_n1764}), .c ({new_AGEMA_signal_4034, new_AGEMA_signal_4033, rd_I_n2197}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U771 ( .a ({new_AGEMA_signal_3154, new_AGEMA_signal_3153, rd_I_n1693}), .b ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, rd_I_n1692}), .c ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, rd_I_n1764}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U770 ( .a ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, rd_I_n1795}), .b ({state_in_s2[186], state_in_s1[186], state_in_s0[186]}), .c ({new_AGEMA_signal_4036, new_AGEMA_signal_4035, rd_I_n2199}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U768 ( .a ({state_in_s2[81], state_in_s1[81], state_in_s0[81]}), .b ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, rd_I_n1690}), .c ({new_AGEMA_signal_4038, new_AGEMA_signal_4037, rd_I_n2065}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U766 ( .a ({new_AGEMA_signal_3586, new_AGEMA_signal_3585, rd_I_n2078}), .b ({state_in_s2[326], state_in_s1[326], state_in_s0[326]}), .c ({new_AGEMA_signal_4040, new_AGEMA_signal_4039, rd_I_n2067}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U765 ( .a ({state_in_s2[177], state_in_s1[177], state_in_s0[177]}), .b ({new_AGEMA_signal_3460, new_AGEMA_signal_3459, rd_I_n1931}), .c ({new_AGEMA_signal_4042, new_AGEMA_signal_4041, rd_I_n2064}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U764 ( .a ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, rd_I_n1712}), .b ({new_AGEMA_signal_3390, new_AGEMA_signal_3389, rd_I_n1689}), .c ({new_AGEMA_signal_3460, new_AGEMA_signal_3459, rd_I_n1931}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U763 ( .a ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, rd_I_n1688}), .b ({state_in_s2[259], state_in_s1[259], state_in_s0[259]}), .c ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, rd_I_n1712}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U762 ( .a ({state_in_s2[3], state_in_s1[3], state_in_s0[3]}), .b ({state_in_s2[131], state_in_s1[131], state_in_s0[131]}), .c ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, rd_I_n1688}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U759 ( .a ({new_AGEMA_signal_4332, new_AGEMA_signal_4331, rd_I_n2284}), .b ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, rd_I_n1686}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U752 ( .a ({state_in_s2[92], state_in_s1[92], state_in_s0[92]}), .b ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, rd_I_n1679}), .c ({new_AGEMA_signal_4044, new_AGEMA_signal_4043, rd_I_n2319}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U751 ( .a ({state_in_s2[188], state_in_s1[188], state_in_s0[188]}), .b ({new_AGEMA_signal_3474, new_AGEMA_signal_3473, rd_I_n1927}), .c ({new_AGEMA_signal_4046, new_AGEMA_signal_4045, rd_I_n2322}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U750 ( .a ({state_in_s2[337], state_in_s1[337], state_in_s0[337]}), .b ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, rd_I_n1690}), .c ({new_AGEMA_signal_4048, new_AGEMA_signal_4047, rd_I_n2320}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U747 ( .a ({new_AGEMA_signal_4212, new_AGEMA_signal_4211, rd_I_n1806}), .b ({new_AGEMA_signal_5036, new_AGEMA_signal_5035, rd_I_n1677}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U742 ( .a ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, rd_I_n1822}), .b ({state_in_s2[265], state_in_s1[265], state_in_s0[265]}), .c ({new_AGEMA_signal_4050, new_AGEMA_signal_4049, rd_I_n2583}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U741 ( .a ({new_AGEMA_signal_4052, new_AGEMA_signal_4051, rd_I_n1674}), .b ({1'b0, 1'b0, rc[20]}), .c ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, rd_I_n2586}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U740 ( .a ({state_in_s2[20], state_in_s1[20], state_in_s0[20]}), .b ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, rd_I_n2102}), .c ({new_AGEMA_signal_4052, new_AGEMA_signal_4051, rd_I_n1674}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U739 ( .a ({new_AGEMA_signal_3286, new_AGEMA_signal_3285, rd_I_n1673}), .b ({new_AGEMA_signal_2952, new_AGEMA_signal_2951, rd_I_n1672}), .c ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, rd_I_n2102}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U738 ( .a ({state_in_s2[244], state_in_s1[244], state_in_s0[244]}), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, rd_I_n1671}), .c ({new_AGEMA_signal_4054, new_AGEMA_signal_4053, rd_I_n2584}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U736 ( .a ({state_in_s2[235], state_in_s1[235], state_in_s0[235]}), .b ({new_AGEMA_signal_3514, new_AGEMA_signal_3513, rd_I_n1669}), .c ({new_AGEMA_signal_4056, new_AGEMA_signal_4055, rd_I_n2580}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U734 ( .a ({state_in_s2[11], state_in_s1[11], state_in_s0[11]}), .b ({new_AGEMA_signal_4058, new_AGEMA_signal_4057, rd_I_n1668}), .c ({new_AGEMA_signal_5042, new_AGEMA_signal_5041, rd_I_n2582}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U733 ( .a ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, rd_I_n2098}), .b ({1'b0, 1'b0, rc[11]}), .c ({new_AGEMA_signal_4058, new_AGEMA_signal_4057, rd_I_n1668}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U732 ( .a ({new_AGEMA_signal_3318, new_AGEMA_signal_3317, rd_I_n1667}), .b ({new_AGEMA_signal_2952, new_AGEMA_signal_2951, rd_I_n1672}), .c ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, rd_I_n2098}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U731 ( .a ({state_in_s2[102], state_in_s1[102], state_in_s0[102]}), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, rd_I_n1666}), .c ({new_AGEMA_signal_2952, new_AGEMA_signal_2951, rd_I_n1672}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U730 ( .a ({state_in_s2[358], state_in_s1[358], state_in_s0[358]}), .b ({state_in_s2[230], state_in_s1[230], state_in_s0[230]}), .c ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, rd_I_n1666}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U729 ( .a ({state_in_s2[256], state_in_s1[256], state_in_s0[256]}), .b ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, rd_I_n2015}), .c ({new_AGEMA_signal_4060, new_AGEMA_signal_4059, rd_I_n2579}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U728 ( .a ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, rd_I_n1665}), .b ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, rd_I_n1664}), .c ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, rd_I_n2015}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U726 ( .a ({state_in_s2[363], state_in_s1[363], state_in_s0[363]}), .b ({new_AGEMA_signal_3514, new_AGEMA_signal_3513, rd_I_n1669}), .c ({new_AGEMA_signal_4062, new_AGEMA_signal_4061, rd_I_n1904}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U724 ( .a ({state_in_s2[214], state_in_s1[214], state_in_s0[214]}), .b ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, rd_I_n1896}), .c ({new_AGEMA_signal_4064, new_AGEMA_signal_4063, rd_I_n1906}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U723 ( .a ({state_in_s2[118], state_in_s1[118], state_in_s0[118]}), .b ({new_AGEMA_signal_3468, new_AGEMA_signal_3467, rd_I_n1876}), .c ({new_AGEMA_signal_4066, new_AGEMA_signal_4065, rd_I_n1903}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U722 ( .a ({new_AGEMA_signal_3016, new_AGEMA_signal_3015, rd_I_n1662}), .b ({new_AGEMA_signal_3330, new_AGEMA_signal_3329, rd_I_n1661}), .c ({new_AGEMA_signal_3468, new_AGEMA_signal_3467, rd_I_n1876}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U719 ( .a ({state_in_s2[127], state_in_s1[127], state_in_s0[127]}), .b ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, rd_I_n1874}), .c ({new_AGEMA_signal_4068, new_AGEMA_signal_4067, rd_I_n1899}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U718 ( .a ({state_in_s2[223], state_in_s1[223], state_in_s0[223]}), .b ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, rd_I_n1800}), .c ({new_AGEMA_signal_4070, new_AGEMA_signal_4069, rd_I_n1902}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U717 ( .a ({state_in_s2[372], state_in_s1[372], state_in_s0[372]}), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, rd_I_n1671}), .c ({new_AGEMA_signal_4072, new_AGEMA_signal_4071, rd_I_n1900}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U712 ( .a ({new_AGEMA_signal_4450, new_AGEMA_signal_4449, rd_I_n1654}), .b ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, rd_I_n1656}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U709 ( .a ({state_in_s2[302], state_in_s1[302], state_in_s0[302]}), .b ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, rd_I_n1751}), .c ({new_AGEMA_signal_4074, new_AGEMA_signal_4073, rd_I_n1839}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U708 ( .a ({state_in_s2[57], state_in_s1[57], state_in_s0[57]}), .b ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, rd_I_n1833}), .c ({new_AGEMA_signal_4076, new_AGEMA_signal_4075, rd_I_n1842}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U707 ( .a ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, rd_I_n1652}), .b ({state_in_s2[153], state_in_s1[153], state_in_s0[153]}), .c ({new_AGEMA_signal_4078, new_AGEMA_signal_4077, rd_I_n1840}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U704 ( .a ({state_in_s2[293], state_in_s1[293], state_in_s0[293]}), .b ({new_AGEMA_signal_3676, new_AGEMA_signal_3675, rd_I_n1650}), .c ({new_AGEMA_signal_4080, new_AGEMA_signal_4079, rd_I_n2312}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U703 ( .a ({state_in_s2[48], state_in_s1[48], state_in_s0[48]}), .b ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, rd_I_n1830}), .c ({new_AGEMA_signal_4082, new_AGEMA_signal_4081, rd_I_n2310}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U702 ( .a ({state_in_s2[144], state_in_s1[144], state_in_s0[144]}), .b ({new_AGEMA_signal_3678, new_AGEMA_signal_3677, rd_I_n1649}), .c ({new_AGEMA_signal_4084, new_AGEMA_signal_4083, rd_I_n2309}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U700 ( .a ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, rd_I_n1652}), .b ({state_in_s2[281], state_in_s1[281], state_in_s0[281]}), .c ({new_AGEMA_signal_4086, new_AGEMA_signal_4085, rd_I_n2152}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U698 ( .a ({state_in_s2[228], state_in_s1[228], state_in_s0[228]}), .b ({new_AGEMA_signal_3666, new_AGEMA_signal_3665, rd_I_n1723}), .c ({new_AGEMA_signal_4088, new_AGEMA_signal_4087, rd_I_n2153}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U697 ( .a ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, rd_I_n1647}), .b ({new_AGEMA_signal_3618, new_AGEMA_signal_3617, rd_I_n1834}), .c ({new_AGEMA_signal_4090, new_AGEMA_signal_4089, rd_I_n2155}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U696 ( .a ({state_in_s2[4], state_in_s1[4], state_in_s0[4]}), .b ({1'b0, 1'b0, rc[4]}), .c ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, rd_I_n1647}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U694 ( .a ({state_in_s2[272], state_in_s1[272], state_in_s0[272]}), .b ({new_AGEMA_signal_3678, new_AGEMA_signal_3677, rd_I_n1649}), .c ({new_AGEMA_signal_4092, new_AGEMA_signal_4091, rd_I_n1862}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U692 ( .a ({state_in_s2[251], state_in_s1[251], state_in_s0[251]}), .b ({new_AGEMA_signal_3588, new_AGEMA_signal_3587, rd_I_n1645}), .c ({new_AGEMA_signal_4094, new_AGEMA_signal_4093, rd_I_n1863}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U691 ( .a ({1'b0, 1'b0, rc[27]}), .b ({new_AGEMA_signal_4096, new_AGEMA_signal_4095, rd_I_n1644}), .c ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, rd_I_n1865}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U690 ( .a ({new_AGEMA_signal_3592, new_AGEMA_signal_3591, rd_I_n1831}), .b ({state_in_s2[27], state_in_s1[27], state_in_s0[27]}), .c ({new_AGEMA_signal_4096, new_AGEMA_signal_4095, rd_I_n1644}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U687 ( .a ({new_AGEMA_signal_4170, new_AGEMA_signal_4169, rd_I_n1748}), .b ({new_AGEMA_signal_5060, new_AGEMA_signal_5059, rd_I_n1642}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U683 ( .a ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, rd_I_n1639}), .b ({state_in_s2[334], state_in_s1[334], state_in_s0[334]}), .c ({new_AGEMA_signal_4098, new_AGEMA_signal_4097, rd_I_n2230}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U681 ( .a ({state_in_s2[185], state_in_s1[185], state_in_s0[185]}), .b ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, rd_I_n1833}), .c ({new_AGEMA_signal_4100, new_AGEMA_signal_4099, rd_I_n2231}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U680 ( .a ({new_AGEMA_signal_3106, new_AGEMA_signal_3105, rd_I_n1638}), .b ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, rd_I_n1739}), .c ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, rd_I_n1833}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U679 ( .a ({state_in_s2[148], state_in_s1[148], state_in_s0[148]}), .b ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, rd_I_n1637}), .c ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, rd_I_n1739}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U678 ( .a ({state_in_s2[276], state_in_s1[276], state_in_s0[276]}), .b ({state_in_s2[20], state_in_s1[20], state_in_s0[20]}), .c ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, rd_I_n1637}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U677 ( .a ({new_AGEMA_signal_3658, new_AGEMA_signal_3657, rd_I_n2214}), .b ({state_in_s2[89], state_in_s1[89], state_in_s0[89]}), .c ({new_AGEMA_signal_4102, new_AGEMA_signal_4101, rd_I_n2233}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U674 ( .a ({state_in_s2[231], state_in_s1[231], state_in_s0[231]}), .b ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, rd_I_n1735}), .c ({new_AGEMA_signal_4104, new_AGEMA_signal_4103, rd_I_n2397}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U673 ( .a ({state_in_s2[284], state_in_s1[284], state_in_s0[284]}), .b ({new_AGEMA_signal_3472, new_AGEMA_signal_3471, rd_I_n1936}), .c ({new_AGEMA_signal_4106, new_AGEMA_signal_4105, rd_I_n2395}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U672 ( .a ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, rd_I_n1635}), .b ({new_AGEMA_signal_3072, new_AGEMA_signal_3071, rd_I_n1634}), .c ({new_AGEMA_signal_3472, new_AGEMA_signal_3471, rd_I_n1936}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U671 ( .a ({new_AGEMA_signal_3628, new_AGEMA_signal_3627, rd_I_n1633}), .b ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, rd_I_n1632}), .c ({new_AGEMA_signal_4108, new_AGEMA_signal_4107, rd_I_n2394}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U670 ( .a ({state_in_s2[7], state_in_s1[7], state_in_s0[7]}), .b ({1'b0, 1'b0, rc[7]}), .c ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, rd_I_n1632}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U668 ( .a ({state_in_s2[135], state_in_s1[135], state_in_s0[135]}), .b ({new_AGEMA_signal_3628, new_AGEMA_signal_3627, rd_I_n1633}), .c ({new_AGEMA_signal_4110, new_AGEMA_signal_4109, rd_I_n2420}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U666 ( .a ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, rd_I_n1630}), .b ({state_in_s2[39], state_in_s1[39], state_in_s0[39]}), .c ({new_AGEMA_signal_4112, new_AGEMA_signal_4111, rd_I_n2422}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U665 ( .a ({state_in_s2[316], state_in_s1[316], state_in_s0[316]}), .b ({new_AGEMA_signal_3474, new_AGEMA_signal_3473, rd_I_n1927}), .c ({new_AGEMA_signal_4114, new_AGEMA_signal_4113, rd_I_n2419}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U664 ( .a ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, rd_I_n1629}), .b ({new_AGEMA_signal_3084, new_AGEMA_signal_3083, rd_I_n1628}), .c ({new_AGEMA_signal_3474, new_AGEMA_signal_3473, rd_I_n1927}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U657 ( .a ({state_in_s2[287], state_in_s1[287], state_in_s0[287]}), .b ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, rd_I_n2083}), .c ({new_AGEMA_signal_4116, new_AGEMA_signal_4115, rd_I_n2603}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U656 ( .a ({new_AGEMA_signal_3118, new_AGEMA_signal_3117, rd_I_n1624}), .b ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, rd_I_n1877}), .c ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, rd_I_n2083}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U655 ( .a ({state_in_s2[241], state_in_s1[241], state_in_s0[241]}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, rd_I_n1623}), .c ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, rd_I_n1877}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U654 ( .a ({state_in_s2[113], state_in_s1[113], state_in_s0[113]}), .b ({state_in_s2[369], state_in_s1[369], state_in_s0[369]}), .c ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, rd_I_n1623}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U653 ( .a ({state_in_s2[10], state_in_s1[10], state_in_s0[10]}), .b ({new_AGEMA_signal_4118, new_AGEMA_signal_4117, rd_I_n1622}), .c ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, rd_I_n2601}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U652 ( .a ({new_AGEMA_signal_3478, new_AGEMA_signal_3477, rd_I_n2011}), .b ({1'b0, 1'b0, rc[10]}), .c ({new_AGEMA_signal_4118, new_AGEMA_signal_4117, rd_I_n1622}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U651 ( .a ({new_AGEMA_signal_3076, new_AGEMA_signal_3075, rd_I_n1621}), .b ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, rd_I_n1767}), .c ({new_AGEMA_signal_3478, new_AGEMA_signal_3477, rd_I_n2011}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U650 ( .a ({state_in_s2[252], state_in_s1[252], state_in_s0[252]}), .b ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, rd_I_n1620}), .c ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, rd_I_n1767}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U649 ( .a ({state_in_s2[124], state_in_s1[124], state_in_s0[124]}), .b ({state_in_s2[380], state_in_s1[380], state_in_s0[380]}), .c ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, rd_I_n1620}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U648 ( .a ({state_in_s2[234], state_in_s1[234], state_in_s0[234]}), .b ({new_AGEMA_signal_3526, new_AGEMA_signal_3525, rd_I_n1619}), .c ({new_AGEMA_signal_4120, new_AGEMA_signal_4119, rd_I_n2600}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U646 ( .a ({state_in_s2[362], state_in_s1[362], state_in_s0[362]}), .b ({new_AGEMA_signal_3526, new_AGEMA_signal_3525, rd_I_n1619}), .c ({new_AGEMA_signal_4122, new_AGEMA_signal_4121, rd_I_n2556}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U644 ( .a ({state_in_s2[213], state_in_s1[213], state_in_s0[213]}), .b ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, rd_I_n1845}), .c ({new_AGEMA_signal_4124, new_AGEMA_signal_4123, rd_I_n2557}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U643 ( .a ({state_in_s2[117], state_in_s1[117], state_in_s0[117]}), .b ({new_AGEMA_signal_3480, new_AGEMA_signal_3479, rd_I_n1947}), .c ({new_AGEMA_signal_4126, new_AGEMA_signal_4125, rd_I_n2559}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U642 ( .a ({new_AGEMA_signal_3064, new_AGEMA_signal_3063, rd_I_n1617}), .b ({new_AGEMA_signal_2968, new_AGEMA_signal_2967, rd_I_n1616}), .c ({new_AGEMA_signal_3480, new_AGEMA_signal_3479, rd_I_n1947}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U639 ( .a ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, rd_I_n1630}), .b ({state_in_s2[167], state_in_s1[167], state_in_s0[167]}), .c ({new_AGEMA_signal_4128, new_AGEMA_signal_4127, rd_I_n2413}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U638 ( .a ({state_in_s2[348], state_in_s1[348], state_in_s0[348]}), .b ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, rd_I_n1679}), .c ({new_AGEMA_signal_4130, new_AGEMA_signal_4129, rd_I_n2411}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U637 ( .a ({state_in_s2[71], state_in_s1[71], state_in_s0[71]}), .b ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, rd_I_n1614}), .c ({new_AGEMA_signal_4132, new_AGEMA_signal_4131, rd_I_n2410}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U635 ( .a ({state_in_s2[199], state_in_s1[199], state_in_s0[199]}), .b ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, rd_I_n1614}), .c ({new_AGEMA_signal_4134, new_AGEMA_signal_4133, rd_I_n2400}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U633 ( .a ({state_in_s2[103], state_in_s1[103], state_in_s0[103]}), .b ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, rd_I_n1735}), .c ({new_AGEMA_signal_4136, new_AGEMA_signal_4135, rd_I_n2402}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U632 ( .a ({new_AGEMA_signal_3414, new_AGEMA_signal_3413, rd_I_n1612}), .b ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, rd_I_n1611}), .c ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, rd_I_n1735}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U631 ( .a ({new_AGEMA_signal_3580, new_AGEMA_signal_3579, rd_I_n1938}), .b ({state_in_s2[380], state_in_s1[380], state_in_s0[380]}), .c ({new_AGEMA_signal_4138, new_AGEMA_signal_4137, rd_I_n2399}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U628 ( .a ({state_in_s2[82], state_in_s1[82], state_in_s0[82]}), .b ({new_AGEMA_signal_3484, new_AGEMA_signal_3483, rd_I_n1733}), .c ({new_AGEMA_signal_4140, new_AGEMA_signal_4139, rd_I_n2164}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U627 ( .a ({new_AGEMA_signal_3146, new_AGEMA_signal_3145, rd_I_n1609}), .b ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, rd_I_n1608}), .c ({new_AGEMA_signal_3484, new_AGEMA_signal_3483, rd_I_n1733}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U626 ( .a ({state_in_s2[178], state_in_s1[178], state_in_s0[178]}), .b ({new_AGEMA_signal_3634, new_AGEMA_signal_3633, rd_I_n1989}), .c ({new_AGEMA_signal_4142, new_AGEMA_signal_4141, rd_I_n2167}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U625 ( .a ({state_in_s2[327], state_in_s1[327], state_in_s0[327]}), .b ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, rd_I_n1614}), .c ({new_AGEMA_signal_4144, new_AGEMA_signal_4143, rd_I_n2165}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U624 ( .a ({new_AGEMA_signal_3042, new_AGEMA_signal_3041, rd_I_n1607}), .b ({new_AGEMA_signal_3142, new_AGEMA_signal_3141, rd_I_n1606}), .c ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, rd_I_n1614}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U621 ( .a ({state_in_s2[172], state_in_s1[172], state_in_s0[172]}), .b ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, rd_I_n1923}), .c ({new_AGEMA_signal_4146, new_AGEMA_signal_4145, rd_I_n2050}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U620 ( .a ({new_AGEMA_signal_3022, new_AGEMA_signal_3021, rd_I_n1604}), .b ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, rd_I_n1603}), .c ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, rd_I_n1923}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U619 ( .a ({state_in_s2[321], state_in_s1[321], state_in_s0[321]}), .b ({new_AGEMA_signal_3490, new_AGEMA_signal_3489, rd_I_n1893}), .c ({new_AGEMA_signal_4148, new_AGEMA_signal_4147, rd_I_n2048}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U618 ( .a ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, rd_I_n1602}), .b ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, rd_I_n1601}), .c ({new_AGEMA_signal_3490, new_AGEMA_signal_3489, rd_I_n1893}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U617 ( .a ({state_in_s2[76], state_in_s1[76], state_in_s0[76]}), .b ({new_AGEMA_signal_3496, new_AGEMA_signal_3495, rd_I_n1600}), .c ({new_AGEMA_signal_4150, new_AGEMA_signal_4149, rd_I_n2047}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U615 ( .a ({state_in_s2[204], state_in_s1[204], state_in_s0[204]}), .b ({new_AGEMA_signal_3496, new_AGEMA_signal_3495, rd_I_n1600}), .c ({new_AGEMA_signal_4152, new_AGEMA_signal_4151, rd_I_n2235}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U613 ( .a ({state_in_s2[108], state_in_s1[108], state_in_s0[108]}), .b ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, rd_I_n1772}), .c ({new_AGEMA_signal_4154, new_AGEMA_signal_4153, rd_I_n2236}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U612 ( .a ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, rd_I_n1598}), .b ({new_AGEMA_signal_2968, new_AGEMA_signal_2967, rd_I_n1616}), .c ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, rd_I_n1772}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U611 ( .a ({state_in_s2[199], state_in_s1[199], state_in_s0[199]}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, rd_I_n1597}), .c ({new_AGEMA_signal_2968, new_AGEMA_signal_2967, rd_I_n1616}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U610 ( .a ({state_in_s2[327], state_in_s1[327], state_in_s0[327]}), .b ({state_in_s2[71], state_in_s1[71], state_in_s0[71]}), .c ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, rd_I_n1597}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U609 ( .a ({state_in_s2[353], state_in_s1[353], state_in_s0[353]}), .b ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, rd_I_n2243}), .c ({new_AGEMA_signal_4156, new_AGEMA_signal_4155, rd_I_n2238}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U608 ( .a ({new_AGEMA_signal_3174, new_AGEMA_signal_3173, rd_I_n1596}), .b ({new_AGEMA_signal_3012, new_AGEMA_signal_3011, rd_I_n1595}), .c ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, rd_I_n2243}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U606 ( .a ({state_in_s2[332], state_in_s1[332], state_in_s0[332]}), .b ({new_AGEMA_signal_3496, new_AGEMA_signal_3495, rd_I_n1600}), .c ({new_AGEMA_signal_4158, new_AGEMA_signal_4157, rd_I_n1959}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U605 ( .a ({new_AGEMA_signal_3178, new_AGEMA_signal_3177, rd_I_n1593}), .b ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, rd_I_n1592}), .c ({new_AGEMA_signal_3496, new_AGEMA_signal_3495, rd_I_n1600}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U603 ( .a ({state_in_s2[183], state_in_s1[183], state_in_s0[183]}), .b ({new_AGEMA_signal_3498, new_AGEMA_signal_3497, rd_I_n1743}), .c ({new_AGEMA_signal_4160, new_AGEMA_signal_4159, rd_I_n1960}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U602 ( .a ({new_AGEMA_signal_2986, new_AGEMA_signal_2985, rd_I_n1591}), .b ({new_AGEMA_signal_2970, new_AGEMA_signal_2969, rd_I_n1844}), .c ({new_AGEMA_signal_3498, new_AGEMA_signal_3497, rd_I_n1743}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U601 ( .a ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, rd_I_n1590}), .b ({state_in_s2[18], state_in_s1[18], state_in_s0[18]}), .c ({new_AGEMA_signal_2970, new_AGEMA_signal_2969, rd_I_n1844}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U600 ( .a ({state_in_s2[274], state_in_s1[274], state_in_s0[274]}), .b ({state_in_s2[146], state_in_s1[146], state_in_s0[146]}), .c ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, rd_I_n1590}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U599 ( .a ({state_in_s2[87], state_in_s1[87], state_in_s0[87]}), .b ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, rd_I_n1950}), .c ({new_AGEMA_signal_4162, new_AGEMA_signal_4161, rd_I_n1962}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U598 ( .a ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, rd_I_n1589}), .b ({new_AGEMA_signal_3198, new_AGEMA_signal_3197, rd_I_n1588}), .c ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, rd_I_n1950}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U596 ( .a ({new_AGEMA_signal_3606, new_AGEMA_signal_3605, rd_I_n1586}), .b ({state_in_s2[67], state_in_s1[67], state_in_s0[67]}), .c ({new_AGEMA_signal_4164, new_AGEMA_signal_4163, rd_I_n2191}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U594 ( .a ({state_in_s2[163], state_in_s1[163], state_in_s0[163]}), .b ({new_AGEMA_signal_3502, new_AGEMA_signal_3501, rd_I_n1920}), .c ({new_AGEMA_signal_4166, new_AGEMA_signal_4165, rd_I_n2194}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U593 ( .a ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, rd_I_n1585}), .b ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, rd_I_n1603}), .c ({new_AGEMA_signal_3502, new_AGEMA_signal_3501, rd_I_n1920}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U592 ( .a ({state_in_s2[30], state_in_s1[30], state_in_s0[30]}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, rd_I_n1584}), .c ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, rd_I_n1603}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U591 ( .a ({state_in_s2[286], state_in_s1[286], state_in_s0[286]}), .b ({state_in_s2[158], state_in_s1[158], state_in_s0[158]}), .c ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, rd_I_n1584}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U590 ( .a ({state_in_s2[344], state_in_s1[344], state_in_s0[344]}), .b ({new_AGEMA_signal_3504, new_AGEMA_signal_3503, rd_I_n1812}), .c ({new_AGEMA_signal_4168, new_AGEMA_signal_4167, rd_I_n2192}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U589 ( .a ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, rd_I_n1692}), .b ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, rd_I_n1601}), .c ({new_AGEMA_signal_3504, new_AGEMA_signal_3503, rd_I_n1812}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U588 ( .a ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, rd_I_n1583}), .b ({state_in_s2[179], state_in_s1[179], state_in_s0[179]}), .c ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, rd_I_n1601}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U587 ( .a ({state_in_s2[307], state_in_s1[307], state_in_s0[307]}), .b ({state_in_s2[51], state_in_s1[51], state_in_s0[51]}), .c ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, rd_I_n1583}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U586 ( .a ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, rd_I_n1582}), .b ({state_in_s2[298], state_in_s1[298], state_in_s0[298]}), .c ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, rd_I_n1692}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U585 ( .a ({state_in_s2[170], state_in_s1[170], state_in_s0[170]}), .b ({state_in_s2[42], state_in_s1[42], state_in_s0[42]}), .c ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, rd_I_n1582}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U582 ( .a ({new_AGEMA_signal_4344, new_AGEMA_signal_4343, rd_I_n2288}), .b ({new_AGEMA_signal_5092, new_AGEMA_signal_5091, rd_I_n1580}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U580 ( .a ({new_AGEMA_signal_3606, new_AGEMA_signal_3605, rd_I_n1586}), .b ({state_in_s2[323], state_in_s1[323], state_in_s0[323]}), .c ({new_AGEMA_signal_4170, new_AGEMA_signal_4169, rd_I_n1748}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U578 ( .a ({state_in_s2[174], state_in_s1[174], state_in_s0[174]}), .b ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, rd_I_n1751}), .c ({new_AGEMA_signal_4172, new_AGEMA_signal_4171, rd_I_n1750}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U577 ( .a ({new_AGEMA_signal_3402, new_AGEMA_signal_3401, rd_I_n1578}), .b ({new_AGEMA_signal_2986, new_AGEMA_signal_2985, rd_I_n1591}), .c ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, rd_I_n1751}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U576 ( .a ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, rd_I_n1577}), .b ({state_in_s2[137], state_in_s1[137], state_in_s0[137]}), .c ({new_AGEMA_signal_2986, new_AGEMA_signal_2985, rd_I_n1591}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U575 ( .a ({state_in_s2[9], state_in_s1[9], state_in_s0[9]}), .b ({state_in_s2[265], state_in_s1[265], state_in_s0[265]}), .c ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, rd_I_n1577}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U574 ( .a ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, rd_I_n1639}), .b ({state_in_s2[78], state_in_s1[78], state_in_s0[78]}), .c ({new_AGEMA_signal_4174, new_AGEMA_signal_4173, rd_I_n1747}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U572 ( .a ({state_in_s2[75], state_in_s1[75], state_in_s0[75]}), .b ({new_AGEMA_signal_3516, new_AGEMA_signal_3515, rd_I_n1575}), .c ({new_AGEMA_signal_4176, new_AGEMA_signal_4175, rd_I_n2087}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U570 ( .a ({state_in_s2[320], state_in_s1[320], state_in_s0[320]}), .b ({new_AGEMA_signal_3508, new_AGEMA_signal_3507, rd_I_n1948}), .c ({new_AGEMA_signal_4178, new_AGEMA_signal_4177, rd_I_n2088}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U569 ( .a ({new_AGEMA_signal_3046, new_AGEMA_signal_3045, rd_I_n1574}), .b ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, rd_I_n1589}), .c ({new_AGEMA_signal_3508, new_AGEMA_signal_3507, rd_I_n1948}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U568 ( .a ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, rd_I_n1573}), .b ({state_in_s2[306], state_in_s1[306], state_in_s0[306]}), .c ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, rd_I_n1589}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U567 ( .a ({state_in_s2[50], state_in_s1[50], state_in_s0[50]}), .b ({state_in_s2[178], state_in_s1[178], state_in_s0[178]}), .c ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, rd_I_n1573}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U566 ( .a ({state_in_s2[171], state_in_s1[171], state_in_s0[171]}), .b ({new_AGEMA_signal_3510, new_AGEMA_signal_3509, rd_I_n2096}), .c ({new_AGEMA_signal_4180, new_AGEMA_signal_4179, rd_I_n2090}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U565 ( .a ({new_AGEMA_signal_3058, new_AGEMA_signal_3057, rd_I_n1572}), .b ({new_AGEMA_signal_2994, new_AGEMA_signal_2993, rd_I_n1740}), .c ({new_AGEMA_signal_3510, new_AGEMA_signal_3509, rd_I_n2096}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U564 ( .a ({state_in_s2[157], state_in_s1[157], state_in_s0[157]}), .b ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, rd_I_n1571}), .c ({new_AGEMA_signal_2994, new_AGEMA_signal_2993, rd_I_n1740}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U563 ( .a ({state_in_s2[29], state_in_s1[29], state_in_s0[29]}), .b ({state_in_s2[285], state_in_s1[285], state_in_s0[285]}), .c ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, rd_I_n1571}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U560 ( .a ({state_in_s2[352], state_in_s1[352], state_in_s0[352]}), .b ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, rd_I_n1946}), .c ({new_AGEMA_signal_4182, new_AGEMA_signal_4181, rd_I_n1943}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U559 ( .a ({new_AGEMA_signal_3306, new_AGEMA_signal_3305, rd_I_n1569}), .b ({new_AGEMA_signal_3094, new_AGEMA_signal_3093, rd_I_n1568}), .c ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, rd_I_n1946}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U558 ( .a ({state_in_s2[107], state_in_s1[107], state_in_s0[107]}), .b ({new_AGEMA_signal_3514, new_AGEMA_signal_3513, rd_I_n1669}), .c ({new_AGEMA_signal_4184, new_AGEMA_signal_4183, rd_I_n1941}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U557 ( .a ({new_AGEMA_signal_3322, new_AGEMA_signal_3321, rd_I_n1567}), .b ({new_AGEMA_signal_3030, new_AGEMA_signal_3029, rd_I_n1566}), .c ({new_AGEMA_signal_3514, new_AGEMA_signal_3513, rd_I_n1669}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U556 ( .a ({state_in_s2[203], state_in_s1[203], state_in_s0[203]}), .b ({new_AGEMA_signal_3516, new_AGEMA_signal_3515, rd_I_n1575}), .c ({new_AGEMA_signal_4186, new_AGEMA_signal_4185, rd_I_n1940}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U554 ( .a ({state_in_s2[331], state_in_s1[331], state_in_s0[331]}), .b ({new_AGEMA_signal_3516, new_AGEMA_signal_3515, rd_I_n1575}), .c ({new_AGEMA_signal_4188, new_AGEMA_signal_4187, rd_I_n2136}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U553 ( .a ({new_AGEMA_signal_3310, new_AGEMA_signal_3309, rd_I_n1564}), .b ({new_AGEMA_signal_3054, new_AGEMA_signal_3053, rd_I_n1563}), .c ({new_AGEMA_signal_3516, new_AGEMA_signal_3515, rd_I_n1575}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U551 ( .a ({state_in_s2[182], state_in_s1[182], state_in_s0[182]}), .b ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, rd_I_n2132}), .c ({new_AGEMA_signal_4190, new_AGEMA_signal_4189, rd_I_n2138}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U550 ( .a ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, rd_I_n1802}), .b ({new_AGEMA_signal_2998, new_AGEMA_signal_2997, rd_I_n1720}), .c ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, rd_I_n2132}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U549 ( .a ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, rd_I_n1562}), .b ({state_in_s2[264], state_in_s1[264], state_in_s0[264]}), .c ({new_AGEMA_signal_2998, new_AGEMA_signal_2997, rd_I_n1720}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U548 ( .a ({state_in_s2[8], state_in_s1[8], state_in_s0[8]}), .b ({state_in_s2[136], state_in_s1[136], state_in_s0[136]}), .c ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, rd_I_n1562}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U547 ( .a ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, rd_I_n1561}), .b ({state_in_s2[273], state_in_s1[273], state_in_s0[273]}), .c ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, rd_I_n1802}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U546 ( .a ({state_in_s2[17], state_in_s1[17], state_in_s0[17]}), .b ({state_in_s2[145], state_in_s1[145], state_in_s0[145]}), .c ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, rd_I_n1561}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U545 ( .a ({state_in_s2[86], state_in_s1[86], state_in_s0[86]}), .b ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, rd_I_n1896}), .c ({new_AGEMA_signal_4192, new_AGEMA_signal_4191, rd_I_n2135}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U544 ( .a ({new_AGEMA_signal_3006, new_AGEMA_signal_3005, rd_I_n1560}), .b ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, rd_I_n1559}), .c ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, rd_I_n1896}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U542 ( .a ({state_in_s2[74], state_in_s1[74], state_in_s0[74]}), .b ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, rd_I_n1557}), .c ({new_AGEMA_signal_4194, new_AGEMA_signal_4193, rd_I_n2005}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U540 ( .a ({state_in_s2[351], state_in_s1[351], state_in_s0[351]}), .b ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, rd_I_n1800}), .c ({new_AGEMA_signal_4196, new_AGEMA_signal_4195, rd_I_n2006}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U539 ( .a ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, rd_I_n1556}), .b ({new_AGEMA_signal_3006, new_AGEMA_signal_3005, rd_I_n1560}), .c ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, rd_I_n1800}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U538 ( .a ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, rd_I_n1555}), .b ({state_in_s2[305], state_in_s1[305], state_in_s0[305]}), .c ({new_AGEMA_signal_3006, new_AGEMA_signal_3005, rd_I_n1560}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U537 ( .a ({state_in_s2[177], state_in_s1[177], state_in_s0[177]}), .b ({state_in_s2[49], state_in_s1[49], state_in_s0[49]}), .c ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, rd_I_n1555}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U536 ( .a ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, rd_I_n2010}), .b ({state_in_s2[170], state_in_s1[170], state_in_s0[170]}), .c ({new_AGEMA_signal_4198, new_AGEMA_signal_4197, rd_I_n2008}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U535 ( .a ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, rd_I_n1554}), .b ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, rd_I_n1894}), .c ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, rd_I_n2010}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U534 ( .a ({state_in_s2[28], state_in_s1[28], state_in_s0[28]}), .b ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, rd_I_n1553}), .c ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, rd_I_n1894}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U533 ( .a ({state_in_s2[156], state_in_s1[156], state_in_s0[156]}), .b ({state_in_s2[284], state_in_s1[284], state_in_s0[284]}), .c ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, rd_I_n1553}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U531 ( .a ({state_in_s2[202], state_in_s1[202], state_in_s0[202]}), .b ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, rd_I_n1557}), .c ({new_AGEMA_signal_4200, new_AGEMA_signal_4199, rd_I_n1868}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U529 ( .a ({state_in_s2[106], state_in_s1[106], state_in_s0[106]}), .b ({new_AGEMA_signal_3526, new_AGEMA_signal_3525, rd_I_n1619}), .c ({new_AGEMA_signal_4202, new_AGEMA_signal_4201, rd_I_n1869}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U528 ( .a ({new_AGEMA_signal_3130, new_AGEMA_signal_3129, rd_I_n1551}), .b ({new_AGEMA_signal_3012, new_AGEMA_signal_3011, rd_I_n1595}), .c ({new_AGEMA_signal_3526, new_AGEMA_signal_3525, rd_I_n1619}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U527 ( .a ({state_in_s2[348], state_in_s1[348], state_in_s0[348]}), .b ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, rd_I_n1550}), .c ({new_AGEMA_signal_3012, new_AGEMA_signal_3011, rd_I_n1595}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U526 ( .a ({state_in_s2[220], state_in_s1[220], state_in_s0[220]}), .b ({state_in_s2[92], state_in_s1[92], state_in_s0[92]}), .c ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, rd_I_n1550}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U525 ( .a ({state_in_s2[383], state_in_s1[383], state_in_s0[383]}), .b ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, rd_I_n1874}), .c ({new_AGEMA_signal_4204, new_AGEMA_signal_4203, rd_I_n1871}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U524 ( .a ({new_AGEMA_signal_3016, new_AGEMA_signal_3015, rd_I_n1662}), .b ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, rd_I_n1549}), .c ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, rd_I_n1874}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U523 ( .a ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, rd_I_n1548}), .b ({state_in_s2[81], state_in_s1[81], state_in_s0[81]}), .c ({new_AGEMA_signal_3016, new_AGEMA_signal_3015, rd_I_n1662}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U522 ( .a ({state_in_s2[209], state_in_s1[209], state_in_s0[209]}), .b ({state_in_s2[337], state_in_s1[337], state_in_s0[337]}), .c ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, rd_I_n1548}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U520 ( .a ({state_in_s2[330], state_in_s1[330], state_in_s0[330]}), .b ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, rd_I_n1557}), .c ({new_AGEMA_signal_4206, new_AGEMA_signal_4205, rd_I_n2056}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U519 ( .a ({new_AGEMA_signal_3126, new_AGEMA_signal_3125, rd_I_n1546}), .b ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, rd_I_n1602}), .c ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, rd_I_n1557}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U518 ( .a ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, rd_I_n1545}), .b ({state_in_s2[188], state_in_s1[188], state_in_s0[188]}), .c ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, rd_I_n1602}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U517 ( .a ({state_in_s2[316], state_in_s1[316], state_in_s0[316]}), .b ({state_in_s2[60], state_in_s1[60], state_in_s0[60]}), .c ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, rd_I_n1545}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U515 ( .a ({state_in_s2[181], state_in_s1[181], state_in_s0[181]}), .b ({new_AGEMA_signal_3532, new_AGEMA_signal_3531, rd_I_n2016}), .c ({new_AGEMA_signal_4208, new_AGEMA_signal_4207, rd_I_n2058}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U514 ( .a ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, rd_I_n1544}), .b ({new_AGEMA_signal_3022, new_AGEMA_signal_3021, rd_I_n1604}), .c ({new_AGEMA_signal_3532, new_AGEMA_signal_3531, rd_I_n2016}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U513 ( .a ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, rd_I_n1543}), .b ({state_in_s2[7], state_in_s1[7], state_in_s0[7]}), .c ({new_AGEMA_signal_3022, new_AGEMA_signal_3021, rd_I_n1604}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U512 ( .a ({state_in_s2[263], state_in_s1[263], state_in_s0[263]}), .b ({state_in_s2[135], state_in_s1[135], state_in_s0[135]}), .c ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, rd_I_n1543}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U511 ( .a ({state_in_s2[85], state_in_s1[85], state_in_s0[85]}), .b ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, rd_I_n1845}), .c ({new_AGEMA_signal_4210, new_AGEMA_signal_4209, rd_I_n2055}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U510 ( .a ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, rd_I_n1542}), .b ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, rd_I_n1592}), .c ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, rd_I_n1845}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U509 ( .a ({state_in_s2[167], state_in_s1[167], state_in_s0[167]}), .b ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, rd_I_n1541}), .c ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, rd_I_n1592}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U508 ( .a ({state_in_s2[295], state_in_s1[295], state_in_s0[295]}), .b ({state_in_s2[39], state_in_s1[39], state_in_s0[39]}), .c ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, rd_I_n1541}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U502 ( .a ({state_in_s2[361], state_in_s1[361], state_in_s0[361]}), .b ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, rd_I_n1537}), .c ({new_AGEMA_signal_4212, new_AGEMA_signal_4211, rd_I_n1806}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U500 ( .a ({state_in_s2[212], state_in_s1[212], state_in_s0[212]}), .b ({new_AGEMA_signal_3544, new_AGEMA_signal_3543, rd_I_n1803}), .c ({new_AGEMA_signal_4214, new_AGEMA_signal_4213, rd_I_n1808}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U499 ( .a ({state_in_s2[116], state_in_s1[116], state_in_s0[116]}), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, rd_I_n1671}), .c ({new_AGEMA_signal_4216, new_AGEMA_signal_4215, rd_I_n1805}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U498 ( .a ({new_AGEMA_signal_3294, new_AGEMA_signal_3293, rd_I_n1536}), .b ({new_AGEMA_signal_3030, new_AGEMA_signal_3029, rd_I_n1566}), .c ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, rd_I_n1671}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U497 ( .a ({state_in_s2[70], state_in_s1[70], state_in_s0[70]}), .b ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, rd_I_n1535}), .c ({new_AGEMA_signal_3030, new_AGEMA_signal_3029, rd_I_n1566}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U496 ( .a ({state_in_s2[198], state_in_s1[198], state_in_s0[198]}), .b ({state_in_s2[326], state_in_s1[326], state_in_s0[326]}), .c ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, rd_I_n1535}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U494 ( .a ({state_in_s2[73], state_in_s1[73], state_in_s0[73]}), .b ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, rd_I_n1533}), .c ({new_AGEMA_signal_4218, new_AGEMA_signal_4217, rd_I_n2477}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U492 ( .a ({state_in_s2[169], state_in_s1[169], state_in_s0[169]}), .b ({new_AGEMA_signal_3538, new_AGEMA_signal_3537, rd_I_n2101}), .c ({new_AGEMA_signal_4220, new_AGEMA_signal_4219, rd_I_n2480}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U491 ( .a ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, rd_I_n1532}), .b ({new_AGEMA_signal_3034, new_AGEMA_signal_3033, rd_I_n1843}), .c ({new_AGEMA_signal_3538, new_AGEMA_signal_3537, rd_I_n2101}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U490 ( .a ({state_in_s2[27], state_in_s1[27], state_in_s0[27]}), .b ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, rd_I_n1531}), .c ({new_AGEMA_signal_3034, new_AGEMA_signal_3033, rd_I_n1843}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U489 ( .a ({state_in_s2[283], state_in_s1[283], state_in_s0[283]}), .b ({state_in_s2[155], state_in_s1[155], state_in_s0[155]}), .c ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, rd_I_n1531}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U488 ( .a ({state_in_s2[350], state_in_s1[350], state_in_s0[350]}), .b ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, rd_I_n1849}), .c ({new_AGEMA_signal_4222, new_AGEMA_signal_4221, rd_I_n2478}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U487 ( .a ({new_AGEMA_signal_3042, new_AGEMA_signal_3041, rd_I_n1607}), .b ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, rd_I_n1542}), .c ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, rd_I_n1849}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U486 ( .a ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, rd_I_n1530}), .b ({state_in_s2[304], state_in_s1[304], state_in_s0[304]}), .c ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, rd_I_n1542}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U485 ( .a ({state_in_s2[176], state_in_s1[176], state_in_s0[176]}), .b ({state_in_s2[48], state_in_s1[48], state_in_s0[48]}), .c ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, rd_I_n1530}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U484 ( .a ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, rd_I_n1529}), .b ({state_in_s2[185], state_in_s1[185], state_in_s0[185]}), .c ({new_AGEMA_signal_3042, new_AGEMA_signal_3041, rd_I_n1607}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U483 ( .a ({state_in_s2[57], state_in_s1[57], state_in_s0[57]}), .b ({state_in_s2[313], state_in_s1[313], state_in_s0[313]}), .c ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, rd_I_n1529}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U480 ( .a ({state_in_s2[382], state_in_s1[382], state_in_s0[382]}), .b ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, rd_I_n1850}), .c ({new_AGEMA_signal_4224, new_AGEMA_signal_4223, rd_I_n2544}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U479 ( .a ({state_in_s2[105], state_in_s1[105], state_in_s0[105]}), .b ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, rd_I_n1537}), .c ({new_AGEMA_signal_4226, new_AGEMA_signal_4225, rd_I_n2542}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U478 ( .a ({state_in_s2[201], state_in_s1[201], state_in_s0[201]}), .b ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, rd_I_n1533}), .c ({new_AGEMA_signal_4228, new_AGEMA_signal_4227, rd_I_n2541}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U476 ( .a ({state_in_s2[329], state_in_s1[329], state_in_s0[329]}), .b ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, rd_I_n1533}), .c ({new_AGEMA_signal_4230, new_AGEMA_signal_4229, rd_I_n2093}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U475 ( .a ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, rd_I_n1608}), .b ({new_AGEMA_signal_3046, new_AGEMA_signal_3045, rd_I_n1574}), .c ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, rd_I_n1533}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U474 ( .a ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, rd_I_n1526}), .b ({state_in_s2[315], state_in_s1[315], state_in_s0[315]}), .c ({new_AGEMA_signal_3046, new_AGEMA_signal_3045, rd_I_n1574}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U473 ( .a ({state_in_s2[59], state_in_s1[59], state_in_s0[59]}), .b ({state_in_s2[187], state_in_s1[187], state_in_s0[187]}), .c ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, rd_I_n1526}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U472 ( .a ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, rd_I_n1525}), .b ({state_in_s2[36], state_in_s1[36], state_in_s0[36]}), .c ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, rd_I_n1608}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U471 ( .a ({state_in_s2[292], state_in_s1[292], state_in_s0[292]}), .b ({state_in_s2[164], state_in_s1[164], state_in_s0[164]}), .c ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, rd_I_n1525}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U469 ( .a ({state_in_s2[84], state_in_s1[84], state_in_s0[84]}), .b ({new_AGEMA_signal_3544, new_AGEMA_signal_3543, rd_I_n1803}), .c ({new_AGEMA_signal_4232, new_AGEMA_signal_4231, rd_I_n2092}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U468 ( .a ({new_AGEMA_signal_3102, new_AGEMA_signal_3101, rd_I_n1524}), .b ({new_AGEMA_signal_3054, new_AGEMA_signal_3053, rd_I_n1563}), .c ({new_AGEMA_signal_3544, new_AGEMA_signal_3543, rd_I_n1803}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U467 ( .a ({state_in_s2[38], state_in_s1[38], state_in_s0[38]}), .b ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, rd_I_n1523}), .c ({new_AGEMA_signal_3054, new_AGEMA_signal_3053, rd_I_n1563}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U466 ( .a ({state_in_s2[166], state_in_s1[166], state_in_s0[166]}), .b ({state_in_s2[294], state_in_s1[294], state_in_s0[294]}), .c ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, rd_I_n1523}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U465 ( .a ({state_in_s2[180], state_in_s1[180], state_in_s0[180]}), .b ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, rd_I_n2100}), .c ({new_AGEMA_signal_4234, new_AGEMA_signal_4233, rd_I_n2095}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U464 ( .a ({new_AGEMA_signal_3060, new_AGEMA_signal_3059, rd_I_n1731}), .b ({new_AGEMA_signal_3058, new_AGEMA_signal_3057, rd_I_n1572}), .c ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, rd_I_n2100}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U463 ( .a ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, rd_I_n1522}), .b ({state_in_s2[134], state_in_s1[134], state_in_s0[134]}), .c ({new_AGEMA_signal_3058, new_AGEMA_signal_3057, rd_I_n1572}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U462 ( .a ({state_in_s2[6], state_in_s1[6], state_in_s0[6]}), .b ({state_in_s2[262], state_in_s1[262], state_in_s0[262]}), .c ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, rd_I_n1522}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U461 ( .a ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, rd_I_n1521}), .b ({state_in_s2[15], state_in_s1[15], state_in_s0[15]}), .c ({new_AGEMA_signal_3060, new_AGEMA_signal_3059, rd_I_n1731}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U460 ( .a ({state_in_s2[271], state_in_s1[271], state_in_s0[271]}), .b ({state_in_s2[143], state_in_s1[143], state_in_s0[143]}), .c ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, rd_I_n1521}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U457 ( .a ({state_in_s2[254], state_in_s1[254], state_in_s0[254]}), .b ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, rd_I_n1850}), .c ({new_AGEMA_signal_4236, new_AGEMA_signal_4235, rd_I_n2554}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U456 ( .a ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, rd_I_n1611}), .b ({new_AGEMA_signal_3064, new_AGEMA_signal_3063, rd_I_n1617}), .c ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, rd_I_n1850}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U455 ( .a ({state_in_s2[336], state_in_s1[336], state_in_s0[336]}), .b ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, rd_I_n1519}), .c ({new_AGEMA_signal_3064, new_AGEMA_signal_3063, rd_I_n1617}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U454 ( .a ({state_in_s2[208], state_in_s1[208], state_in_s0[208]}), .b ({state_in_s2[80], state_in_s1[80], state_in_s0[80]}), .c ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, rd_I_n1519}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U453 ( .a ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, rd_I_n1518}), .b ({state_in_s2[89], state_in_s1[89], state_in_s0[89]}), .c ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, rd_I_n1611}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U452 ( .a ({state_in_s2[217], state_in_s1[217], state_in_s0[217]}), .b ({state_in_s2[345], state_in_s1[345], state_in_s0[345]}), .c ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, rd_I_n1518}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U451 ( .a ({state_in_s2[275], state_in_s1[275], state_in_s0[275]}), .b ({new_AGEMA_signal_3550, new_AGEMA_signal_3549, rd_I_n2043}), .c ({new_AGEMA_signal_4238, new_AGEMA_signal_4237, rd_I_n2552}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U450 ( .a ({new_AGEMA_signal_3076, new_AGEMA_signal_3075, rd_I_n1621}), .b ({new_AGEMA_signal_3072, new_AGEMA_signal_3071, rd_I_n1634}), .c ({new_AGEMA_signal_3550, new_AGEMA_signal_3549, rd_I_n2043}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U449 ( .a ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, rd_I_n1517}), .b ({state_in_s2[238], state_in_s1[238], state_in_s0[238]}), .c ({new_AGEMA_signal_3072, new_AGEMA_signal_3071, rd_I_n1634}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U448 ( .a ({state_in_s2[366], state_in_s1[366], state_in_s0[366]}), .b ({state_in_s2[110], state_in_s1[110], state_in_s0[110]}), .c ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, rd_I_n1517}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U447 ( .a ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, rd_I_n1516}), .b ({state_in_s2[357], state_in_s1[357], state_in_s0[357]}), .c ({new_AGEMA_signal_3076, new_AGEMA_signal_3075, rd_I_n1621}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U446 ( .a ({state_in_s2[229], state_in_s1[229], state_in_s0[229]}), .b ({state_in_s2[101], state_in_s1[101], state_in_s0[101]}), .c ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, rd_I_n1516}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U445 ( .a ({new_AGEMA_signal_4240, new_AGEMA_signal_4239, rd_I_n1515}), .b ({state_in_s2[30], state_in_s1[30], state_in_s0[30]}), .c ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, rd_I_n2551}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U444 ( .a ({new_AGEMA_signal_3556, new_AGEMA_signal_3555, rd_I_n1514}), .b ({1'b0, 1'b0, rc[30]}), .c ({new_AGEMA_signal_4240, new_AGEMA_signal_4239, rd_I_n1515}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U442 ( .a ({new_AGEMA_signal_3556, new_AGEMA_signal_3555, rd_I_n1514}), .b ({state_in_s2[158], state_in_s1[158], state_in_s0[158]}), .c ({new_AGEMA_signal_4242, new_AGEMA_signal_4241, rd_I_n2424}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U440 ( .a ({state_in_s2[62], state_in_s1[62], state_in_s0[62]}), .b ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, rd_I_n1823}), .c ({new_AGEMA_signal_4244, new_AGEMA_signal_4243, rd_I_n2426}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U439 ( .a ({new_AGEMA_signal_3270, new_AGEMA_signal_3269, rd_I_n1512}), .b ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, rd_I_n1544}), .c ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, rd_I_n1823}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U438 ( .a ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, rd_I_n1511}), .b ({state_in_s2[272], state_in_s1[272], state_in_s0[272]}), .c ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, rd_I_n1544}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U437 ( .a ({state_in_s2[16], state_in_s1[16], state_in_s0[16]}), .b ({state_in_s2[144], state_in_s1[144], state_in_s0[144]}), .c ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, rd_I_n1511}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U436 ( .a ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, rd_I_n2029}), .b ({state_in_s2[307], state_in_s1[307], state_in_s0[307]}), .c ({new_AGEMA_signal_4246, new_AGEMA_signal_4245, rd_I_n2423}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U435 ( .a ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, rd_I_n1554}), .b ({new_AGEMA_signal_3084, new_AGEMA_signal_3083, rd_I_n1628}), .c ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, rd_I_n2029}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U434 ( .a ({state_in_s2[142], state_in_s1[142], state_in_s0[142]}), .b ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, rd_I_n1510}), .c ({new_AGEMA_signal_3084, new_AGEMA_signal_3083, rd_I_n1628}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U433 ( .a ({state_in_s2[270], state_in_s1[270], state_in_s0[270]}), .b ({state_in_s2[14], state_in_s1[14], state_in_s0[14]}), .c ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, rd_I_n1510}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U432 ( .a ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, rd_I_n1509}), .b ({state_in_s2[5], state_in_s1[5], state_in_s0[5]}), .c ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, rd_I_n1554}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U431 ( .a ({state_in_s2[261], state_in_s1[261], state_in_s0[261]}), .b ({state_in_s2[133], state_in_s1[133], state_in_s0[133]}), .c ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, rd_I_n1509}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U429 ( .a ({new_AGEMA_signal_3556, new_AGEMA_signal_3555, rd_I_n1514}), .b ({state_in_s2[286], state_in_s1[286], state_in_s0[286]}), .c ({new_AGEMA_signal_4248, new_AGEMA_signal_4247, rd_I_n1825}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U428 ( .a ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, rd_I_n1507}), .b ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, rd_I_n1885}), .c ({new_AGEMA_signal_3556, new_AGEMA_signal_3555, rd_I_n1514}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U427 ( .a ({state_in_s2[112], state_in_s1[112], state_in_s0[112]}), .b ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, rd_I_n1506}), .c ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, rd_I_n1885}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U426 ( .a ({state_in_s2[240], state_in_s1[240], state_in_s0[240]}), .b ({state_in_s2[368], state_in_s1[368], state_in_s0[368]}), .c ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, rd_I_n1506}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U424 ( .a ({state_in_s2[233], state_in_s1[233], state_in_s0[233]}), .b ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, rd_I_n1537}), .c ({new_AGEMA_signal_4250, new_AGEMA_signal_4249, rd_I_n1827}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U423 ( .a ({new_AGEMA_signal_3262, new_AGEMA_signal_3261, rd_I_n1505}), .b ({new_AGEMA_signal_3094, new_AGEMA_signal_3093, rd_I_n1568}), .c ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, rd_I_n1537}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U422 ( .a ({state_in_s2[91], state_in_s1[91], state_in_s0[91]}), .b ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, rd_I_n1504}), .c ({new_AGEMA_signal_3094, new_AGEMA_signal_3093, rd_I_n1568}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U421 ( .a ({state_in_s2[219], state_in_s1[219], state_in_s0[219]}), .b ({state_in_s2[347], state_in_s1[347], state_in_s0[347]}), .c ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, rd_I_n1504}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U420 ( .a ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, rd_I_n1822}), .b ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, rd_I_n1503}), .c ({new_AGEMA_signal_4252, new_AGEMA_signal_4251, rd_I_n1828}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U419 ( .a ({state_in_s2[9], state_in_s1[9], state_in_s0[9]}), .b ({1'b0, 1'b0, rc[9]}), .c ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, rd_I_n1503}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U418 ( .a ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, rd_I_n1502}), .b ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, rd_I_n1664}), .c ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, rd_I_n1822}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U417 ( .a ({state_in_s2[251], state_in_s1[251], state_in_s0[251]}), .b ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, rd_I_n1501}), .c ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, rd_I_n1664}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U416 ( .a ({state_in_s2[379], state_in_s1[379], state_in_s0[379]}), .b ({state_in_s2[123], state_in_s1[123], state_in_s0[123]}), .c ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, rd_I_n1501}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U414 ( .a ({state_in_s2[125], state_in_s1[125], state_in_s0[125]}), .b ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, rd_I_n1499}), .c ({new_AGEMA_signal_4254, new_AGEMA_signal_4253, rd_I_n2073}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U412 ( .a ({state_in_s2[370], state_in_s1[370], state_in_s0[370]}), .b ({new_AGEMA_signal_3630, new_AGEMA_signal_3629, rd_I_n1734}), .c ({new_AGEMA_signal_4256, new_AGEMA_signal_4255, rd_I_n2074}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U411 ( .a ({state_in_s2[221], state_in_s1[221], state_in_s0[221]}), .b ({new_AGEMA_signal_3562, new_AGEMA_signal_3561, rd_I_n1729}), .c ({new_AGEMA_signal_4258, new_AGEMA_signal_4257, rd_I_n2076}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U410 ( .a ({new_AGEMA_signal_3102, new_AGEMA_signal_3101, rd_I_n1524}), .b ({new_AGEMA_signal_3150, new_AGEMA_signal_3149, rd_I_n1498}), .c ({new_AGEMA_signal_3562, new_AGEMA_signal_3561, rd_I_n1729}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U409 ( .a ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, rd_I_n1497}), .b ({state_in_s2[303], state_in_s1[303], state_in_s0[303]}), .c ({new_AGEMA_signal_3102, new_AGEMA_signal_3101, rd_I_n1524}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U408 ( .a ({state_in_s2[47], state_in_s1[47], state_in_s0[47]}), .b ({state_in_s2[175], state_in_s1[175], state_in_s0[175]}), .c ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, rd_I_n1497}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U401 ( .a ({state_in_s2[165], state_in_s1[165], state_in_s0[165]}), .b ({new_AGEMA_signal_3676, new_AGEMA_signal_3675, rd_I_n1650}), .c ({new_AGEMA_signal_4260, new_AGEMA_signal_4259, rd_I_n2317}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U400 ( .a ({new_AGEMA_signal_3600, new_AGEMA_signal_3599, rd_I_n1694}), .b ({state_in_s2[346], state_in_s1[346], state_in_s0[346]}), .c ({new_AGEMA_signal_4262, new_AGEMA_signal_4261, rd_I_n2315}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U399 ( .a ({state_in_s2[69], state_in_s1[69], state_in_s0[69]}), .b ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, rd_I_n1493}), .c ({new_AGEMA_signal_4264, new_AGEMA_signal_4263, rd_I_n2314}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U395 ( .a ({state_in_s2[325], state_in_s1[325], state_in_s0[325]}), .b ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, rd_I_n1493}), .c ({new_AGEMA_signal_4266, new_AGEMA_signal_4265, rd_I_n2225}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U393 ( .a ({state_in_s2[176], state_in_s1[176], state_in_s0[176]}), .b ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, rd_I_n1830}), .c ({new_AGEMA_signal_4268, new_AGEMA_signal_4267, rd_I_n2226}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U392 ( .a ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, rd_I_n1490}), .b ({new_AGEMA_signal_3106, new_AGEMA_signal_3105, rd_I_n1638}), .c ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, rd_I_n1830}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U391 ( .a ({state_in_s2[139], state_in_s1[139], state_in_s0[139]}), .b ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, rd_I_n1489}), .c ({new_AGEMA_signal_3106, new_AGEMA_signal_3105, rd_I_n1638}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U390 ( .a ({state_in_s2[267], state_in_s1[267], state_in_s0[267]}), .b ({state_in_s2[11], state_in_s1[11], state_in_s0[11]}), .c ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, rd_I_n1489}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U389 ( .a ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, rd_I_n2210}), .b ({state_in_s2[80], state_in_s1[80], state_in_s0[80]}), .c ({new_AGEMA_signal_4270, new_AGEMA_signal_4269, rd_I_n2228}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) rd_I_U386 ( .a ({new_AGEMA_signal_4326, new_AGEMA_signal_4325, rd_I_n1683}), .b ({new_AGEMA_signal_5140, new_AGEMA_signal_5139, rd_I_n1487}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U384 ( .a ({state_in_s2[104], state_in_s1[104], state_in_s0[104]}), .b ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, rd_I_n1485}), .c ({new_AGEMA_signal_4272, new_AGEMA_signal_4271, rd_I_n1706}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U382 ( .a ({state_in_s2[381], state_in_s1[381], state_in_s0[381]}), .b ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, rd_I_n1499}), .c ({new_AGEMA_signal_4274, new_AGEMA_signal_4273, rd_I_n1707}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U381 ( .a ({state_in_s2[200], state_in_s1[200], state_in_s0[200]}), .b ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, rd_I_n1713}), .c ({new_AGEMA_signal_4276, new_AGEMA_signal_4275, rd_I_n1709}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U380 ( .a ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, rd_I_n1556}), .b ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, rd_I_n1484}), .c ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, rd_I_n1713}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U379 ( .a ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, rd_I_n1483}), .b ({state_in_s2[58], state_in_s1[58], state_in_s0[58]}), .c ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, rd_I_n1556}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U378 ( .a ({state_in_s2[314], state_in_s1[314], state_in_s0[314]}), .b ({state_in_s2[186], state_in_s1[186], state_in_s0[186]}), .c ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, rd_I_n1483}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U375 ( .a ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, rd_I_n1702}), .b ({state_in_s2[262], state_in_s1[262], state_in_s0[262]}), .c ({new_AGEMA_signal_4278, new_AGEMA_signal_4277, rd_I_n2107}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U374 ( .a ({new_AGEMA_signal_4280, new_AGEMA_signal_4279, rd_I_n1481}), .b ({1'b0, 1'b0, rc[17]}), .c ({new_AGEMA_signal_5144, new_AGEMA_signal_5143, rd_I_n2110}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U373 ( .a ({state_in_s2[17], state_in_s1[17], state_in_s0[17]}), .b ({new_AGEMA_signal_3568, new_AGEMA_signal_3567, rd_I_n1937}), .c ({new_AGEMA_signal_4280, new_AGEMA_signal_4279, rd_I_n1481}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U372 ( .a ({new_AGEMA_signal_3382, new_AGEMA_signal_3381, rd_I_n1480}), .b ({new_AGEMA_signal_3114, new_AGEMA_signal_3113, rd_I_n1479}), .c ({new_AGEMA_signal_3568, new_AGEMA_signal_3567, rd_I_n1937}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U371 ( .a ({new_AGEMA_signal_3598, new_AGEMA_signal_3597, rd_I_n1478}), .b ({state_in_s2[241], state_in_s1[241], state_in_s0[241]}), .c ({new_AGEMA_signal_4282, new_AGEMA_signal_4281, rd_I_n2108}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U368 ( .a ({state_in_s2[285], state_in_s1[285], state_in_s0[285]}), .b ({new_AGEMA_signal_3636, new_AGEMA_signal_3635, rd_I_n1988}), .c ({new_AGEMA_signal_4284, new_AGEMA_signal_4283, rd_I_n2617}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U367 ( .a ({new_AGEMA_signal_4286, new_AGEMA_signal_4285, rd_I_n1476}), .b ({state_in_s2[8], state_in_s1[8], state_in_s0[8]}), .c ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, rd_I_n2620}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U366 ( .a ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, rd_I_n2354}), .b ({1'b0, 1'b0, rc[8]}), .c ({new_AGEMA_signal_4286, new_AGEMA_signal_4285, rd_I_n1476}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U365 ( .a ({new_AGEMA_signal_3118, new_AGEMA_signal_3117, rd_I_n1624}), .b ({new_AGEMA_signal_3114, new_AGEMA_signal_3113, rd_I_n1479}), .c ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, rd_I_n2354}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U364 ( .a ({state_in_s2[99], state_in_s1[99], state_in_s0[99]}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, rd_I_n1475}), .c ({new_AGEMA_signal_3114, new_AGEMA_signal_3113, rd_I_n1479}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U363 ( .a ({state_in_s2[355], state_in_s1[355], state_in_s0[355]}), .b ({state_in_s2[227], state_in_s1[227], state_in_s0[227]}), .c ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, rd_I_n1475}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U362 ( .a ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, rd_I_n1474}), .b ({state_in_s2[122], state_in_s1[122], state_in_s0[122]}), .c ({new_AGEMA_signal_3118, new_AGEMA_signal_3117, rd_I_n1624}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U361 ( .a ({state_in_s2[250], state_in_s1[250], state_in_s0[250]}), .b ({state_in_s2[378], state_in_s1[378], state_in_s0[378]}), .c ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, rd_I_n1474}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U360 ( .a ({state_in_s2[232], state_in_s1[232], state_in_s0[232]}), .b ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, rd_I_n1485}), .c ({new_AGEMA_signal_4288, new_AGEMA_signal_4287, rd_I_n2618}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U358 ( .a ({state_in_s2[360], state_in_s1[360], state_in_s0[360]}), .b ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, rd_I_n1485}), .c ({new_AGEMA_signal_4290, new_AGEMA_signal_4289, rd_I_n2343}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U357 ( .a ({new_AGEMA_signal_3162, new_AGEMA_signal_3161, rd_I_n1472}), .b ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, rd_I_n1549}), .c ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, rd_I_n1485}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U356 ( .a ({state_in_s2[346], state_in_s1[346], state_in_s0[346]}), .b ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, rd_I_n1471}), .c ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, rd_I_n1549}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U355 ( .a ({state_in_s2[218], state_in_s1[218], state_in_s0[218]}), .b ({state_in_s2[90], state_in_s1[90], state_in_s0[90]}), .c ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, rd_I_n1471}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U353 ( .a ({state_in_s2[211], state_in_s1[211], state_in_s0[211]}), .b ({new_AGEMA_signal_3574, new_AGEMA_signal_3573, rd_I_n1753}), .c ({new_AGEMA_signal_4292, new_AGEMA_signal_4291, rd_I_n2344}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U352 ( .a ({new_AGEMA_signal_3134, new_AGEMA_signal_3133, rd_I_n1470}), .b ({new_AGEMA_signal_3126, new_AGEMA_signal_3125, rd_I_n1546}), .c ({new_AGEMA_signal_3574, new_AGEMA_signal_3573, rd_I_n1753}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U351 ( .a ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, rd_I_n1469}), .b ({state_in_s2[165], state_in_s1[165], state_in_s0[165]}), .c ({new_AGEMA_signal_3126, new_AGEMA_signal_3125, rd_I_n1546}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U350 ( .a ({state_in_s2[37], state_in_s1[37], state_in_s0[37]}), .b ({state_in_s2[293], state_in_s1[293], state_in_s0[293]}), .c ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, rd_I_n1469}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U349 ( .a ({state_in_s2[115], state_in_s1[115], state_in_s0[115]}), .b ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, rd_I_n2044}), .c ({new_AGEMA_signal_4294, new_AGEMA_signal_4293, rd_I_n2346}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U348 ( .a ({new_AGEMA_signal_3138, new_AGEMA_signal_3137, rd_I_n1468}), .b ({new_AGEMA_signal_3130, new_AGEMA_signal_3129, rd_I_n1551}), .c ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, rd_I_n2044}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U347 ( .a ({state_in_s2[69], state_in_s1[69], state_in_s0[69]}), .b ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, rd_I_n1467}), .c ({new_AGEMA_signal_3130, new_AGEMA_signal_3129, rd_I_n1551}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U346 ( .a ({state_in_s2[197], state_in_s1[197], state_in_s0[197]}), .b ({state_in_s2[325], state_in_s1[325], state_in_s0[325]}), .c ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, rd_I_n1467}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U344 ( .a ({new_AGEMA_signal_3598, new_AGEMA_signal_3597, rd_I_n1478}), .b ({state_in_s2[369], state_in_s1[369], state_in_s0[369]}), .c ({new_AGEMA_signal_4296, new_AGEMA_signal_4295, rd_I_n2348}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U342 ( .a ({state_in_s2[220], state_in_s1[220], state_in_s0[220]}), .b ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, rd_I_n1679}), .c ({new_AGEMA_signal_4298, new_AGEMA_signal_4297, rd_I_n2349}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U341 ( .a ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, rd_I_n1465}), .b ({new_AGEMA_signal_3134, new_AGEMA_signal_3133, rd_I_n1470}), .c ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, rd_I_n1679}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U340 ( .a ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, rd_I_n1464}), .b ({state_in_s2[302], state_in_s1[302], state_in_s0[302]}), .c ({new_AGEMA_signal_3134, new_AGEMA_signal_3133, rd_I_n1470}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U339 ( .a ({state_in_s2[46], state_in_s1[46], state_in_s0[46]}), .b ({state_in_s2[174], state_in_s1[174], state_in_s0[174]}), .c ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, rd_I_n1464}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U338 ( .a ({state_in_s2[124], state_in_s1[124], state_in_s0[124]}), .b ({new_AGEMA_signal_3580, new_AGEMA_signal_3579, rd_I_n1938}), .c ({new_AGEMA_signal_4300, new_AGEMA_signal_4299, rd_I_n2351}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U337 ( .a ({new_AGEMA_signal_3138, new_AGEMA_signal_3137, rd_I_n1468}), .b ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, rd_I_n1463}), .c ({new_AGEMA_signal_3580, new_AGEMA_signal_3579, rd_I_n1938}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U336 ( .a ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, rd_I_n1462}), .b ({state_in_s2[334], state_in_s1[334], state_in_s0[334]}), .c ({new_AGEMA_signal_3138, new_AGEMA_signal_3137, rd_I_n1468}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U335 ( .a ({state_in_s2[206], state_in_s1[206], state_in_s0[206]}), .b ({state_in_s2[78], state_in_s1[78], state_in_s0[78]}), .c ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, rd_I_n1462}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U333 ( .a ({state_in_s2[112], state_in_s1[112], state_in_s0[112]}), .b ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, rd_I_n1460}), .c ({new_AGEMA_signal_4302, new_AGEMA_signal_4301, rd_I_n2251}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U331 ( .a ({new_AGEMA_signal_3670, new_AGEMA_signal_3669, rd_I_n1459}), .b ({state_in_s2[357], state_in_s1[357], state_in_s0[357]}), .c ({new_AGEMA_signal_4304, new_AGEMA_signal_4303, rd_I_n2253}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U330 ( .a ({state_in_s2[208], state_in_s1[208], state_in_s0[208]}), .b ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, rd_I_n2210}), .c ({new_AGEMA_signal_4306, new_AGEMA_signal_4305, rd_I_n2250}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U329 ( .a ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, rd_I_n1458}), .b ({new_AGEMA_signal_3142, new_AGEMA_signal_3141, rd_I_n1606}), .c ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, rd_I_n2210}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U328 ( .a ({state_in_s2[162], state_in_s1[162], state_in_s0[162]}), .b ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, rd_I_n1457}), .c ({new_AGEMA_signal_3142, new_AGEMA_signal_3141, rd_I_n1606}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U327 ( .a ({state_in_s2[34], state_in_s1[34], state_in_s0[34]}), .b ({state_in_s2[290], state_in_s1[290], state_in_s0[290]}), .c ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, rd_I_n1457}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U323 ( .a ({state_in_s2[368], state_in_s1[368], state_in_s0[368]}), .b ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, rd_I_n1460}), .c ({new_AGEMA_signal_4308, new_AGEMA_signal_4307, rd_I_n2458}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U321 ( .a ({state_in_s2[219], state_in_s1[219], state_in_s0[219]}), .b ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, rd_I_n2212}), .c ({new_AGEMA_signal_4310, new_AGEMA_signal_4309, rd_I_n2460}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U320 ( .a ({new_AGEMA_signal_3370, new_AGEMA_signal_3369, rd_I_n1454}), .b ({new_AGEMA_signal_3146, new_AGEMA_signal_3145, rd_I_n1609}), .c ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, rd_I_n2212}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U319 ( .a ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, rd_I_n1453}), .b ({state_in_s2[45], state_in_s1[45], state_in_s0[45]}), .c ({new_AGEMA_signal_3146, new_AGEMA_signal_3145, rd_I_n1609}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U318 ( .a ({state_in_s2[173], state_in_s1[173], state_in_s0[173]}), .b ({state_in_s2[301], state_in_s1[301], state_in_s0[301]}), .c ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, rd_I_n1453}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U317 ( .a ({state_in_s2[123], state_in_s1[123], state_in_s0[123]}), .b ({new_AGEMA_signal_3588, new_AGEMA_signal_3587, rd_I_n1645}), .c ({new_AGEMA_signal_4312, new_AGEMA_signal_4311, rd_I_n2457}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U314 ( .a ({state_in_s2[198], state_in_s1[198], state_in_s0[198]}), .b ({new_AGEMA_signal_3586, new_AGEMA_signal_3585, rd_I_n2078}), .c ({new_AGEMA_signal_4314, new_AGEMA_signal_4313, rd_I_n2071}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U313 ( .a ({new_AGEMA_signal_3154, new_AGEMA_signal_3153, rd_I_n1693}), .b ({new_AGEMA_signal_3150, new_AGEMA_signal_3149, rd_I_n1498}), .c ({new_AGEMA_signal_3586, new_AGEMA_signal_3585, rd_I_n2078}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U312 ( .a ({state_in_s2[312], state_in_s1[312], state_in_s0[312]}), .b ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, rd_I_n1451}), .c ({new_AGEMA_signal_3150, new_AGEMA_signal_3149, rd_I_n1498}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U311 ( .a ({state_in_s2[184], state_in_s1[184], state_in_s0[184]}), .b ({state_in_s2[56], state_in_s1[56], state_in_s0[56]}), .c ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, rd_I_n1451}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U310 ( .a ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, rd_I_n1450}), .b ({state_in_s2[161], state_in_s1[161], state_in_s0[161]}), .c ({new_AGEMA_signal_3154, new_AGEMA_signal_3153, rd_I_n1693}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U309 ( .a ({state_in_s2[33], state_in_s1[33], state_in_s0[33]}), .b ({state_in_s2[289], state_in_s1[289], state_in_s0[289]}), .c ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, rd_I_n1450}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U308 ( .a ({state_in_s2[379], state_in_s1[379], state_in_s0[379]}), .b ({new_AGEMA_signal_3588, new_AGEMA_signal_3587, rd_I_n1645}), .c ({new_AGEMA_signal_4316, new_AGEMA_signal_4315, rd_I_n2069}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U307 ( .a ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, rd_I_n1449}), .b ({new_AGEMA_signal_3258, new_AGEMA_signal_3257, rd_I_n1448}), .c ({new_AGEMA_signal_3588, new_AGEMA_signal_3587, rd_I_n1645}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U306 ( .a ({state_in_s2[102], state_in_s1[102], state_in_s0[102]}), .b ({new_AGEMA_signal_3594, new_AGEMA_signal_3593, rd_I_n1447}), .c ({new_AGEMA_signal_4318, new_AGEMA_signal_4317, rd_I_n2068}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U304 ( .a ({state_in_s2[230], state_in_s1[230], state_in_s0[230]}), .b ({new_AGEMA_signal_3594, new_AGEMA_signal_3593, rd_I_n1447}), .c ({new_AGEMA_signal_4320, new_AGEMA_signal_4319, rd_I_n1856}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U302 ( .a ({new_AGEMA_signal_4322, new_AGEMA_signal_4321, rd_I_n1445}), .b ({1'b0, 1'b0, rc[6]}), .c ({new_AGEMA_signal_5160, new_AGEMA_signal_5159, rd_I_n1857}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U301 ( .a ({state_in_s2[6], state_in_s1[6], state_in_s0[6]}), .b ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, rd_I_n1702}), .c ({new_AGEMA_signal_4322, new_AGEMA_signal_4321, rd_I_n1445}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U300 ( .a ({new_AGEMA_signal_3282, new_AGEMA_signal_3281, rd_I_n1444}), .b ({new_AGEMA_signal_3246, new_AGEMA_signal_3245, rd_I_n1443}), .c ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, rd_I_n1702}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U299 ( .a ({state_in_s2[283], state_in_s1[283], state_in_s0[283]}), .b ({new_AGEMA_signal_3592, new_AGEMA_signal_3591, rd_I_n1831}), .c ({new_AGEMA_signal_4324, new_AGEMA_signal_4323, rd_I_n1859}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U298 ( .a ({new_AGEMA_signal_3298, new_AGEMA_signal_3297, rd_I_n1442}), .b ({new_AGEMA_signal_3214, new_AGEMA_signal_3213, rd_I_n1441}), .c ({new_AGEMA_signal_3592, new_AGEMA_signal_3591, rd_I_n1831}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U296 ( .a ({state_in_s2[358], state_in_s1[358], state_in_s0[358]}), .b ({new_AGEMA_signal_3594, new_AGEMA_signal_3593, rd_I_n1447}), .c ({new_AGEMA_signal_4326, new_AGEMA_signal_4325, rd_I_n1683}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U295 ( .a ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, rd_I_n1439}), .b ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, rd_I_n1438}), .c ({new_AGEMA_signal_3594, new_AGEMA_signal_3593, rd_I_n1447}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U293 ( .a ({state_in_s2[209], state_in_s1[209], state_in_s0[209]}), .b ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, rd_I_n1690}), .c ({new_AGEMA_signal_4328, new_AGEMA_signal_4327, rd_I_n1685}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U292 ( .a ({new_AGEMA_signal_3166, new_AGEMA_signal_3165, rd_I_n1437}), .b ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, rd_I_n1484}), .c ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, rd_I_n1690}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U291 ( .a ({state_in_s2[35], state_in_s1[35], state_in_s0[35]}), .b ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, rd_I_n1436}), .c ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, rd_I_n1484}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U290 ( .a ({state_in_s2[291], state_in_s1[291], state_in_s0[291]}), .b ({state_in_s2[163], state_in_s1[163], state_in_s0[163]}), .c ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, rd_I_n1436}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U289 ( .a ({state_in_s2[113], state_in_s1[113], state_in_s0[113]}), .b ({new_AGEMA_signal_3598, new_AGEMA_signal_3597, rd_I_n1478}), .c ({new_AGEMA_signal_4330, new_AGEMA_signal_4329, rd_I_n1682}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U288 ( .a ({new_AGEMA_signal_3238, new_AGEMA_signal_3237, rd_I_n1435}), .b ({new_AGEMA_signal_3162, new_AGEMA_signal_3161, rd_I_n1472}), .c ({new_AGEMA_signal_3598, new_AGEMA_signal_3597, rd_I_n1478}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U287 ( .a ({state_in_s2[67], state_in_s1[67], state_in_s0[67]}), .b ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, rd_I_n1434}), .c ({new_AGEMA_signal_3162, new_AGEMA_signal_3161, rd_I_n1472}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U286 ( .a ({state_in_s2[195], state_in_s1[195], state_in_s0[195]}), .b ({state_in_s2[323], state_in_s1[323], state_in_s0[323]}), .c ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, rd_I_n1434}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U284 ( .a ({state_in_s2[122], state_in_s1[122], state_in_s0[122]}), .b ({new_AGEMA_signal_3624, new_AGEMA_signal_3623, rd_I_n1432}), .c ({new_AGEMA_signal_4332, new_AGEMA_signal_4331, rd_I_n2284}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U282 ( .a ({state_in_s2[367], state_in_s1[367], state_in_s0[367]}), .b ({new_AGEMA_signal_3616, new_AGEMA_signal_3615, rd_I_n1724}), .c ({new_AGEMA_signal_4334, new_AGEMA_signal_4333, rd_I_n2286}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U281 ( .a ({state_in_s2[218], state_in_s1[218], state_in_s0[218]}), .b ({new_AGEMA_signal_3600, new_AGEMA_signal_3599, rd_I_n1694}), .c ({new_AGEMA_signal_4336, new_AGEMA_signal_4335, rd_I_n2283}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U280 ( .a ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, rd_I_n1431}), .b ({new_AGEMA_signal_3166, new_AGEMA_signal_3165, rd_I_n1437}), .c ({new_AGEMA_signal_3600, new_AGEMA_signal_3599, rd_I_n1694}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U279 ( .a ({state_in_s2[44], state_in_s1[44], state_in_s0[44]}), .b ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, rd_I_n1430}), .c ({new_AGEMA_signal_3166, new_AGEMA_signal_3165, rd_I_n1437}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U278 ( .a ({state_in_s2[300], state_in_s1[300], state_in_s0[300]}), .b ({state_in_s2[172], state_in_s1[172], state_in_s0[172]}), .c ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, rd_I_n1430}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U274 ( .a ({state_in_s2[378], state_in_s1[378], state_in_s0[378]}), .b ({new_AGEMA_signal_3624, new_AGEMA_signal_3623, rd_I_n1432}), .c ({new_AGEMA_signal_4338, new_AGEMA_signal_4337, rd_I_n2259}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U272 ( .a ({state_in_s2[197], state_in_s1[197], state_in_s0[197]}), .b ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, rd_I_n1493}), .c ({new_AGEMA_signal_4340, new_AGEMA_signal_4339, rd_I_n2260}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U271 ( .a ({new_AGEMA_signal_3202, new_AGEMA_signal_3201, rd_I_n1427}), .b ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, rd_I_n1465}), .c ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, rd_I_n1493}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U270 ( .a ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, rd_I_n1426}), .b ({state_in_s2[311], state_in_s1[311], state_in_s0[311]}), .c ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, rd_I_n1465}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U269 ( .a ({state_in_s2[55], state_in_s1[55], state_in_s0[55]}), .b ({state_in_s2[183], state_in_s1[183], state_in_s0[183]}), .c ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, rd_I_n1426}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U268 ( .a ({new_AGEMA_signal_3670, new_AGEMA_signal_3669, rd_I_n1459}), .b ({state_in_s2[101], state_in_s1[101], state_in_s0[101]}), .c ({new_AGEMA_signal_4342, new_AGEMA_signal_4341, rd_I_n2262}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U266 ( .a ({new_AGEMA_signal_3612, new_AGEMA_signal_3611, rd_I_n1424}), .b ({state_in_s2[99], state_in_s1[99], state_in_s0[99]}), .c ({new_AGEMA_signal_4344, new_AGEMA_signal_4343, rd_I_n2288}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U264 ( .a ({state_in_s2[376], state_in_s1[376], state_in_s0[376]}), .b ({new_AGEMA_signal_3604, new_AGEMA_signal_3603, rd_I_n2143}), .c ({new_AGEMA_signal_4346, new_AGEMA_signal_4345, rd_I_n2290}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U263 ( .a ({new_AGEMA_signal_3210, new_AGEMA_signal_3209, rd_I_n1423}), .b ({new_AGEMA_signal_3174, new_AGEMA_signal_3173, rd_I_n1596}), .c ({new_AGEMA_signal_3604, new_AGEMA_signal_3603, rd_I_n2143}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U262 ( .a ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, rd_I_n1422}), .b ({state_in_s2[211], state_in_s1[211], state_in_s0[211]}), .c ({new_AGEMA_signal_3174, new_AGEMA_signal_3173, rd_I_n1596}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U261 ( .a ({state_in_s2[83], state_in_s1[83], state_in_s0[83]}), .b ({state_in_s2[339], state_in_s1[339], state_in_s0[339]}), .c ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, rd_I_n1422}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U260 ( .a ({state_in_s2[195], state_in_s1[195], state_in_s0[195]}), .b ({new_AGEMA_signal_3606, new_AGEMA_signal_3605, rd_I_n1586}), .c ({new_AGEMA_signal_4348, new_AGEMA_signal_4347, rd_I_n2287}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U259 ( .a ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, rd_I_n1431}), .b ({new_AGEMA_signal_3178, new_AGEMA_signal_3177, rd_I_n1593}), .c ({new_AGEMA_signal_3606, new_AGEMA_signal_3605, rd_I_n1586}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U258 ( .a ({state_in_s2[190], state_in_s1[190], state_in_s0[190]}), .b ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, rd_I_n1421}), .c ({new_AGEMA_signal_3178, new_AGEMA_signal_3177, rd_I_n1593}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U257 ( .a ({state_in_s2[318], state_in_s1[318], state_in_s0[318]}), .b ({state_in_s2[62], state_in_s1[62], state_in_s0[62]}), .c ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, rd_I_n1421}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U256 ( .a ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, rd_I_n1420}), .b ({state_in_s2[53], state_in_s1[53], state_in_s0[53]}), .c ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, rd_I_n1431}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U255 ( .a ({state_in_s2[309], state_in_s1[309], state_in_s0[309]}), .b ({state_in_s2[181], state_in_s1[181], state_in_s0[181]}), .c ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, rd_I_n1420}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U252 ( .a ({state_in_s2[280], state_in_s1[280], state_in_s0[280]}), .b ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, rd_I_n2141}), .c ({new_AGEMA_signal_4350, new_AGEMA_signal_4349, rd_I_n2378}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U251 ( .a ({new_AGEMA_signal_3250, new_AGEMA_signal_3249, rd_I_n1418}), .b ({new_AGEMA_signal_3186, new_AGEMA_signal_3185, rd_I_n1768}), .c ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, rd_I_n2141}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U250 ( .a ({state_in_s2[371], state_in_s1[371], state_in_s0[371]}), .b ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, rd_I_n1417}), .c ({new_AGEMA_signal_3186, new_AGEMA_signal_3185, rd_I_n1768}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U249 ( .a ({state_in_s2[243], state_in_s1[243], state_in_s0[243]}), .b ({state_in_s2[115], state_in_s1[115], state_in_s0[115]}), .c ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, rd_I_n1417}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U248 ( .a ({state_in_s2[3], state_in_s1[3], state_in_s0[3]}), .b ({new_AGEMA_signal_4352, new_AGEMA_signal_4351, rd_I_n1416}), .c ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, rd_I_n2376}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U247 ( .a ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, rd_I_n1919}), .b ({1'b0, 1'b0, rc[3]}), .c ({new_AGEMA_signal_4352, new_AGEMA_signal_4351, rd_I_n1416}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U246 ( .a ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, rd_I_n1415}), .b ({new_AGEMA_signal_3190, new_AGEMA_signal_3189, rd_I_n1770}), .c ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, rd_I_n1919}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U245 ( .a ({state_in_s2[382], state_in_s1[382], state_in_s0[382]}), .b ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, rd_I_n1414}), .c ({new_AGEMA_signal_3190, new_AGEMA_signal_3189, rd_I_n1770}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U244 ( .a ({state_in_s2[126], state_in_s1[126], state_in_s0[126]}), .b ({state_in_s2[254], state_in_s1[254], state_in_s0[254]}), .c ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, rd_I_n1414}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U243 ( .a ({new_AGEMA_signal_3612, new_AGEMA_signal_3611, rd_I_n1424}), .b ({state_in_s2[227], state_in_s1[227], state_in_s0[227]}), .c ({new_AGEMA_signal_4354, new_AGEMA_signal_4353, rd_I_n2375}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U241 ( .a ({state_in_s2[355], state_in_s1[355], state_in_s0[355]}), .b ({new_AGEMA_signal_3612, new_AGEMA_signal_3611, rd_I_n1424}), .c ({new_AGEMA_signal_4356, new_AGEMA_signal_4355, rd_I_n1976}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U240 ( .a ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, rd_I_n1412}), .b ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, rd_I_n1598}), .c ({new_AGEMA_signal_3612, new_AGEMA_signal_3611, rd_I_n1424}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U239 ( .a ({state_in_s2[350], state_in_s1[350], state_in_s0[350]}), .b ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, rd_I_n1411}), .c ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, rd_I_n1598}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U238 ( .a ({state_in_s2[222], state_in_s1[222], state_in_s0[222]}), .b ({state_in_s2[94], state_in_s1[94], state_in_s0[94]}), .c ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, rd_I_n1411}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U236 ( .a ({state_in_s2[110], state_in_s1[110], state_in_s0[110]}), .b ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, rd_I_n1913}), .c ({new_AGEMA_signal_4358, new_AGEMA_signal_4357, rd_I_n1979}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U235 ( .a ({state_in_s2[206], state_in_s1[206], state_in_s0[206]}), .b ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, rd_I_n1639}), .c ({new_AGEMA_signal_4360, new_AGEMA_signal_4359, rd_I_n1978}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U234 ( .a ({new_AGEMA_signal_3202, new_AGEMA_signal_3201, rd_I_n1427}), .b ({new_AGEMA_signal_3198, new_AGEMA_signal_3197, rd_I_n1588}), .c ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, rd_I_n1639}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U233 ( .a ({state_in_s2[169], state_in_s1[169], state_in_s0[169]}), .b ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, rd_I_n1410}), .c ({new_AGEMA_signal_3198, new_AGEMA_signal_3197, rd_I_n1588}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U232 ( .a ({state_in_s2[297], state_in_s1[297], state_in_s0[297]}), .b ({state_in_s2[41], state_in_s1[41], state_in_s0[41]}), .c ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, rd_I_n1410}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U231 ( .a ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, rd_I_n1409}), .b ({state_in_s2[160], state_in_s1[160], state_in_s0[160]}), .c ({new_AGEMA_signal_3202, new_AGEMA_signal_3201, rd_I_n1427}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U230 ( .a ({state_in_s2[288], state_in_s1[288], state_in_s0[288]}), .b ({state_in_s2[32], state_in_s1[32], state_in_s0[32]}), .c ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, rd_I_n1409}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U227 ( .a ({state_in_s2[239], state_in_s1[239], state_in_s0[239]}), .b ({new_AGEMA_signal_3616, new_AGEMA_signal_3615, rd_I_n1724}), .c ({new_AGEMA_signal_4362, new_AGEMA_signal_4361, rd_I_n2294}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U226 ( .a ({new_AGEMA_signal_3210, new_AGEMA_signal_3209, rd_I_n1423}), .b ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, rd_I_n1438}), .c ({new_AGEMA_signal_3616, new_AGEMA_signal_3615, rd_I_n1724}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U225 ( .a ({state_in_s2[65], state_in_s1[65], state_in_s0[65]}), .b ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, rd_I_n1407}), .c ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, rd_I_n1438}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U224 ( .a ({state_in_s2[321], state_in_s1[321], state_in_s0[321]}), .b ({state_in_s2[193], state_in_s1[193], state_in_s0[193]}), .c ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, rd_I_n1407}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U223 ( .a ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, rd_I_n1406}), .b ({state_in_s2[74], state_in_s1[74], state_in_s0[74]}), .c ({new_AGEMA_signal_3210, new_AGEMA_signal_3209, rd_I_n1423}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U222 ( .a ({state_in_s2[202], state_in_s1[202], state_in_s0[202]}), .b ({state_in_s2[330], state_in_s1[330], state_in_s0[330]}), .c ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, rd_I_n1406}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U221 ( .a ({state_in_s2[260], state_in_s1[260], state_in_s0[260]}), .b ({new_AGEMA_signal_3618, new_AGEMA_signal_3617, rd_I_n1834}), .c ({new_AGEMA_signal_4364, new_AGEMA_signal_4363, rd_I_n2292}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U220 ( .a ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, rd_I_n1788}), .b ({new_AGEMA_signal_3214, new_AGEMA_signal_3213, rd_I_n1441}), .c ({new_AGEMA_signal_3618, new_AGEMA_signal_3617, rd_I_n1834}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U219 ( .a ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, rd_I_n1405}), .b ({state_in_s2[374], state_in_s1[374], state_in_s0[374]}), .c ({new_AGEMA_signal_3214, new_AGEMA_signal_3213, rd_I_n1441}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U218 ( .a ({state_in_s2[246], state_in_s1[246], state_in_s0[246]}), .b ({state_in_s2[118], state_in_s1[118], state_in_s0[118]}), .c ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, rd_I_n1405}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U217 ( .a ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, rd_I_n1404}), .b ({state_in_s2[127], state_in_s1[127], state_in_s0[127]}), .c ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, rd_I_n1788}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U216 ( .a ({state_in_s2[255], state_in_s1[255], state_in_s0[255]}), .b ({state_in_s2[383], state_in_s1[383], state_in_s0[383]}), .c ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, rd_I_n1404}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U215 ( .a ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, rd_I_n1403}), .b ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, rd_I_n1402}), .c ({new_AGEMA_signal_4366, new_AGEMA_signal_4365, rd_I_n2291}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U214 ( .a ({state_in_s2[15], state_in_s1[15], state_in_s0[15]}), .b ({1'b0, 1'b0, rc[15]}), .c ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, rd_I_n1402}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U211 ( .a ({state_in_s2[292], state_in_s1[292], state_in_s0[292]}), .b ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, rd_I_n2215}), .c ({new_AGEMA_signal_4368, new_AGEMA_signal_4367, rd_I_n2269}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U210 ( .a ({new_AGEMA_signal_3226, new_AGEMA_signal_3225, rd_I_n1698}), .b ({new_AGEMA_signal_3222, new_AGEMA_signal_3221, rd_I_n1719}), .c ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, rd_I_n2215}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U209 ( .a ({state_in_s2[287], state_in_s1[287], state_in_s0[287]}), .b ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, rd_I_n1400}), .c ({new_AGEMA_signal_3222, new_AGEMA_signal_3221, rd_I_n1719}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U208 ( .a ({state_in_s2[31], state_in_s1[31], state_in_s0[31]}), .b ({state_in_s2[159], state_in_s1[159], state_in_s0[159]}), .c ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, rd_I_n1400}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U207 ( .a ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, rd_I_n1399}), .b ({state_in_s2[278], state_in_s1[278], state_in_s0[278]}), .c ({new_AGEMA_signal_3226, new_AGEMA_signal_3225, rd_I_n1698}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U206 ( .a ({state_in_s2[22], state_in_s1[22], state_in_s0[22]}), .b ({state_in_s2[150], state_in_s1[150], state_in_s0[150]}), .c ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, rd_I_n1399}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U205 ( .a ({state_in_s2[47], state_in_s1[47], state_in_s0[47]}), .b ({new_AGEMA_signal_3622, new_AGEMA_signal_3621, rd_I_n1793}), .c ({new_AGEMA_signal_4370, new_AGEMA_signal_4369, rd_I_n2267}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U204 ( .a ({new_AGEMA_signal_3234, new_AGEMA_signal_3233, rd_I_n1716}), .b ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, rd_I_n1701}), .c ({new_AGEMA_signal_3622, new_AGEMA_signal_3621, rd_I_n1793}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U203 ( .a ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, rd_I_n1398}), .b ({state_in_s2[257], state_in_s1[257], state_in_s0[257]}), .c ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, rd_I_n1701}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U202 ( .a ({state_in_s2[1], state_in_s1[1], state_in_s0[1]}), .b ({state_in_s2[129], state_in_s1[129], state_in_s0[129]}), .c ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, rd_I_n1398}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U201 ( .a ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, rd_I_n1397}), .b ({state_in_s2[138], state_in_s1[138], state_in_s0[138]}), .c ({new_AGEMA_signal_3234, new_AGEMA_signal_3233, rd_I_n1716}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U200 ( .a ({state_in_s2[10], state_in_s1[10], state_in_s0[10]}), .b ({state_in_s2[266], state_in_s1[266], state_in_s0[266]}), .c ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, rd_I_n1397}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U199 ( .a ({state_in_s2[143], state_in_s1[143], state_in_s0[143]}), .b ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, rd_I_n1403}), .c ({new_AGEMA_signal_4372, new_AGEMA_signal_4371, rd_I_n2266}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U196 ( .a ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, rd_I_n1395}), .b ({new_AGEMA_signal_3672, new_AGEMA_signal_3671, rd_I_n1794}), .c ({new_AGEMA_signal_4374, new_AGEMA_signal_4373, rd_I_n2001}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U195 ( .a ({state_in_s2[26], state_in_s1[26], state_in_s0[26]}), .b ({1'b0, 1'b0, rc[26]}), .c ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, rd_I_n1395}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U194 ( .a ({state_in_s2[250], state_in_s1[250], state_in_s0[250]}), .b ({new_AGEMA_signal_3624, new_AGEMA_signal_3623, rd_I_n1432}), .c ({new_AGEMA_signal_4376, new_AGEMA_signal_4375, rd_I_n1999}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U193 ( .a ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, rd_I_n1412}), .b ({new_AGEMA_signal_3238, new_AGEMA_signal_3237, rd_I_n1435}), .c ({new_AGEMA_signal_3624, new_AGEMA_signal_3623, rd_I_n1432}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U192 ( .a ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, rd_I_n1394}), .b ({state_in_s2[76], state_in_s1[76], state_in_s0[76]}), .c ({new_AGEMA_signal_3238, new_AGEMA_signal_3237, rd_I_n1435}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U191 ( .a ({state_in_s2[332], state_in_s1[332], state_in_s0[332]}), .b ({state_in_s2[204], state_in_s1[204], state_in_s0[204]}), .c ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, rd_I_n1394}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U190 ( .a ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, rd_I_n1393}), .b ({state_in_s2[85], state_in_s1[85], state_in_s0[85]}), .c ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, rd_I_n1412}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U189 ( .a ({state_in_s2[213], state_in_s1[213], state_in_s0[213]}), .b ({state_in_s2[341], state_in_s1[341], state_in_s0[341]}), .c ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, rd_I_n1393}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U188 ( .a ({state_in_s2[271], state_in_s1[271], state_in_s0[271]}), .b ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, rd_I_n1403}), .c ({new_AGEMA_signal_4378, new_AGEMA_signal_4377, rd_I_n1998}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U187 ( .a ({new_AGEMA_signal_3250, new_AGEMA_signal_3249, rd_I_n1418}), .b ({new_AGEMA_signal_3246, new_AGEMA_signal_3245, rd_I_n1443}), .c ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, rd_I_n1403}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U186 ( .a ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, rd_I_n1392}), .b ({state_in_s2[97], state_in_s1[97], state_in_s0[97]}), .c ({new_AGEMA_signal_3246, new_AGEMA_signal_3245, rd_I_n1443}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U185 ( .a ({state_in_s2[225], state_in_s1[225], state_in_s0[225]}), .b ({state_in_s2[353], state_in_s1[353], state_in_s0[353]}), .c ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, rd_I_n1392}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U184 ( .a ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, rd_I_n1391}), .b ({state_in_s2[106], state_in_s1[106], state_in_s0[106]}), .c ({new_AGEMA_signal_3250, new_AGEMA_signal_3249, rd_I_n1418}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U183 ( .a ({state_in_s2[234], state_in_s1[234], state_in_s0[234]}), .b ({state_in_s2[362], state_in_s1[362], state_in_s0[362]}), .c ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, rd_I_n1391}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U181 ( .a ({new_AGEMA_signal_3640, new_AGEMA_signal_3639, rd_I_n1389}), .b ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, rd_I_n1388}), .c ({new_AGEMA_signal_4380, new_AGEMA_signal_4379, rd_I_n1777}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U180 ( .a ({state_in_s2[18], state_in_s1[18], state_in_s0[18]}), .b ({1'b0, 1'b0, rc[18]}), .c ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, rd_I_n1388}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U178 ( .a ({state_in_s2[263], state_in_s1[263], state_in_s0[263]}), .b ({new_AGEMA_signal_3628, new_AGEMA_signal_3627, rd_I_n1633}), .c ({new_AGEMA_signal_4382, new_AGEMA_signal_4381, rd_I_n1778}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U177 ( .a ({new_AGEMA_signal_3406, new_AGEMA_signal_3405, rd_I_n1387}), .b ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, rd_I_n1507}), .c ({new_AGEMA_signal_3628, new_AGEMA_signal_3627, rd_I_n1633}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U176 ( .a ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, rd_I_n1386}), .b ({state_in_s2[121], state_in_s1[121], state_in_s0[121]}), .c ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, rd_I_n1507}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U175 ( .a ({state_in_s2[377], state_in_s1[377], state_in_s0[377]}), .b ({state_in_s2[249], state_in_s1[249], state_in_s0[249]}), .c ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, rd_I_n1386}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U174 ( .a ({state_in_s2[242], state_in_s1[242], state_in_s0[242]}), .b ({new_AGEMA_signal_3630, new_AGEMA_signal_3629, rd_I_n1734}), .c ({new_AGEMA_signal_4384, new_AGEMA_signal_4383, rd_I_n1780}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U173 ( .a ({new_AGEMA_signal_3262, new_AGEMA_signal_3261, rd_I_n1505}), .b ({new_AGEMA_signal_3258, new_AGEMA_signal_3257, rd_I_n1448}), .c ({new_AGEMA_signal_3630, new_AGEMA_signal_3629, rd_I_n1734}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U172 ( .a ({state_in_s2[77], state_in_s1[77], state_in_s0[77]}), .b ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, rd_I_n1385}), .c ({new_AGEMA_signal_3258, new_AGEMA_signal_3257, rd_I_n1448}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U171 ( .a ({state_in_s2[205], state_in_s1[205], state_in_s0[205]}), .b ({state_in_s2[333], state_in_s1[333], state_in_s0[333]}), .c ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, rd_I_n1385}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U170 ( .a ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, rd_I_n1384}), .b ({state_in_s2[68], state_in_s1[68], state_in_s0[68]}), .c ({new_AGEMA_signal_3262, new_AGEMA_signal_3261, rd_I_n1505}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U169 ( .a ({state_in_s2[196], state_in_s1[196], state_in_s0[196]}), .b ({state_in_s2[324], state_in_s1[324], state_in_s0[324]}), .c ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, rd_I_n1384}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U166 ( .a ({state_in_s2[295], state_in_s1[295], state_in_s0[295]}), .b ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, rd_I_n1630}), .c ({new_AGEMA_signal_4386, new_AGEMA_signal_4385, rd_I_n2408}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U165 ( .a ({new_AGEMA_signal_3270, new_AGEMA_signal_3269, rd_I_n1512}), .b ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, rd_I_n1490}), .c ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, rd_I_n1630}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U164 ( .a ({state_in_s2[258], state_in_s1[258], state_in_s0[258]}), .b ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, rd_I_n1382}), .c ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, rd_I_n1490}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U163 ( .a ({state_in_s2[2], state_in_s1[2], state_in_s0[2]}), .b ({state_in_s2[130], state_in_s1[130], state_in_s0[130]}), .c ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, rd_I_n1382}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U162 ( .a ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, rd_I_n1381}), .b ({state_in_s2[281], state_in_s1[281], state_in_s0[281]}), .c ({new_AGEMA_signal_3270, new_AGEMA_signal_3269, rd_I_n1512}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U161 ( .a ({state_in_s2[25], state_in_s1[25], state_in_s0[25]}), .b ({state_in_s2[153], state_in_s1[153], state_in_s0[153]}), .c ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, rd_I_n1381}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U160 ( .a ({state_in_s2[50], state_in_s1[50], state_in_s0[50]}), .b ({new_AGEMA_signal_3634, new_AGEMA_signal_3633, rd_I_n1989}), .c ({new_AGEMA_signal_4388, new_AGEMA_signal_4387, rd_I_n2406}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U159 ( .a ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, rd_I_n1532}), .b ({new_AGEMA_signal_3274, new_AGEMA_signal_3273, rd_I_n1699}), .c ({new_AGEMA_signal_3634, new_AGEMA_signal_3633, rd_I_n1989}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U158 ( .a ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, rd_I_n1380}), .b ({state_in_s2[13], state_in_s1[13], state_in_s0[13]}), .c ({new_AGEMA_signal_3274, new_AGEMA_signal_3273, rd_I_n1699}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U157 ( .a ({state_in_s2[141], state_in_s1[141], state_in_s0[141]}), .b ({state_in_s2[269], state_in_s1[269], state_in_s0[269]}), .c ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, rd_I_n1380}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U156 ( .a ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, rd_I_n1379}), .b ({state_in_s2[132], state_in_s1[132], state_in_s0[132]}), .c ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, rd_I_n1532}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U155 ( .a ({state_in_s2[4], state_in_s1[4], state_in_s0[4]}), .b ({state_in_s2[260], state_in_s1[260], state_in_s0[260]}), .c ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, rd_I_n1379}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U154 ( .a ({state_in_s2[146], state_in_s1[146], state_in_s0[146]}), .b ({new_AGEMA_signal_3640, new_AGEMA_signal_3639, rd_I_n1389}), .c ({new_AGEMA_signal_4390, new_AGEMA_signal_4389, rd_I_n2405}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U151 ( .a ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, rd_I_n1377}), .b ({new_AGEMA_signal_3636, new_AGEMA_signal_3635, rd_I_n1988}), .c ({new_AGEMA_signal_4392, new_AGEMA_signal_4391, rd_I_n1994}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U150 ( .a ({new_AGEMA_signal_3286, new_AGEMA_signal_3285, rd_I_n1673}), .b ({new_AGEMA_signal_3282, new_AGEMA_signal_3281, rd_I_n1444}), .c ({new_AGEMA_signal_3636, new_AGEMA_signal_3635, rd_I_n1988}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U149 ( .a ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, rd_I_n1376}), .b ({state_in_s2[120], state_in_s1[120], state_in_s0[120]}), .c ({new_AGEMA_signal_3282, new_AGEMA_signal_3281, rd_I_n1444}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U148 ( .a ({state_in_s2[376], state_in_s1[376], state_in_s0[376]}), .b ({state_in_s2[248], state_in_s1[248], state_in_s0[248]}), .c ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, rd_I_n1376}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U147 ( .a ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, rd_I_n1375}), .b ({state_in_s2[239], state_in_s1[239], state_in_s0[239]}), .c ({new_AGEMA_signal_3286, new_AGEMA_signal_3285, rd_I_n1673}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U146 ( .a ({state_in_s2[367], state_in_s1[367], state_in_s0[367]}), .b ({state_in_s2[111], state_in_s1[111], state_in_s0[111]}), .c ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, rd_I_n1375}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U145 ( .a ({state_in_s2[29], state_in_s1[29], state_in_s0[29]}), .b ({1'b0, 1'b0, rc[29]}), .c ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, rd_I_n1377}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U144 ( .a ({state_in_s2[253], state_in_s1[253], state_in_s0[253]}), .b ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, rd_I_n1499}), .c ({new_AGEMA_signal_4394, new_AGEMA_signal_4393, rd_I_n1992}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U143 ( .a ({new_AGEMA_signal_3294, new_AGEMA_signal_3293, rd_I_n1536}), .b ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, rd_I_n1439}), .c ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, rd_I_n1499}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U142 ( .a ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, rd_I_n1374}), .b ({state_in_s2[88], state_in_s1[88], state_in_s0[88]}), .c ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, rd_I_n1439}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U141 ( .a ({state_in_s2[216], state_in_s1[216], state_in_s0[216]}), .b ({state_in_s2[344], state_in_s1[344], state_in_s0[344]}), .c ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, rd_I_n1374}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U140 ( .a ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, rd_I_n1373}), .b ({state_in_s2[207], state_in_s1[207], state_in_s0[207]}), .c ({new_AGEMA_signal_3294, new_AGEMA_signal_3293, rd_I_n1536}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U139 ( .a ({state_in_s2[335], state_in_s1[335], state_in_s0[335]}), .b ({state_in_s2[79], state_in_s1[79], state_in_s0[79]}), .c ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, rd_I_n1373}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U138 ( .a ({state_in_s2[274], state_in_s1[274], state_in_s0[274]}), .b ({new_AGEMA_signal_3640, new_AGEMA_signal_3639, rd_I_n1389}), .c ({new_AGEMA_signal_4396, new_AGEMA_signal_4395, rd_I_n1991}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U137 ( .a ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, rd_I_n1502}), .b ({new_AGEMA_signal_3298, new_AGEMA_signal_3297, rd_I_n1442}), .c ({new_AGEMA_signal_3640, new_AGEMA_signal_3639, rd_I_n1389}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U136 ( .a ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, rd_I_n1372}), .b ({state_in_s2[237], state_in_s1[237], state_in_s0[237]}), .c ({new_AGEMA_signal_3298, new_AGEMA_signal_3297, rd_I_n1442}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U135 ( .a ({state_in_s2[109], state_in_s1[109], state_in_s0[109]}), .b ({state_in_s2[365], state_in_s1[365], state_in_s0[365]}), .c ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, rd_I_n1372}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U134 ( .a ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, rd_I_n1371}), .b ({state_in_s2[356], state_in_s1[356], state_in_s0[356]}), .c ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, rd_I_n1502}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U133 ( .a ({state_in_s2[100], state_in_s1[100], state_in_s0[100]}), .b ({state_in_s2[228], state_in_s1[228], state_in_s0[228]}), .c ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, rd_I_n1371}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U131 ( .a ({state_in_s2[98], state_in_s1[98], state_in_s0[98]}), .b ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, rd_I_n1369}), .c ({new_AGEMA_signal_4398, new_AGEMA_signal_4397, rd_I_n2112}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U129 ( .a ({state_in_s2[375], state_in_s1[375], state_in_s0[375]}), .b ({new_AGEMA_signal_3642, new_AGEMA_signal_3641, rd_I_n1917}), .c ({new_AGEMA_signal_4400, new_AGEMA_signal_4399, rd_I_n2113}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U128 ( .a ({new_AGEMA_signal_3334, new_AGEMA_signal_3333, rd_I_n1368}), .b ({new_AGEMA_signal_3306, new_AGEMA_signal_3305, rd_I_n1569}), .c ({new_AGEMA_signal_3642, new_AGEMA_signal_3641, rd_I_n1917}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U127 ( .a ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, rd_I_n1367}), .b ({state_in_s2[338], state_in_s1[338], state_in_s0[338]}), .c ({new_AGEMA_signal_3306, new_AGEMA_signal_3305, rd_I_n1569}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U126 ( .a ({state_in_s2[82], state_in_s1[82], state_in_s0[82]}), .b ({state_in_s2[210], state_in_s1[210], state_in_s0[210]}), .c ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, rd_I_n1367}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U125 ( .a ({state_in_s2[194], state_in_s1[194], state_in_s0[194]}), .b ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, rd_I_n1951}), .c ({new_AGEMA_signal_4402, new_AGEMA_signal_4401, rd_I_n2115}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U124 ( .a ({new_AGEMA_signal_3310, new_AGEMA_signal_3309, rd_I_n1564}), .b ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, rd_I_n1366}), .c ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, rd_I_n1951}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U123 ( .a ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, rd_I_n1365}), .b ({state_in_s2[189], state_in_s1[189], state_in_s0[189]}), .c ({new_AGEMA_signal_3310, new_AGEMA_signal_3309, rd_I_n1564}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U122 ( .a ({state_in_s2[317], state_in_s1[317], state_in_s0[317]}), .b ({state_in_s2[61], state_in_s1[61], state_in_s0[61]}), .c ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, rd_I_n1365}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U119 ( .a ({state_in_s2[279], state_in_s1[279], state_in_s0[279]}), .b ({new_AGEMA_signal_3646, new_AGEMA_signal_3645, rd_I_n1915}), .c ({new_AGEMA_signal_4404, new_AGEMA_signal_4403, rd_I_n2498}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U118 ( .a ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, rd_I_n1665}), .b ({new_AGEMA_signal_3346, new_AGEMA_signal_3345, rd_I_n1363}), .c ({new_AGEMA_signal_3646, new_AGEMA_signal_3645, rd_I_n1915}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U117 ( .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, rd_I_n1362}), .b ({state_in_s2[370], state_in_s1[370], state_in_s0[370]}), .c ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, rd_I_n1665}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U116 ( .a ({state_in_s2[242], state_in_s1[242], state_in_s0[242]}), .b ({state_in_s2[114], state_in_s1[114], state_in_s0[114]}), .c ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, rd_I_n1362}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U115 ( .a ({new_AGEMA_signal_3648, new_AGEMA_signal_3647, rd_I_n1786}), .b ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, rd_I_n1361}), .c ({new_AGEMA_signal_4406, new_AGEMA_signal_4405, rd_I_n2496}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U114 ( .a ({1'b0, 1'b0, rc[2]}), .b ({state_in_s2[2], state_in_s1[2], state_in_s0[2]}), .c ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, rd_I_n1361}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U113 ( .a ({new_AGEMA_signal_3318, new_AGEMA_signal_3317, rd_I_n1667}), .b ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, rd_I_n1360}), .c ({new_AGEMA_signal_3648, new_AGEMA_signal_3647, rd_I_n1786}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U112 ( .a ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, rd_I_n1359}), .b ({state_in_s2[253], state_in_s1[253], state_in_s0[253]}), .c ({new_AGEMA_signal_3318, new_AGEMA_signal_3317, rd_I_n1667}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U111 ( .a ({state_in_s2[381], state_in_s1[381], state_in_s0[381]}), .b ({state_in_s2[125], state_in_s1[125], state_in_s0[125]}), .c ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, rd_I_n1359}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U110 ( .a ({state_in_s2[226], state_in_s1[226], state_in_s0[226]}), .b ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, rd_I_n1369}), .c ({new_AGEMA_signal_4408, new_AGEMA_signal_4407, rd_I_n2495}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U108 ( .a ({state_in_s2[354], state_in_s1[354], state_in_s0[354]}), .b ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, rd_I_n1369}), .c ({new_AGEMA_signal_4410, new_AGEMA_signal_4409, rd_I_n1815}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U107 ( .a ({new_AGEMA_signal_3354, new_AGEMA_signal_3353, rd_I_n1357}), .b ({new_AGEMA_signal_3322, new_AGEMA_signal_3321, rd_I_n1567}), .c ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, rd_I_n1369}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U106 ( .a ({state_in_s2[93], state_in_s1[93], state_in_s0[93]}), .b ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, rd_I_n1356}), .c ({new_AGEMA_signal_3322, new_AGEMA_signal_3321, rd_I_n1567}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U105 ( .a ({state_in_s2[221], state_in_s1[221], state_in_s0[221]}), .b ({state_in_s2[349], state_in_s1[349], state_in_s0[349]}), .c ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, rd_I_n1356}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U103 ( .a ({state_in_s2[205], state_in_s1[205], state_in_s0[205]}), .b ({new_AGEMA_signal_3652, new_AGEMA_signal_3651, rd_I_n1721}), .c ({new_AGEMA_signal_4412, new_AGEMA_signal_4411, rd_I_n1816}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U102 ( .a ({new_AGEMA_signal_3366, new_AGEMA_signal_3365, rd_I_n1355}), .b ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, rd_I_n1559}), .c ({new_AGEMA_signal_3652, new_AGEMA_signal_3651, rd_I_n1721}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U101 ( .a ({state_in_s2[296], state_in_s1[296], state_in_s0[296]}), .b ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, rd_I_n1354}), .c ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, rd_I_n1559}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U100 ( .a ({state_in_s2[40], state_in_s1[40], state_in_s0[40]}), .b ({state_in_s2[168], state_in_s1[168], state_in_s0[168]}), .c ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, rd_I_n1354}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U99 ( .a ({state_in_s2[109], state_in_s1[109], state_in_s0[109]}), .b ({new_AGEMA_signal_3654, new_AGEMA_signal_3653, rd_I_n1811}), .c ({new_AGEMA_signal_4414, new_AGEMA_signal_4413, rd_I_n1818}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U98 ( .a ({new_AGEMA_signal_3358, new_AGEMA_signal_3357, rd_I_n1353}), .b ({new_AGEMA_signal_3330, new_AGEMA_signal_3329, rd_I_n1661}), .c ({new_AGEMA_signal_3654, new_AGEMA_signal_3653, rd_I_n1811}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U97 ( .a ({state_in_s2[328], state_in_s1[328], state_in_s0[328]}), .b ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, rd_I_n1352}), .c ({new_AGEMA_signal_3330, new_AGEMA_signal_3329, rd_I_n1661}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U96 ( .a ({state_in_s2[200], state_in_s1[200], state_in_s0[200]}), .b ({state_in_s2[72], state_in_s1[72], state_in_s0[72]}), .c ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, rd_I_n1352}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U94 ( .a ({new_AGEMA_signal_3664, new_AGEMA_signal_3663, rd_I_n1350}), .b ({state_in_s2[121], state_in_s1[121], state_in_s0[121]}), .c ({new_AGEMA_signal_4416, new_AGEMA_signal_4415, rd_I_n2220}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U92 ( .a ({state_in_s2[366], state_in_s1[366], state_in_s0[366]}), .b ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, rd_I_n1913}), .c ({new_AGEMA_signal_4418, new_AGEMA_signal_4417, rd_I_n2221}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U91 ( .a ({new_AGEMA_signal_3378, new_AGEMA_signal_3377, rd_I_n1349}), .b ({new_AGEMA_signal_3334, new_AGEMA_signal_3333, rd_I_n1368}), .c ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, rd_I_n1913}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U90 ( .a ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, rd_I_n1348}), .b ({state_in_s2[73], state_in_s1[73], state_in_s0[73]}), .c ({new_AGEMA_signal_3334, new_AGEMA_signal_3333, rd_I_n1368}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U89 ( .a ({state_in_s2[201], state_in_s1[201], state_in_s0[201]}), .b ({state_in_s2[329], state_in_s1[329], state_in_s0[329]}), .c ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, rd_I_n1348}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U88 ( .a ({state_in_s2[217], state_in_s1[217], state_in_s0[217]}), .b ({new_AGEMA_signal_3658, new_AGEMA_signal_3657, rd_I_n2214}), .c ({new_AGEMA_signal_4420, new_AGEMA_signal_4419, rd_I_n2223}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U87 ( .a ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, rd_I_n1458}), .b ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, rd_I_n1366}), .c ({new_AGEMA_signal_3658, new_AGEMA_signal_3657, rd_I_n2214}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U86 ( .a ({state_in_s2[180], state_in_s1[180], state_in_s0[180]}), .b ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, rd_I_n1347}), .c ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, rd_I_n1366}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U85 ( .a ({state_in_s2[308], state_in_s1[308], state_in_s0[308]}), .b ({state_in_s2[52], state_in_s1[52], state_in_s0[52]}), .c ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, rd_I_n1347}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U84 ( .a ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, rd_I_n1346}), .b ({state_in_s2[171], state_in_s1[171], state_in_s0[171]}), .c ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, rd_I_n1458}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U83 ( .a ({state_in_s2[299], state_in_s1[299], state_in_s0[299]}), .b ({state_in_s2[43], state_in_s1[43], state_in_s0[43]}), .c ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, rd_I_n1346}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U80 ( .a ({new_AGEMA_signal_3660, new_AGEMA_signal_3659, rd_I_n1911}), .b ({state_in_s2[270], state_in_s1[270], state_in_s0[270]}), .c ({new_AGEMA_signal_4422, new_AGEMA_signal_4421, rd_I_n2493}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U79 ( .a ({new_AGEMA_signal_3426, new_AGEMA_signal_3425, rd_I_n1344}), .b ({new_AGEMA_signal_3346, new_AGEMA_signal_3345, rd_I_n1363}), .c ({new_AGEMA_signal_3660, new_AGEMA_signal_3659, rd_I_n1911}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U78 ( .a ({state_in_s2[233], state_in_s1[233], state_in_s0[233]}), .b ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, rd_I_n1343}), .c ({new_AGEMA_signal_3346, new_AGEMA_signal_3345, rd_I_n1363}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U77 ( .a ({state_in_s2[105], state_in_s1[105], state_in_s0[105]}), .b ({state_in_s2[361], state_in_s1[361], state_in_s0[361]}), .c ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, rd_I_n1343}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U76 ( .a ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, rd_I_n1652}), .b ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, rd_I_n1342}), .c ({new_AGEMA_signal_4424, new_AGEMA_signal_4423, rd_I_n2491}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U75 ( .a ({1'b0, 1'b0, rc[25]}), .b ({state_in_s2[25], state_in_s1[25], state_in_s0[25]}), .c ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, rd_I_n1342}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U74 ( .a ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, rd_I_n1341}), .b ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, rd_I_n1360}), .c ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, rd_I_n1652}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U73 ( .a ({state_in_s2[372], state_in_s1[372], state_in_s0[372]}), .b ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, rd_I_n1340}), .c ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, rd_I_n1360}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U72 ( .a ({state_in_s2[244], state_in_s1[244], state_in_s0[244]}), .b ({state_in_s2[116], state_in_s1[116], state_in_s0[116]}), .c ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, rd_I_n1340}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U71 ( .a ({new_AGEMA_signal_3664, new_AGEMA_signal_3663, rd_I_n1350}), .b ({state_in_s2[249], state_in_s1[249], state_in_s0[249]}), .c ({new_AGEMA_signal_4426, new_AGEMA_signal_4425, rd_I_n2490}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U69 ( .a ({state_in_s2[377], state_in_s1[377], state_in_s0[377]}), .b ({new_AGEMA_signal_3664, new_AGEMA_signal_3663, rd_I_n1350}), .c ({new_AGEMA_signal_4428, new_AGEMA_signal_4427, rd_I_n2454}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U68 ( .a ({new_AGEMA_signal_3418, new_AGEMA_signal_3417, rd_I_n1338}), .b ({new_AGEMA_signal_3354, new_AGEMA_signal_3353, rd_I_n1357}), .c ({new_AGEMA_signal_3664, new_AGEMA_signal_3663, rd_I_n1350}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U67 ( .a ({state_in_s2[84], state_in_s1[84], state_in_s0[84]}), .b ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, rd_I_n1337}), .c ({new_AGEMA_signal_3354, new_AGEMA_signal_3353, rd_I_n1357}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U66 ( .a ({state_in_s2[212], state_in_s1[212], state_in_s0[212]}), .b ({state_in_s2[340], state_in_s1[340], state_in_s0[340]}), .c ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, rd_I_n1337}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U64 ( .a ({state_in_s2[100], state_in_s1[100], state_in_s0[100]}), .b ({new_AGEMA_signal_3666, new_AGEMA_signal_3665, rd_I_n1723}), .c ({new_AGEMA_signal_4430, new_AGEMA_signal_4429, rd_I_n2453}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U63 ( .a ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, rd_I_n1449}), .b ({new_AGEMA_signal_3358, new_AGEMA_signal_3357, rd_I_n1353}), .c ({new_AGEMA_signal_3666, new_AGEMA_signal_3665, rd_I_n1723}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U62 ( .a ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, rd_I_n1336}), .b ({state_in_s2[351], state_in_s1[351], state_in_s0[351]}), .c ({new_AGEMA_signal_3358, new_AGEMA_signal_3357, rd_I_n1353}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U61 ( .a ({state_in_s2[223], state_in_s1[223], state_in_s0[223]}), .b ({state_in_s2[95], state_in_s1[95], state_in_s0[95]}), .c ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, rd_I_n1336}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U60 ( .a ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, rd_I_n1335}), .b ({state_in_s2[86], state_in_s1[86], state_in_s0[86]}), .c ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, rd_I_n1449}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U59 ( .a ({state_in_s2[214], state_in_s1[214], state_in_s0[214]}), .b ({state_in_s2[342], state_in_s1[342], state_in_s0[342]}), .c ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, rd_I_n1335}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U58 ( .a ({state_in_s2[196], state_in_s1[196], state_in_s0[196]}), .b ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, rd_I_n2216}), .c ({new_AGEMA_signal_4432, new_AGEMA_signal_4431, rd_I_n2456}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U57 ( .a ({new_AGEMA_signal_3370, new_AGEMA_signal_3369, rd_I_n1454}), .b ({new_AGEMA_signal_3366, new_AGEMA_signal_3365, rd_I_n1355}), .c ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, rd_I_n2216}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U56 ( .a ({state_in_s2[191], state_in_s1[191], state_in_s0[191]}), .b ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, rd_I_n1334}), .c ({new_AGEMA_signal_3366, new_AGEMA_signal_3365, rd_I_n1355}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U55 ( .a ({state_in_s2[63], state_in_s1[63], state_in_s0[63]}), .b ({state_in_s2[319], state_in_s1[319], state_in_s0[319]}), .c ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, rd_I_n1334}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U54 ( .a ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, rd_I_n1333}), .b ({state_in_s2[182], state_in_s1[182], state_in_s0[182]}), .c ({new_AGEMA_signal_3370, new_AGEMA_signal_3369, rd_I_n1454}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U53 ( .a ({state_in_s2[54], state_in_s1[54], state_in_s0[54]}), .b ({state_in_s2[310], state_in_s1[310], state_in_s0[310]}), .c ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, rd_I_n1333}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U50 ( .a ({state_in_s2[229], state_in_s1[229], state_in_s0[229]}), .b ({new_AGEMA_signal_3670, new_AGEMA_signal_3669, rd_I_n1459}), .c ({new_AGEMA_signal_4434, new_AGEMA_signal_4433, rd_I_n2257}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U49 ( .a ({new_AGEMA_signal_3378, new_AGEMA_signal_3377, rd_I_n1349}), .b ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, rd_I_n1463}), .c ({new_AGEMA_signal_3670, new_AGEMA_signal_3669, rd_I_n1459}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U48 ( .a ({state_in_s2[215], state_in_s1[215], state_in_s0[215]}), .b ({new_AGEMA_signal_2842, new_AGEMA_signal_2841, rd_I_n1331}), .c ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, rd_I_n1463}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U47 ( .a ({state_in_s2[87], state_in_s1[87], state_in_s0[87]}), .b ({state_in_s2[343], state_in_s1[343], state_in_s0[343]}), .c ({new_AGEMA_signal_2842, new_AGEMA_signal_2841, rd_I_n1331}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U46 ( .a ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, rd_I_n1330}), .b ({state_in_s2[64], state_in_s1[64], state_in_s0[64]}), .c ({new_AGEMA_signal_3378, new_AGEMA_signal_3377, rd_I_n1349}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U45 ( .a ({state_in_s2[192], state_in_s1[192], state_in_s0[192]}), .b ({state_in_s2[320], state_in_s1[320], state_in_s0[320]}), .c ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, rd_I_n1330}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U44 ( .a ({state_in_s2[282], state_in_s1[282], state_in_s0[282]}), .b ({new_AGEMA_signal_3672, new_AGEMA_signal_3671, rd_I_n1794}), .c ({new_AGEMA_signal_4436, new_AGEMA_signal_4435, rd_I_n2255}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U43 ( .a ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, rd_I_n1415}), .b ({new_AGEMA_signal_3382, new_AGEMA_signal_3381, rd_I_n1480}), .c ({new_AGEMA_signal_3672, new_AGEMA_signal_3671, rd_I_n1794}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U42 ( .a ({new_AGEMA_signal_2854, new_AGEMA_signal_2853, rd_I_n1329}), .b ({state_in_s2[108], state_in_s1[108], state_in_s0[108]}), .c ({new_AGEMA_signal_3382, new_AGEMA_signal_3381, rd_I_n1480}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U41 ( .a ({state_in_s2[236], state_in_s1[236], state_in_s0[236]}), .b ({state_in_s2[364], state_in_s1[364], state_in_s0[364]}), .c ({new_AGEMA_signal_2854, new_AGEMA_signal_2853, rd_I_n1329}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U40 ( .a ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, rd_I_n1328}), .b ({state_in_s2[373], state_in_s1[373], state_in_s0[373]}), .c ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, rd_I_n1415}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U39 ( .a ({state_in_s2[117], state_in_s1[117], state_in_s0[117]}), .b ({state_in_s2[245], state_in_s1[245], state_in_s0[245]}), .c ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, rd_I_n1328}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U38 ( .a ({new_AGEMA_signal_3682, new_AGEMA_signal_3681, rd_I_n1327}), .b ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, rd_I_n1326}), .c ({new_AGEMA_signal_4438, new_AGEMA_signal_4437, rd_I_n2254}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U37 ( .a ({state_in_s2[5], state_in_s1[5], state_in_s0[5]}), .b ({1'b0, 1'b0, rc[5]}), .c ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, rd_I_n1326}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U34 ( .a ({state_in_s2[314], state_in_s1[314], state_in_s0[314]}), .b ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, rd_I_n1795}), .c ({new_AGEMA_signal_4440, new_AGEMA_signal_4439, rd_I_n2323}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U33 ( .a ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, rd_I_n1585}), .b ({new_AGEMA_signal_3390, new_AGEMA_signal_3389, rd_I_n1689}), .c ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, rd_I_n1795}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U32 ( .a ({state_in_s2[140], state_in_s1[140], state_in_s0[140]}), .b ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, rd_I_n1324}), .c ({new_AGEMA_signal_3390, new_AGEMA_signal_3389, rd_I_n1689}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U31 ( .a ({state_in_s2[12], state_in_s1[12], state_in_s0[12]}), .b ({state_in_s2[268], state_in_s1[268], state_in_s0[268]}), .c ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, rd_I_n1324}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U30 ( .a ({new_AGEMA_signal_2874, new_AGEMA_signal_2873, rd_I_n1323}), .b ({state_in_s2[149], state_in_s1[149], state_in_s0[149]}), .c ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, rd_I_n1585}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U29 ( .a ({state_in_s2[21], state_in_s1[21], state_in_s0[21]}), .b ({state_in_s2[277], state_in_s1[277], state_in_s0[277]}), .c ({new_AGEMA_signal_2874, new_AGEMA_signal_2873, rd_I_n1323}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U28 ( .a ({state_in_s2[37], state_in_s1[37], state_in_s0[37]}), .b ({new_AGEMA_signal_3676, new_AGEMA_signal_3675, rd_I_n1650}), .c ({new_AGEMA_signal_4442, new_AGEMA_signal_4441, rd_I_n2326}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U27 ( .a ({new_AGEMA_signal_3402, new_AGEMA_signal_3401, rd_I_n1578}), .b ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, rd_I_n1629}), .c ({new_AGEMA_signal_3676, new_AGEMA_signal_3675, rd_I_n1650}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U26 ( .a ({new_AGEMA_signal_2880, new_AGEMA_signal_2879, rd_I_n1322}), .b ({state_in_s2[279], state_in_s1[279], state_in_s0[279]}), .c ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, rd_I_n1629}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U25 ( .a ({state_in_s2[23], state_in_s1[23], state_in_s0[23]}), .b ({state_in_s2[151], state_in_s1[151], state_in_s0[151]}), .c ({new_AGEMA_signal_2880, new_AGEMA_signal_2879, rd_I_n1322}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U24 ( .a ({new_AGEMA_signal_2886, new_AGEMA_signal_2885, rd_I_n1321}), .b ({state_in_s2[128], state_in_s1[128], state_in_s0[128]}), .c ({new_AGEMA_signal_3402, new_AGEMA_signal_3401, rd_I_n1578}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U23 ( .a ({state_in_s2[256], state_in_s1[256], state_in_s0[256]}), .b ({state_in_s2[0], state_in_s1[0], state_in_s0[0]}), .c ({new_AGEMA_signal_2886, new_AGEMA_signal_2885, rd_I_n1321}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U22 ( .a ({state_in_s2[133], state_in_s1[133], state_in_s0[133]}), .b ({new_AGEMA_signal_3682, new_AGEMA_signal_3681, rd_I_n1327}), .c ({new_AGEMA_signal_4444, new_AGEMA_signal_4443, rd_I_n2324}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U19 ( .a ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, rd_I_n1319}), .b ({new_AGEMA_signal_3678, new_AGEMA_signal_3677, rd_I_n1649}), .c ({new_AGEMA_signal_4446, new_AGEMA_signal_4445, rd_I_n1657}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U18 ( .a ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, rd_I_n1341}), .b ({new_AGEMA_signal_3406, new_AGEMA_signal_3405, rd_I_n1387}), .c ({new_AGEMA_signal_3678, new_AGEMA_signal_3677, rd_I_n1649}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U17 ( .a ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, rd_I_n1318}), .b ({state_in_s2[98], state_in_s1[98], state_in_s0[98]}), .c ({new_AGEMA_signal_3406, new_AGEMA_signal_3405, rd_I_n1387}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U16 ( .a ({state_in_s2[226], state_in_s1[226], state_in_s0[226]}), .b ({state_in_s2[354], state_in_s1[354], state_in_s0[354]}), .c ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, rd_I_n1318}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U15 ( .a ({new_AGEMA_signal_2898, new_AGEMA_signal_2897, rd_I_n1317}), .b ({state_in_s2[107], state_in_s1[107], state_in_s0[107]}), .c ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, rd_I_n1341}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U14 ( .a ({state_in_s2[235], state_in_s1[235], state_in_s0[235]}), .b ({state_in_s2[363], state_in_s1[363], state_in_s0[363]}), .c ({new_AGEMA_signal_2898, new_AGEMA_signal_2897, rd_I_n1317}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U13 ( .a ({state_in_s2[16], state_in_s1[16], state_in_s0[16]}), .b ({1'b0, 1'b0, rc[16]}), .c ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, rd_I_n1319}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U12 ( .a ({state_in_s2[240], state_in_s1[240], state_in_s0[240]}), .b ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, rd_I_n1460}), .c ({new_AGEMA_signal_4448, new_AGEMA_signal_4447, rd_I_n1655}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U11 ( .a ({new_AGEMA_signal_3418, new_AGEMA_signal_3417, rd_I_n1338}), .b ({new_AGEMA_signal_3414, new_AGEMA_signal_3413, rd_I_n1612}), .c ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, rd_I_n1460}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U10 ( .a ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, rd_I_n1316}), .b ({state_in_s2[66], state_in_s1[66], state_in_s0[66]}), .c ({new_AGEMA_signal_3414, new_AGEMA_signal_3413, rd_I_n1612}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U9 ( .a ({state_in_s2[194], state_in_s1[194], state_in_s0[194]}), .b ({state_in_s2[322], state_in_s1[322], state_in_s0[322]}), .c ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, rd_I_n1316}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U8 ( .a ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, rd_I_n1315}), .b ({state_in_s2[75], state_in_s1[75], state_in_s0[75]}), .c ({new_AGEMA_signal_3418, new_AGEMA_signal_3417, rd_I_n1338}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U7 ( .a ({state_in_s2[203], state_in_s1[203], state_in_s0[203]}), .b ({state_in_s2[331], state_in_s1[331], state_in_s0[331]}), .c ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, rd_I_n1315}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U6 ( .a ({state_in_s2[261], state_in_s1[261], state_in_s0[261]}), .b ({new_AGEMA_signal_3682, new_AGEMA_signal_3681, rd_I_n1327}), .c ({new_AGEMA_signal_4450, new_AGEMA_signal_4449, rd_I_n1654}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U5 ( .a ({new_AGEMA_signal_3426, new_AGEMA_signal_3425, rd_I_n1344}), .b ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, rd_I_n1635}), .c ({new_AGEMA_signal_3682, new_AGEMA_signal_3681, rd_I_n1327}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U4 ( .a ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, rd_I_n1314}), .b ({state_in_s2[375], state_in_s1[375], state_in_s0[375]}), .c ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, rd_I_n1635}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U3 ( .a ({state_in_s2[247], state_in_s1[247], state_in_s0[247]}), .b ({state_in_s2[119], state_in_s1[119], state_in_s0[119]}), .c ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, rd_I_n1314}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U2 ( .a ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, rd_I_n1313}), .b ({state_in_s2[224], state_in_s1[224], state_in_s0[224]}), .c ({new_AGEMA_signal_3426, new_AGEMA_signal_3425, rd_I_n1344}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1 ( .a ({state_in_s2[96], state_in_s1[96], state_in_s0[96]}), .b ({state_in_s2[352], state_in_s1[352], state_in_s0[352]}), .c ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, rd_I_n1313}) ) ;
    //ClockGatingController #(2) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1696 ( .a ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, rd_I_n2624}), .b ({new_AGEMA_signal_4452, new_AGEMA_signal_4451, rd_I_n2623}), .c ({state_out_s2[31], state_out_s1[31], state_out_s0[31]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1695 ( .a ({new_AGEMA_signal_3876, new_AGEMA_signal_3875, rd_I_n2622}), .b ({new_AGEMA_signal_3880, new_AGEMA_signal_3879, rd_I_n2621}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_4452, new_AGEMA_signal_4451, rd_I_n2623}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1694 ( .a ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, rd_I_n2620}), .b ({new_AGEMA_signal_4454, new_AGEMA_signal_4453, rd_I_n2619}), .c ({state_out_s2[8], state_out_s1[8], state_out_s0[8]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1693 ( .a ({new_AGEMA_signal_4288, new_AGEMA_signal_4287, rd_I_n2618}), .b ({new_AGEMA_signal_4284, new_AGEMA_signal_4283, rd_I_n2617}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_4454, new_AGEMA_signal_4453, rd_I_n2619}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1692 ( .a ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, rd_I_n2616}), .b ({new_AGEMA_signal_4456, new_AGEMA_signal_4455, rd_I_n2615}), .c ({state_out_s2[169], state_out_s1[169], state_out_s0[169]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1691 ( .a ({new_AGEMA_signal_3688, new_AGEMA_signal_3687, rd_I_n2614}), .b ({new_AGEMA_signal_3684, new_AGEMA_signal_3683, rd_I_n2613}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_4456, new_AGEMA_signal_4455, rd_I_n2615}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1690 ( .a ({new_AGEMA_signal_3746, new_AGEMA_signal_3745, rd_I_n2612}), .b ({new_AGEMA_signal_4458, new_AGEMA_signal_4457, rd_I_n2611}), .c ({state_out_s2[160], state_out_s1[160], state_out_s0[160]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1689 ( .a ({new_AGEMA_signal_3748, new_AGEMA_signal_3747, rd_I_n2610}), .b ({new_AGEMA_signal_3744, new_AGEMA_signal_3743, rd_I_n2609}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_4458, new_AGEMA_signal_4457, rd_I_n2611}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1688 ( .a ({new_AGEMA_signal_3758, new_AGEMA_signal_3757, rd_I_n2608}), .b ({new_AGEMA_signal_4460, new_AGEMA_signal_4459, rd_I_n2607}), .c ({state_out_s2[347], state_out_s1[347], state_out_s0[347]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1687 ( .a ({new_AGEMA_signal_3760, new_AGEMA_signal_3759, rd_I_n2606}), .b ({new_AGEMA_signal_3756, new_AGEMA_signal_3755, rd_I_n2605}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_4460, new_AGEMA_signal_4459, rd_I_n2607}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1686 ( .a ({new_AGEMA_signal_5216, new_AGEMA_signal_5215, rd_I_n2604}), .b ({new_AGEMA_signal_4116, new_AGEMA_signal_4115, rd_I_n2603}), .c ({state_out_s2[338], state_out_s1[338], state_out_s0[338]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1685 ( .a ({new_AGEMA_signal_4462, new_AGEMA_signal_4461, rd_I_n2602}), .b ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, rd_I_n2601}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_5216, new_AGEMA_signal_5215, rd_I_n2604}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1683 ( .a ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, rd_I_n2599}), .b ({new_AGEMA_signal_4464, new_AGEMA_signal_4463, rd_I_n2598}), .c ({state_out_s2[22], state_out_s1[22], state_out_s0[22]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1682 ( .a ({new_AGEMA_signal_3874, new_AGEMA_signal_3873, rd_I_n2597}), .b ({new_AGEMA_signal_3870, new_AGEMA_signal_3869, rd_I_n2596}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_4464, new_AGEMA_signal_4463, rd_I_n2598}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1681 ( .a ({new_AGEMA_signal_3740, new_AGEMA_signal_3739, rd_I_n2595}), .b ({new_AGEMA_signal_4466, new_AGEMA_signal_4465, rd_I_n2594}), .c ({state_out_s2[183], state_out_s1[183], state_out_s0[183]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1680 ( .a ({new_AGEMA_signal_3742, new_AGEMA_signal_3741, rd_I_n2593}), .b ({new_AGEMA_signal_3738, new_AGEMA_signal_3737, rd_I_n2592}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_4466, new_AGEMA_signal_4465, rd_I_n2594}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1679 ( .a ({new_AGEMA_signal_5222, new_AGEMA_signal_5221, rd_I_n2591}), .b ({new_AGEMA_signal_3694, new_AGEMA_signal_3693, rd_I_n2590}), .c ({state_out_s2[329], state_out_s1[329], state_out_s0[329]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1678 ( .a ({new_AGEMA_signal_4468, new_AGEMA_signal_4467, rd_I_n2589}), .b ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, rd_I_n2588}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_5222, new_AGEMA_signal_5221, rd_I_n2591}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1676 ( .a ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, rd_I_n2586}), .b ({new_AGEMA_signal_4470, new_AGEMA_signal_4469, rd_I_n2585}), .c ({state_out_s2[20], state_out_s1[20], state_out_s0[20]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1675 ( .a ({new_AGEMA_signal_4054, new_AGEMA_signal_4053, rd_I_n2584}), .b ({new_AGEMA_signal_4050, new_AGEMA_signal_4049, rd_I_n2583}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_4470, new_AGEMA_signal_4469, rd_I_n2585}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1674 ( .a ({new_AGEMA_signal_5042, new_AGEMA_signal_5041, rd_I_n2582}), .b ({new_AGEMA_signal_4472, new_AGEMA_signal_4471, rd_I_n2581}), .c ({state_out_s2[11], state_out_s1[11], state_out_s0[11]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1673 ( .a ({new_AGEMA_signal_4056, new_AGEMA_signal_4055, rd_I_n2580}), .b ({new_AGEMA_signal_4060, new_AGEMA_signal_4059, rd_I_n2579}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_4472, new_AGEMA_signal_4471, rd_I_n2581}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1672 ( .a ({new_AGEMA_signal_5228, new_AGEMA_signal_5227, rd_I_n2578}), .b ({new_AGEMA_signal_3726, new_AGEMA_signal_3725, rd_I_n2577}), .c ({state_out_s2[181], state_out_s1[181], state_out_s0[181]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1671 ( .a ({new_AGEMA_signal_4474, new_AGEMA_signal_4473, rd_I_n2576}), .b ({new_AGEMA_signal_3728, new_AGEMA_signal_3727, rd_I_n2575}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_5228, new_AGEMA_signal_5227, rd_I_n2578}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1669 ( .a ({new_AGEMA_signal_5230, new_AGEMA_signal_5229, rd_I_n2573}), .b ({new_AGEMA_signal_3732, new_AGEMA_signal_3731, rd_I_n2572}), .c ({state_out_s2[172], state_out_s1[172], state_out_s0[172]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1668 ( .a ({new_AGEMA_signal_4476, new_AGEMA_signal_4475, rd_I_n2571}), .b ({new_AGEMA_signal_3734, new_AGEMA_signal_3733, rd_I_n2570}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_5230, new_AGEMA_signal_5229, rd_I_n2573}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1666 ( .a ({new_AGEMA_signal_5232, new_AGEMA_signal_5231, rd_I_n2568}), .b ({new_AGEMA_signal_3870, new_AGEMA_signal_3869, rd_I_n2596}), .c ({state_out_s2[350], state_out_s1[350], state_out_s0[350]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1665 ( .a ({new_AGEMA_signal_4478, new_AGEMA_signal_4477, rd_I_n2567}), .b ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, rd_I_n2599}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_5232, new_AGEMA_signal_5231, rd_I_n2568}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1663 ( .a ({new_AGEMA_signal_5234, new_AGEMA_signal_5233, rd_I_n2566}), .b ({new_AGEMA_signal_3880, new_AGEMA_signal_3879, rd_I_n2621}), .c ({state_out_s2[327], state_out_s1[327], state_out_s0[327]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1662 ( .a ({new_AGEMA_signal_4480, new_AGEMA_signal_4479, rd_I_n2565}), .b ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, rd_I_n2624}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_5234, new_AGEMA_signal_5233, rd_I_n2566}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1660 ( .a ({new_AGEMA_signal_3890, new_AGEMA_signal_3889, rd_I_n2564}), .b ({new_AGEMA_signal_4482, new_AGEMA_signal_4481, rd_I_n2563}), .c ({state_out_s2[126], state_out_s1[126], state_out_s0[126]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1659 ( .a ({new_AGEMA_signal_3892, new_AGEMA_signal_3891, rd_I_n2562}), .b ({new_AGEMA_signal_3888, new_AGEMA_signal_3887, rd_I_n2561}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_4482, new_AGEMA_signal_4481, rd_I_n2563}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1658 ( .a ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, rd_I_n2560}), .b ({new_AGEMA_signal_4126, new_AGEMA_signal_4125, rd_I_n2559}), .c ({state_out_s2[117], state_out_s1[117], state_out_s0[117]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1657 ( .a ({new_AGEMA_signal_4484, new_AGEMA_signal_4483, rd_I_n2558}), .b ({new_AGEMA_signal_4124, new_AGEMA_signal_4123, rd_I_n2557}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, rd_I_n2560}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1655 ( .a ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, rd_I_n2555}), .b ({new_AGEMA_signal_4236, new_AGEMA_signal_4235, rd_I_n2554}), .c ({state_out_s2[159], state_out_s1[159], state_out_s0[159]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1654 ( .a ({new_AGEMA_signal_5240, new_AGEMA_signal_5239, rd_I_n2553}), .b ({new_AGEMA_signal_4238, new_AGEMA_signal_4237, rd_I_n2552}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, rd_I_n2555}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1652 ( .a ({new_AGEMA_signal_5242, new_AGEMA_signal_5241, rd_I_n2550}), .b ({new_AGEMA_signal_3852, new_AGEMA_signal_3851, rd_I_n2549}), .c ({state_out_s2[150], state_out_s1[150], state_out_s0[150]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1651 ( .a ({new_AGEMA_signal_4486, new_AGEMA_signal_4485, rd_I_n2548}), .b ({new_AGEMA_signal_3854, new_AGEMA_signal_3853, rd_I_n2547}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_5242, new_AGEMA_signal_5241, rd_I_n2550}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1649 ( .a ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, rd_I_n2545}), .b ({new_AGEMA_signal_4224, new_AGEMA_signal_4223, rd_I_n2544}), .c ({state_out_s2[305], state_out_s1[305], state_out_s0[305]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1648 ( .a ({new_AGEMA_signal_4488, new_AGEMA_signal_4487, rd_I_n2543}), .b ({new_AGEMA_signal_4226, new_AGEMA_signal_4225, rd_I_n2542}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, rd_I_n2545}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1646 ( .a ({new_AGEMA_signal_3800, new_AGEMA_signal_3799, rd_I_n2540}), .b ({new_AGEMA_signal_4490, new_AGEMA_signal_4489, rd_I_n2539}), .c ({state_out_s2[296], state_out_s1[296], state_out_s0[296]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1645 ( .a ({new_AGEMA_signal_3802, new_AGEMA_signal_3801, rd_I_n2538}), .b ({new_AGEMA_signal_3798, new_AGEMA_signal_3797, rd_I_n2537}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_4490, new_AGEMA_signal_4489, rd_I_n2539}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1644 ( .a ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, rd_I_n2601}), .b ({new_AGEMA_signal_4492, new_AGEMA_signal_4491, rd_I_n2536}), .c ({state_out_s2[10], state_out_s1[10], state_out_s0[10]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1643 ( .a ({new_AGEMA_signal_4120, new_AGEMA_signal_4119, rd_I_n2600}), .b ({new_AGEMA_signal_4116, new_AGEMA_signal_4115, rd_I_n2603}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_4492, new_AGEMA_signal_4491, rd_I_n2536}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1642 ( .a ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, rd_I_n2588}), .b ({new_AGEMA_signal_4494, new_AGEMA_signal_4493, rd_I_n2535}), .c ({state_out_s2[1], state_out_s1[1], state_out_s0[1]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1641 ( .a ({new_AGEMA_signal_3690, new_AGEMA_signal_3689, rd_I_n2587}), .b ({new_AGEMA_signal_3694, new_AGEMA_signal_3693, rd_I_n2590}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_4494, new_AGEMA_signal_4493, rd_I_n2535}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1640 ( .a ({new_AGEMA_signal_5252, new_AGEMA_signal_5251, rd_I_n2534}), .b ({new_AGEMA_signal_3774, new_AGEMA_signal_3773, rd_I_n2533}), .c ({state_out_s2[171], state_out_s1[171], state_out_s0[171]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1639 ( .a ({new_AGEMA_signal_4496, new_AGEMA_signal_4495, rd_I_n2532}), .b ({new_AGEMA_signal_3776, new_AGEMA_signal_3775, rd_I_n2531}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_5252, new_AGEMA_signal_5251, rd_I_n2534}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1637 ( .a ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, rd_I_n2529}), .b ({new_AGEMA_signal_4498, new_AGEMA_signal_4497, rd_I_n2528}), .c ({state_out_s2[162], state_out_s1[162], state_out_s0[162]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1636 ( .a ({new_AGEMA_signal_3718, new_AGEMA_signal_3717, rd_I_n2527}), .b ({new_AGEMA_signal_3714, new_AGEMA_signal_3713, rd_I_n2526}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_4498, new_AGEMA_signal_4497, rd_I_n2528}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1635 ( .a ({new_AGEMA_signal_3854, new_AGEMA_signal_3853, rd_I_n2547}), .b ({new_AGEMA_signal_4500, new_AGEMA_signal_4499, rd_I_n2525}), .c ({state_out_s2[349], state_out_s1[349], state_out_s0[349]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1634 ( .a ({new_AGEMA_signal_3856, new_AGEMA_signal_3855, rd_I_n2546}), .b ({new_AGEMA_signal_3852, new_AGEMA_signal_3851, rd_I_n2549}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_4500, new_AGEMA_signal_4499, rd_I_n2525}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1633 ( .a ({new_AGEMA_signal_5258, new_AGEMA_signal_5257, rd_I_n2524}), .b ({new_AGEMA_signal_3946, new_AGEMA_signal_3945, rd_I_n2523}), .c ({state_out_s2[340], state_out_s1[340], state_out_s0[340]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1632 ( .a ({new_AGEMA_signal_4502, new_AGEMA_signal_4501, rd_I_n2522}), .b ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, rd_I_n2521}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_5258, new_AGEMA_signal_5257, rd_I_n2524}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1630 ( .a ({new_AGEMA_signal_5260, new_AGEMA_signal_5259, rd_I_n2519}), .b ({new_AGEMA_signal_4856, new_AGEMA_signal_4855, rd_I_n2518}), .c ({state_out_s2[23], state_out_s1[23], state_out_s0[23]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1629 ( .a ({new_AGEMA_signal_4504, new_AGEMA_signal_4503, rd_I_n2517}), .b ({new_AGEMA_signal_3836, new_AGEMA_signal_3835, rd_I_n2516}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_5260, new_AGEMA_signal_5259, rd_I_n2519}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1627 ( .a ({new_AGEMA_signal_5262, new_AGEMA_signal_5261, rd_I_n2514}), .b ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, rd_I_n2513}), .c ({state_out_s2[14], state_out_s1[14], state_out_s0[14]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1626 ( .a ({new_AGEMA_signal_4506, new_AGEMA_signal_4505, rd_I_n2512}), .b ({new_AGEMA_signal_3842, new_AGEMA_signal_3841, rd_I_n2511}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_5262, new_AGEMA_signal_5261, rd_I_n2514}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1624 ( .a ({new_AGEMA_signal_5264, new_AGEMA_signal_5263, rd_I_n2509}), .b ({new_AGEMA_signal_3972, new_AGEMA_signal_3971, rd_I_n2508}), .c ({state_out_s2[184], state_out_s1[184], state_out_s0[184]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1623 ( .a ({new_AGEMA_signal_4508, new_AGEMA_signal_4507, rd_I_n2507}), .b ({new_AGEMA_signal_3974, new_AGEMA_signal_3973, rd_I_n2506}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_5264, new_AGEMA_signal_5263, rd_I_n2509}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1621 ( .a ({new_AGEMA_signal_5266, new_AGEMA_signal_5265, rd_I_n2504}), .b ({new_AGEMA_signal_3966, new_AGEMA_signal_3965, rd_I_n2503}), .c ({state_out_s2[175], state_out_s1[175], state_out_s0[175]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1620 ( .a ({new_AGEMA_signal_4510, new_AGEMA_signal_4509, rd_I_n2502}), .b ({new_AGEMA_signal_3968, new_AGEMA_signal_3967, rd_I_n2501}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_5266, new_AGEMA_signal_5265, rd_I_n2504}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1618 ( .a ({new_AGEMA_signal_5268, new_AGEMA_signal_5267, rd_I_n2499}), .b ({new_AGEMA_signal_4404, new_AGEMA_signal_4403, rd_I_n2498}), .c ({state_out_s2[330], state_out_s1[330], state_out_s0[330]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1617 ( .a ({new_AGEMA_signal_4512, new_AGEMA_signal_4511, rd_I_n2497}), .b ({new_AGEMA_signal_4406, new_AGEMA_signal_4405, rd_I_n2496}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_5268, new_AGEMA_signal_5267, rd_I_n2499}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1615 ( .a ({new_AGEMA_signal_5270, new_AGEMA_signal_5269, rd_I_n2494}), .b ({new_AGEMA_signal_4422, new_AGEMA_signal_4421, rd_I_n2493}), .c ({state_out_s2[321], state_out_s1[321], state_out_s0[321]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1614 ( .a ({new_AGEMA_signal_4514, new_AGEMA_signal_4513, rd_I_n2492}), .b ({new_AGEMA_signal_4424, new_AGEMA_signal_4423, rd_I_n2491}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_5270, new_AGEMA_signal_5269, rd_I_n2494}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1612 ( .a ({new_AGEMA_signal_3914, new_AGEMA_signal_3913, rd_I_n2489}), .b ({new_AGEMA_signal_4516, new_AGEMA_signal_4515, rd_I_n2488}), .c ({state_out_s2[41], state_out_s1[41], state_out_s0[41]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1611 ( .a ({new_AGEMA_signal_3916, new_AGEMA_signal_3915, rd_I_n2487}), .b ({new_AGEMA_signal_3912, new_AGEMA_signal_3911, rd_I_n2486}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_4516, new_AGEMA_signal_4515, rd_I_n2488}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1610 ( .a ({new_AGEMA_signal_3770, new_AGEMA_signal_3769, rd_I_n2485}), .b ({new_AGEMA_signal_4518, new_AGEMA_signal_4517, rd_I_n2484}), .c ({state_out_s2[32], state_out_s1[32], state_out_s0[32]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1609 ( .a ({new_AGEMA_signal_3772, new_AGEMA_signal_3771, rd_I_n2483}), .b ({new_AGEMA_signal_3768, new_AGEMA_signal_3767, rd_I_n2482}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_4518, new_AGEMA_signal_4517, rd_I_n2484}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1608 ( .a ({new_AGEMA_signal_5276, new_AGEMA_signal_5275, rd_I_n2481}), .b ({new_AGEMA_signal_4220, new_AGEMA_signal_4219, rd_I_n2480}), .c ({state_out_s2[202], state_out_s1[202], state_out_s0[202]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1607 ( .a ({new_AGEMA_signal_4520, new_AGEMA_signal_4519, rd_I_n2479}), .b ({new_AGEMA_signal_4222, new_AGEMA_signal_4221, rd_I_n2478}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_5276, new_AGEMA_signal_5275, rd_I_n2481}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1605 ( .a ({new_AGEMA_signal_3896, new_AGEMA_signal_3895, rd_I_n2476}), .b ({new_AGEMA_signal_4522, new_AGEMA_signal_4521, rd_I_n2475}), .c ({state_out_s2[193], state_out_s1[193], state_out_s0[193]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1604 ( .a ({new_AGEMA_signal_3894, new_AGEMA_signal_3893, rd_I_n2474}), .b ({new_AGEMA_signal_3898, new_AGEMA_signal_3897, rd_I_n2473}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_4522, new_AGEMA_signal_4521, rd_I_n2475}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1603 ( .a ({new_AGEMA_signal_3728, new_AGEMA_signal_3727, rd_I_n2575}), .b ({new_AGEMA_signal_4524, new_AGEMA_signal_4523, rd_I_n2472}), .c ({state_out_s2[380], state_out_s1[380], state_out_s0[380]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1602 ( .a ({new_AGEMA_signal_3730, new_AGEMA_signal_3729, rd_I_n2574}), .b ({new_AGEMA_signal_3726, new_AGEMA_signal_3725, rd_I_n2577}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_4524, new_AGEMA_signal_4523, rd_I_n2472}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1601 ( .a ({new_AGEMA_signal_3734, new_AGEMA_signal_3733, rd_I_n2570}), .b ({new_AGEMA_signal_4526, new_AGEMA_signal_4525, rd_I_n2471}), .c ({state_out_s2[371], state_out_s1[371], state_out_s0[371]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1600 ( .a ({new_AGEMA_signal_3736, new_AGEMA_signal_3735, rd_I_n2569}), .b ({new_AGEMA_signal_3732, new_AGEMA_signal_3731, rd_I_n2572}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_4526, new_AGEMA_signal_4525, rd_I_n2471}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1599 ( .a ({new_AGEMA_signal_5284, new_AGEMA_signal_5283, rd_I_n2470}), .b ({new_AGEMA_signal_3702, new_AGEMA_signal_3701, rd_I_n2469}), .c ({state_out_s2[91], state_out_s1[91], state_out_s0[91]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1598 ( .a ({new_AGEMA_signal_4528, new_AGEMA_signal_4527, rd_I_n2468}), .b ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, rd_I_n2467}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_5284, new_AGEMA_signal_5283, rd_I_n2470}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1596 ( .a ({new_AGEMA_signal_5286, new_AGEMA_signal_5285, rd_I_n2465}), .b ({new_AGEMA_signal_3696, new_AGEMA_signal_3695, rd_I_n2464}), .c ({state_out_s2[68], state_out_s1[68], state_out_s0[68]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1595 ( .a ({new_AGEMA_signal_4530, new_AGEMA_signal_4529, rd_I_n2463}), .b ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, rd_I_n2462}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_5286, new_AGEMA_signal_5285, rd_I_n2465}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1593 ( .a ({new_AGEMA_signal_4310, new_AGEMA_signal_4309, rd_I_n2460}), .b ({new_AGEMA_signal_4532, new_AGEMA_signal_4531, rd_I_n2459}), .c ({state_out_s2[252], state_out_s1[252], state_out_s0[252]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1592 ( .a ({new_AGEMA_signal_4308, new_AGEMA_signal_4307, rd_I_n2458}), .b ({new_AGEMA_signal_4312, new_AGEMA_signal_4311, rd_I_n2457}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_4532, new_AGEMA_signal_4531, rd_I_n2459}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1591 ( .a ({new_AGEMA_signal_4432, new_AGEMA_signal_4431, rd_I_n2456}), .b ({new_AGEMA_signal_4534, new_AGEMA_signal_4533, rd_I_n2455}), .c ({state_out_s2[229], state_out_s1[229], state_out_s0[229]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1590 ( .a ({new_AGEMA_signal_4428, new_AGEMA_signal_4427, rd_I_n2454}), .b ({new_AGEMA_signal_4430, new_AGEMA_signal_4429, rd_I_n2453}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_4534, new_AGEMA_signal_4533, rd_I_n2455}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1589 ( .a ({new_AGEMA_signal_3956, new_AGEMA_signal_3955, rd_I_n2452}), .b ({new_AGEMA_signal_4536, new_AGEMA_signal_4535, rd_I_n2451}), .c ({state_out_s2[279], state_out_s1[279], state_out_s0[279]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1588 ( .a ({new_AGEMA_signal_3958, new_AGEMA_signal_3957, rd_I_n2450}), .b ({new_AGEMA_signal_3954, new_AGEMA_signal_3953, rd_I_n2449}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_4536, new_AGEMA_signal_4535, rd_I_n2451}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1587 ( .a ({new_AGEMA_signal_3752, new_AGEMA_signal_3751, rd_I_n2448}), .b ({new_AGEMA_signal_4538, new_AGEMA_signal_4537, rd_I_n2447}), .c ({state_out_s2[270], state_out_s1[270], state_out_s0[270]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1586 ( .a ({new_AGEMA_signal_3754, new_AGEMA_signal_3753, rd_I_n2446}), .b ({new_AGEMA_signal_3750, new_AGEMA_signal_3749, rd_I_n2445}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_4538, new_AGEMA_signal_4537, rd_I_n2447}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1585 ( .a ({new_AGEMA_signal_5296, new_AGEMA_signal_5295, rd_I_n2444}), .b ({new_AGEMA_signal_3744, new_AGEMA_signal_3743, rd_I_n2609}), .c ({state_out_s2[63], state_out_s1[63], state_out_s0[63]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1584 ( .a ({new_AGEMA_signal_4540, new_AGEMA_signal_4539, rd_I_n2443}), .b ({new_AGEMA_signal_3746, new_AGEMA_signal_3745, rd_I_n2612}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_5296, new_AGEMA_signal_5295, rd_I_n2444}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1582 ( .a ({new_AGEMA_signal_5298, new_AGEMA_signal_5297, rd_I_n2442}), .b ({new_AGEMA_signal_3684, new_AGEMA_signal_3683, rd_I_n2613}), .c ({state_out_s2[40], state_out_s1[40], state_out_s0[40]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1581 ( .a ({new_AGEMA_signal_4542, new_AGEMA_signal_4541, rd_I_n2441}), .b ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, rd_I_n2616}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_5298, new_AGEMA_signal_5297, rd_I_n2442}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1579 ( .a ({new_AGEMA_signal_5300, new_AGEMA_signal_5299, rd_I_n2440}), .b ({new_AGEMA_signal_4018, new_AGEMA_signal_4017, rd_I_n2439}), .c ({state_out_s2[201], state_out_s1[201], state_out_s0[201]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1578 ( .a ({new_AGEMA_signal_4544, new_AGEMA_signal_4543, rd_I_n2438}), .b ({new_AGEMA_signal_4016, new_AGEMA_signal_4015, rd_I_n2437}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_5300, new_AGEMA_signal_5299, rd_I_n2440}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1576 ( .a ({new_AGEMA_signal_3926, new_AGEMA_signal_3925, rd_I_n2435}), .b ({new_AGEMA_signal_4546, new_AGEMA_signal_4545, rd_I_n2434}), .c ({state_out_s2[192], state_out_s1[192], state_out_s0[192]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1575 ( .a ({new_AGEMA_signal_3924, new_AGEMA_signal_3923, rd_I_n2433}), .b ({new_AGEMA_signal_3928, new_AGEMA_signal_3927, rd_I_n2432}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_4546, new_AGEMA_signal_4545, rd_I_n2434}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1574 ( .a ({new_AGEMA_signal_3764, new_AGEMA_signal_3763, rd_I_n2431}), .b ({new_AGEMA_signal_4548, new_AGEMA_signal_4547, rd_I_n2430}), .c ({state_out_s2[379], state_out_s1[379], state_out_s0[379]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1573 ( .a ({new_AGEMA_signal_3766, new_AGEMA_signal_3765, rd_I_n2429}), .b ({new_AGEMA_signal_3762, new_AGEMA_signal_3761, rd_I_n2428}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_4548, new_AGEMA_signal_4547, rd_I_n2430}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1572 ( .a ({new_AGEMA_signal_3776, new_AGEMA_signal_3775, rd_I_n2531}), .b ({new_AGEMA_signal_4550, new_AGEMA_signal_4549, rd_I_n2427}), .c ({state_out_s2[370], state_out_s1[370], state_out_s0[370]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1571 ( .a ({new_AGEMA_signal_3778, new_AGEMA_signal_3777, rd_I_n2530}), .b ({new_AGEMA_signal_3774, new_AGEMA_signal_3773, rd_I_n2533}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_4550, new_AGEMA_signal_4549, rd_I_n2427}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1570 ( .a ({new_AGEMA_signal_4244, new_AGEMA_signal_4243, rd_I_n2426}), .b ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, rd_I_n2425}), .c ({state_out_s2[62], state_out_s1[62], state_out_s0[62]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1569 ( .a ({new_AGEMA_signal_4242, new_AGEMA_signal_4241, rd_I_n2424}), .b ({new_AGEMA_signal_4246, new_AGEMA_signal_4245, rd_I_n2423}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_4552, new_AGEMA_signal_4551, rd_I_n2425}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1568 ( .a ({new_AGEMA_signal_4112, new_AGEMA_signal_4111, rd_I_n2422}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, rd_I_n2421}), .c ({state_out_s2[39], state_out_s1[39], state_out_s0[39]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1567 ( .a ({new_AGEMA_signal_4110, new_AGEMA_signal_4109, rd_I_n2420}), .b ({new_AGEMA_signal_4114, new_AGEMA_signal_4113, rd_I_n2419}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, rd_I_n2421}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1566 ( .a ({new_AGEMA_signal_3962, new_AGEMA_signal_3961, rd_I_n2418}), .b ({new_AGEMA_signal_4556, new_AGEMA_signal_4555, rd_I_n2417}), .c ({state_out_s2[223], state_out_s1[223], state_out_s0[223]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1565 ( .a ({new_AGEMA_signal_3964, new_AGEMA_signal_3963, rd_I_n2416}), .b ({new_AGEMA_signal_3960, new_AGEMA_signal_3959, rd_I_n2415}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_4556, new_AGEMA_signal_4555, rd_I_n2417}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1564 ( .a ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, rd_I_n2414}), .b ({new_AGEMA_signal_4128, new_AGEMA_signal_4127, rd_I_n2413}), .c ({state_out_s2[200], state_out_s1[200], state_out_s0[200]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1563 ( .a ({new_AGEMA_signal_4558, new_AGEMA_signal_4557, rd_I_n2412}), .b ({new_AGEMA_signal_4130, new_AGEMA_signal_4129, rd_I_n2411}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_5314, new_AGEMA_signal_5313, rd_I_n2414}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1561 ( .a ({new_AGEMA_signal_5316, new_AGEMA_signal_5315, rd_I_n2409}), .b ({new_AGEMA_signal_4386, new_AGEMA_signal_4385, rd_I_n2408}), .c ({state_out_s2[378], state_out_s1[378], state_out_s0[378]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1560 ( .a ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, rd_I_n2407}), .b ({new_AGEMA_signal_4388, new_AGEMA_signal_4387, rd_I_n2406}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_5316, new_AGEMA_signal_5315, rd_I_n2409}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1558 ( .a ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, rd_I_n2404}), .b ({new_AGEMA_signal_3912, new_AGEMA_signal_3911, rd_I_n2486}), .c ({state_out_s2[369], state_out_s1[369], state_out_s0[369]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1557 ( .a ({new_AGEMA_signal_4562, new_AGEMA_signal_4561, rd_I_n2403}), .b ({new_AGEMA_signal_3914, new_AGEMA_signal_3913, rd_I_n2489}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_5318, new_AGEMA_signal_5317, rd_I_n2404}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1555 ( .a ({new_AGEMA_signal_4136, new_AGEMA_signal_4135, rd_I_n2402}), .b ({new_AGEMA_signal_4564, new_AGEMA_signal_4563, rd_I_n2401}), .c ({state_out_s2[103], state_out_s1[103], state_out_s0[103]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1554 ( .a ({new_AGEMA_signal_4134, new_AGEMA_signal_4133, rd_I_n2400}), .b ({new_AGEMA_signal_4138, new_AGEMA_signal_4137, rd_I_n2399}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_4564, new_AGEMA_signal_4563, rd_I_n2401}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1553 ( .a ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, rd_I_n2398}), .b ({new_AGEMA_signal_4104, new_AGEMA_signal_4103, rd_I_n2397}), .c ({state_out_s2[136], state_out_s1[136], state_out_s0[136]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1552 ( .a ({new_AGEMA_signal_4566, new_AGEMA_signal_4565, rd_I_n2396}), .b ({new_AGEMA_signal_4106, new_AGEMA_signal_4105, rd_I_n2395}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, rd_I_n2398}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1550 ( .a ({new_AGEMA_signal_5324, new_AGEMA_signal_5323, rd_I_n2393}), .b ({new_AGEMA_signal_3984, new_AGEMA_signal_3983, rd_I_n2392}), .c ({state_out_s2[314], state_out_s1[314], state_out_s0[314]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1549 ( .a ({new_AGEMA_signal_4568, new_AGEMA_signal_4567, rd_I_n2391}), .b ({new_AGEMA_signal_3986, new_AGEMA_signal_3985, rd_I_n2390}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_5324, new_AGEMA_signal_5323, rd_I_n2393}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1547 ( .a ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, rd_I_n2388}), .b ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, rd_I_n2387}), .c ({state_out_s2[24], state_out_s1[24], state_out_s0[24]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1546 ( .a ({new_AGEMA_signal_4570, new_AGEMA_signal_4569, rd_I_n2386}), .b ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, rd_I_n2385}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_5326, new_AGEMA_signal_5325, rd_I_n2388}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1544 ( .a ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, rd_I_n2383}), .b ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, rd_I_n2382}), .c ({state_out_s2[185], state_out_s1[185], state_out_s0[185]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1543 ( .a ({new_AGEMA_signal_3724, new_AGEMA_signal_3723, rd_I_n2381}), .b ({new_AGEMA_signal_3720, new_AGEMA_signal_3719, rd_I_n2380}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, rd_I_n2382}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1542 ( .a ({new_AGEMA_signal_5330, new_AGEMA_signal_5329, rd_I_n2379}), .b ({new_AGEMA_signal_4350, new_AGEMA_signal_4349, rd_I_n2378}), .c ({state_out_s2[331], state_out_s1[331], state_out_s0[331]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1541 ( .a ({new_AGEMA_signal_4574, new_AGEMA_signal_4573, rd_I_n2377}), .b ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, rd_I_n2376}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_5330, new_AGEMA_signal_5329, rd_I_n2379}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1539 ( .a ({new_AGEMA_signal_3782, new_AGEMA_signal_3781, rd_I_n2374}), .b ({new_AGEMA_signal_4576, new_AGEMA_signal_4575, rd_I_n2373}), .c ({state_out_s2[61], state_out_s1[61], state_out_s0[61]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1538 ( .a ({new_AGEMA_signal_3784, new_AGEMA_signal_3783, rd_I_n2372}), .b ({new_AGEMA_signal_3780, new_AGEMA_signal_3779, rd_I_n2371}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_4576, new_AGEMA_signal_4575, rd_I_n2373}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1537 ( .a ({new_AGEMA_signal_4028, new_AGEMA_signal_4027, rd_I_n2370}), .b ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, rd_I_n2369}), .c ({state_out_s2[38], state_out_s1[38], state_out_s0[38]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1536 ( .a ({new_AGEMA_signal_4026, new_AGEMA_signal_4025, rd_I_n2368}), .b ({new_AGEMA_signal_4030, new_AGEMA_signal_4029, rd_I_n2367}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, rd_I_n2369}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1535 ( .a ({new_AGEMA_signal_3992, new_AGEMA_signal_3991, rd_I_n2366}), .b ({new_AGEMA_signal_4580, new_AGEMA_signal_4579, rd_I_n2365}), .c ({state_out_s2[222], state_out_s1[222], state_out_s0[222]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1534 ( .a ({new_AGEMA_signal_3990, new_AGEMA_signal_3989, rd_I_n2364}), .b ({new_AGEMA_signal_3994, new_AGEMA_signal_3993, rd_I_n2363}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_4580, new_AGEMA_signal_4579, rd_I_n2365}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1533 ( .a ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, rd_I_n2362}), .b ({new_AGEMA_signal_3750, new_AGEMA_signal_3749, rd_I_n2445}), .c ({state_out_s2[199], state_out_s1[199], state_out_s0[199]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1532 ( .a ({new_AGEMA_signal_4582, new_AGEMA_signal_4581, rd_I_n2361}), .b ({new_AGEMA_signal_3752, new_AGEMA_signal_3751, rd_I_n2448}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_5338, new_AGEMA_signal_5337, rd_I_n2362}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1530 ( .a ({new_AGEMA_signal_3812, new_AGEMA_signal_3811, rd_I_n2360}), .b ({new_AGEMA_signal_4584, new_AGEMA_signal_4583, rd_I_n2359}), .c ({state_out_s2[377], state_out_s1[377], state_out_s0[377]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1529 ( .a ({new_AGEMA_signal_3814, new_AGEMA_signal_3813, rd_I_n2358}), .b ({new_AGEMA_signal_3810, new_AGEMA_signal_3809, rd_I_n2357}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_4584, new_AGEMA_signal_4583, rd_I_n2359}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1528 ( .a ({new_AGEMA_signal_3688, new_AGEMA_signal_3687, rd_I_n2614}), .b ({new_AGEMA_signal_4586, new_AGEMA_signal_4585, rd_I_n2356}), .c ({state_out_s2[368], state_out_s1[368], state_out_s0[368]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1527 ( .a ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, rd_I_n2616}), .b ({new_AGEMA_signal_3684, new_AGEMA_signal_3683, rd_I_n2613}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_4586, new_AGEMA_signal_4585, rd_I_n2356}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1523 ( .a ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, rd_I_n2352}), .b ({new_AGEMA_signal_4300, new_AGEMA_signal_4299, rd_I_n2351}), .c ({state_out_s2[124], state_out_s1[124], state_out_s0[124]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1522 ( .a ({new_AGEMA_signal_4588, new_AGEMA_signal_4587, rd_I_n2350}), .b ({new_AGEMA_signal_4298, new_AGEMA_signal_4297, rd_I_n2349}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_5344, new_AGEMA_signal_5343, rd_I_n2352}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1520 ( .a ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, rd_I_n2347}), .b ({new_AGEMA_signal_4294, new_AGEMA_signal_4293, rd_I_n2346}), .c ({state_out_s2[115], state_out_s1[115], state_out_s0[115]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1519 ( .a ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, rd_I_n2345}), .b ({new_AGEMA_signal_4292, new_AGEMA_signal_4291, rd_I_n2344}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, rd_I_n2347}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1517 ( .a ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, rd_I_n2342}), .b ({new_AGEMA_signal_3804, new_AGEMA_signal_3803, rd_I_n2341}), .c ({state_out_s2[157], state_out_s1[157], state_out_s0[157]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1516 ( .a ({new_AGEMA_signal_4592, new_AGEMA_signal_4591, rd_I_n2340}), .b ({new_AGEMA_signal_3806, new_AGEMA_signal_3805, rd_I_n2339}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_5348, new_AGEMA_signal_5347, rd_I_n2342}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1514 ( .a ({new_AGEMA_signal_5350, new_AGEMA_signal_5349, rd_I_n2337}), .b ({new_AGEMA_signal_3756, new_AGEMA_signal_3755, rd_I_n2605}), .c ({state_out_s2[148], state_out_s1[148], state_out_s0[148]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1513 ( .a ({new_AGEMA_signal_4594, new_AGEMA_signal_4593, rd_I_n2336}), .b ({new_AGEMA_signal_3758, new_AGEMA_signal_3757, rd_I_n2608}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_5350, new_AGEMA_signal_5349, rd_I_n2337}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1511 ( .a ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, rd_I_n2335}), .b ({new_AGEMA_signal_4138, new_AGEMA_signal_4137, rd_I_n2399}), .c ({state_out_s2[303], state_out_s1[303], state_out_s0[303]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1510 ( .a ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, rd_I_n2334}), .b ({new_AGEMA_signal_4136, new_AGEMA_signal_4135, rd_I_n2402}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, rd_I_n2335}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1508 ( .a ({new_AGEMA_signal_5354, new_AGEMA_signal_5353, rd_I_n2333}), .b ({new_AGEMA_signal_3888, new_AGEMA_signal_3887, rd_I_n2561}), .c ({state_out_s2[294], state_out_s1[294], state_out_s0[294]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1507 ( .a ({new_AGEMA_signal_4598, new_AGEMA_signal_4597, rd_I_n2332}), .b ({new_AGEMA_signal_3890, new_AGEMA_signal_3889, rd_I_n2564}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_5354, new_AGEMA_signal_5353, rd_I_n2333}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1505 ( .a ({new_AGEMA_signal_5356, new_AGEMA_signal_5355, rd_I_n2331}), .b ({new_AGEMA_signal_3816, new_AGEMA_signal_3815, rd_I_n2330}), .c ({state_out_s2[60], state_out_s1[60], state_out_s0[60]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1504 ( .a ({new_AGEMA_signal_4600, new_AGEMA_signal_4599, rd_I_n2329}), .b ({new_AGEMA_signal_3818, new_AGEMA_signal_3817, rd_I_n2328}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_5356, new_AGEMA_signal_5355, rd_I_n2331}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1502 ( .a ({new_AGEMA_signal_4442, new_AGEMA_signal_4441, rd_I_n2326}), .b ({new_AGEMA_signal_4602, new_AGEMA_signal_4601, rd_I_n2325}), .c ({state_out_s2[37], state_out_s1[37], state_out_s0[37]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1501 ( .a ({new_AGEMA_signal_4444, new_AGEMA_signal_4443, rd_I_n2324}), .b ({new_AGEMA_signal_4440, new_AGEMA_signal_4439, rd_I_n2323}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_4602, new_AGEMA_signal_4601, rd_I_n2325}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1500 ( .a ({new_AGEMA_signal_4046, new_AGEMA_signal_4045, rd_I_n2322}), .b ({new_AGEMA_signal_4604, new_AGEMA_signal_4603, rd_I_n2321}), .c ({state_out_s2[221], state_out_s1[221], state_out_s0[221]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1499 ( .a ({new_AGEMA_signal_4048, new_AGEMA_signal_4047, rd_I_n2320}), .b ({new_AGEMA_signal_4044, new_AGEMA_signal_4043, rd_I_n2319}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_4604, new_AGEMA_signal_4603, rd_I_n2321}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1498 ( .a ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, rd_I_n2318}), .b ({new_AGEMA_signal_4260, new_AGEMA_signal_4259, rd_I_n2317}), .c ({state_out_s2[198], state_out_s1[198], state_out_s0[198]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1497 ( .a ({new_AGEMA_signal_4606, new_AGEMA_signal_4605, rd_I_n2316}), .b ({new_AGEMA_signal_4262, new_AGEMA_signal_4261, rd_I_n2315}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_5362, new_AGEMA_signal_5361, rd_I_n2318}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1495 ( .a ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, rd_I_n2313}), .b ({new_AGEMA_signal_4080, new_AGEMA_signal_4079, rd_I_n2312}), .c ({state_out_s2[376], state_out_s1[376], state_out_s0[376]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1494 ( .a ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, rd_I_n2311}), .b ({new_AGEMA_signal_4082, new_AGEMA_signal_4081, rd_I_n2310}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, rd_I_n2313}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1492 ( .a ({new_AGEMA_signal_5366, new_AGEMA_signal_5365, rd_I_n2308}), .b ({new_AGEMA_signal_4114, new_AGEMA_signal_4113, rd_I_n2419}), .c ({state_out_s2[367], state_out_s1[367], state_out_s0[367]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1491 ( .a ({new_AGEMA_signal_4610, new_AGEMA_signal_4609, rd_I_n2307}), .b ({new_AGEMA_signal_4112, new_AGEMA_signal_4111, rd_I_n2422}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_5366, new_AGEMA_signal_5365, rd_I_n2308}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1489 ( .a ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, rd_I_n2306}), .b ({new_AGEMA_signal_3918, new_AGEMA_signal_3917, rd_I_n2305}), .c ({state_out_s2[120], state_out_s1[120], state_out_s0[120]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1488 ( .a ({new_AGEMA_signal_4612, new_AGEMA_signal_4611, rd_I_n2304}), .b ({new_AGEMA_signal_3920, new_AGEMA_signal_3919, rd_I_n2303}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_5368, new_AGEMA_signal_5367, rd_I_n2306}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1486 ( .a ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, rd_I_n2301}), .b ({new_AGEMA_signal_3996, new_AGEMA_signal_3995, rd_I_n2300}), .c ({state_out_s2[111], state_out_s1[111], state_out_s0[111]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1485 ( .a ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, rd_I_n2299}), .b ({new_AGEMA_signal_3998, new_AGEMA_signal_3997, rd_I_n2298}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, rd_I_n2301}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1483 ( .a ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, rd_I_n2385}), .b ({new_AGEMA_signal_5372, new_AGEMA_signal_5371, rd_I_n2296}), .c ({state_out_s2[153], state_out_s1[153], state_out_s0[153]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1482 ( .a ({new_AGEMA_signal_3708, new_AGEMA_signal_3707, rd_I_n2384}), .b ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, rd_I_n2387}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_5372, new_AGEMA_signal_5371, rd_I_n2296}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1481 ( .a ({new_AGEMA_signal_5374, new_AGEMA_signal_5373, rd_I_n2295}), .b ({new_AGEMA_signal_4362, new_AGEMA_signal_4361, rd_I_n2294}), .c ({state_out_s2[144], state_out_s1[144], state_out_s0[144]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1480 ( .a ({new_AGEMA_signal_4616, new_AGEMA_signal_4615, rd_I_n2293}), .b ({new_AGEMA_signal_4364, new_AGEMA_signal_4363, rd_I_n2292}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_5374, new_AGEMA_signal_5373, rd_I_n2295}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1478 ( .a ({new_AGEMA_signal_4346, new_AGEMA_signal_4345, rd_I_n2290}), .b ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, rd_I_n2289}), .c ({state_out_s2[299], state_out_s1[299], state_out_s0[299]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1477 ( .a ({new_AGEMA_signal_4344, new_AGEMA_signal_4343, rd_I_n2288}), .b ({new_AGEMA_signal_4348, new_AGEMA_signal_4347, rd_I_n2287}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_4618, new_AGEMA_signal_4617, rd_I_n2289}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1476 ( .a ({new_AGEMA_signal_4334, new_AGEMA_signal_4333, rd_I_n2286}), .b ({new_AGEMA_signal_4620, new_AGEMA_signal_4619, rd_I_n2285}), .c ({state_out_s2[290], state_out_s1[290], state_out_s0[290]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1475 ( .a ({new_AGEMA_signal_4332, new_AGEMA_signal_4331, rd_I_n2284}), .b ({new_AGEMA_signal_4336, new_AGEMA_signal_4335, rd_I_n2283}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_4620, new_AGEMA_signal_4619, rd_I_n2285}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1474 ( .a ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, rd_I_n2282}), .b ({new_AGEMA_signal_3906, new_AGEMA_signal_3905, rd_I_n2281}), .c ({state_out_s2[59], state_out_s1[59], state_out_s0[59]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1473 ( .a ({new_AGEMA_signal_4622, new_AGEMA_signal_4621, rd_I_n2280}), .b ({new_AGEMA_signal_3908, new_AGEMA_signal_3907, rd_I_n2279}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_5380, new_AGEMA_signal_5379, rd_I_n2282}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1471 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, rd_I_n2277}), .b ({new_AGEMA_signal_3900, new_AGEMA_signal_3899, rd_I_n2276}), .c ({state_out_s2[36], state_out_s1[36], state_out_s0[36]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1470 ( .a ({new_AGEMA_signal_4624, new_AGEMA_signal_4623, rd_I_n2275}), .b ({new_AGEMA_signal_3902, new_AGEMA_signal_3901, rd_I_n2274}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, rd_I_n2277}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1468 ( .a ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, rd_I_n2467}), .b ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, rd_I_n2272}), .c ({state_out_s2[220], state_out_s1[220], state_out_s0[220]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1467 ( .a ({new_AGEMA_signal_3706, new_AGEMA_signal_3705, rd_I_n2466}), .b ({new_AGEMA_signal_3702, new_AGEMA_signal_3701, rd_I_n2469}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, rd_I_n2272}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1466 ( .a ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, rd_I_n2462}), .b ({new_AGEMA_signal_4628, new_AGEMA_signal_4627, rd_I_n2271}), .c ({state_out_s2[197], state_out_s1[197], state_out_s0[197]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1465 ( .a ({new_AGEMA_signal_3700, new_AGEMA_signal_3699, rd_I_n2461}), .b ({new_AGEMA_signal_3696, new_AGEMA_signal_3695, rd_I_n2464}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_4628, new_AGEMA_signal_4627, rd_I_n2271}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1464 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, rd_I_n2270}), .b ({new_AGEMA_signal_4368, new_AGEMA_signal_4367, rd_I_n2269}), .c ({state_out_s2[375], state_out_s1[375], state_out_s0[375]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1463 ( .a ({new_AGEMA_signal_4630, new_AGEMA_signal_4629, rd_I_n2268}), .b ({new_AGEMA_signal_4370, new_AGEMA_signal_4369, rd_I_n2267}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, rd_I_n2270}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1461 ( .a ({new_AGEMA_signal_5390, new_AGEMA_signal_5389, rd_I_n2265}), .b ({new_AGEMA_signal_4030, new_AGEMA_signal_4029, rd_I_n2367}), .c ({state_out_s2[366], state_out_s1[366], state_out_s0[366]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1460 ( .a ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, rd_I_n2264}), .b ({new_AGEMA_signal_4028, new_AGEMA_signal_4027, rd_I_n2370}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_5390, new_AGEMA_signal_5389, rd_I_n2265}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1458 ( .a ({new_AGEMA_signal_5392, new_AGEMA_signal_5391, rd_I_n2263}), .b ({new_AGEMA_signal_4342, new_AGEMA_signal_4341, rd_I_n2262}), .c ({state_out_s2[101], state_out_s1[101], state_out_s0[101]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1457 ( .a ({new_AGEMA_signal_4634, new_AGEMA_signal_4633, rd_I_n2261}), .b ({new_AGEMA_signal_4340, new_AGEMA_signal_4339, rd_I_n2260}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_5392, new_AGEMA_signal_5391, rd_I_n2263}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1455 ( .a ({new_AGEMA_signal_5394, new_AGEMA_signal_5393, rd_I_n2258}), .b ({new_AGEMA_signal_4434, new_AGEMA_signal_4433, rd_I_n2257}), .c ({state_out_s2[134], state_out_s1[134], state_out_s0[134]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1454 ( .a ({new_AGEMA_signal_4636, new_AGEMA_signal_4635, rd_I_n2256}), .b ({new_AGEMA_signal_4436, new_AGEMA_signal_4435, rd_I_n2255}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_5394, new_AGEMA_signal_5393, rd_I_n2258}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1452 ( .a ({new_AGEMA_signal_4304, new_AGEMA_signal_4303, rd_I_n2253}), .b ({new_AGEMA_signal_4638, new_AGEMA_signal_4637, rd_I_n2252}), .c ({state_out_s2[312], state_out_s1[312], state_out_s0[312]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1451 ( .a ({new_AGEMA_signal_4302, new_AGEMA_signal_4301, rd_I_n2251}), .b ({new_AGEMA_signal_4306, new_AGEMA_signal_4305, rd_I_n2250}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_4638, new_AGEMA_signal_4637, rd_I_n2252}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1450 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, rd_I_n2249}), .b ({new_AGEMA_signal_3882, new_AGEMA_signal_3881, rd_I_n2248}), .c ({state_out_s2[97], state_out_s1[97], state_out_s0[97]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1449 ( .a ({new_AGEMA_signal_4640, new_AGEMA_signal_4639, rd_I_n2247}), .b ({new_AGEMA_signal_3884, new_AGEMA_signal_3883, rd_I_n2246}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_5398, new_AGEMA_signal_5397, rd_I_n2249}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1447 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, rd_I_n2244}), .b ({new_AGEMA_signal_3690, new_AGEMA_signal_3689, rd_I_n2587}), .c ({state_out_s2[130], state_out_s1[130], state_out_s0[130]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1445 ( .a ({new_AGEMA_signal_3694, new_AGEMA_signal_3693, rd_I_n2590}), .b ({new_AGEMA_signal_4642, new_AGEMA_signal_4641, rd_I_n2588}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, rd_I_n2244}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1441 ( .a ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, rd_I_n2239}), .b ({new_AGEMA_signal_4156, new_AGEMA_signal_4155, rd_I_n2238}), .c ({state_out_s2[308], state_out_s1[308], state_out_s0[308]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1440 ( .a ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, rd_I_n2237}), .b ({new_AGEMA_signal_4154, new_AGEMA_signal_4153, rd_I_n2236}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_5402, new_AGEMA_signal_5401, rd_I_n2239}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1438 ( .a ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, rd_I_n2234}), .b ({new_AGEMA_signal_4102, new_AGEMA_signal_4101, rd_I_n2233}), .c ({state_out_s2[89], state_out_s1[89], state_out_s0[89]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1437 ( .a ({new_AGEMA_signal_4646, new_AGEMA_signal_4645, rd_I_n2232}), .b ({new_AGEMA_signal_4100, new_AGEMA_signal_4099, rd_I_n2231}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_5404, new_AGEMA_signal_5403, rd_I_n2234}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1435 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, rd_I_n2229}), .b ({new_AGEMA_signal_4270, new_AGEMA_signal_4269, rd_I_n2228}), .c ({state_out_s2[80], state_out_s1[80], state_out_s0[80]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1434 ( .a ({new_AGEMA_signal_4648, new_AGEMA_signal_4647, rd_I_n2227}), .b ({new_AGEMA_signal_4268, new_AGEMA_signal_4267, rd_I_n2226}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, rd_I_n2229}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1432 ( .a ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, rd_I_n2224}), .b ({new_AGEMA_signal_4420, new_AGEMA_signal_4419, rd_I_n2223}), .c ({state_out_s2[250], state_out_s1[250], state_out_s0[250]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1431 ( .a ({new_AGEMA_signal_4650, new_AGEMA_signal_4649, rd_I_n2222}), .b ({new_AGEMA_signal_4418, new_AGEMA_signal_4417, rd_I_n2221}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_5408, new_AGEMA_signal_5407, rd_I_n2224}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1429 ( .a ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, rd_I_n2219}), .b ({new_AGEMA_signal_4306, new_AGEMA_signal_4305, rd_I_n2250}), .c ({state_out_s2[241], state_out_s1[241], state_out_s0[241]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1428 ( .a ({new_AGEMA_signal_4652, new_AGEMA_signal_4651, rd_I_n2218}), .b ({new_AGEMA_signal_4304, new_AGEMA_signal_4303, rd_I_n2253}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_5410, new_AGEMA_signal_5409, rd_I_n2219}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1426 ( .a ({new_AGEMA_signal_3700, new_AGEMA_signal_3699, rd_I_n2461}), .b ({new_AGEMA_signal_4654, new_AGEMA_signal_4653, rd_I_n2217}), .c ({state_out_s2[268], state_out_s1[268], state_out_s0[268]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1425 ( .a ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, rd_I_n2462}), .b ({new_AGEMA_signal_3696, new_AGEMA_signal_3695, rd_I_n2464}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_4654, new_AGEMA_signal_4653, rd_I_n2217}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1421 ( .a ({new_AGEMA_signal_3706, new_AGEMA_signal_3705, rd_I_n2466}), .b ({new_AGEMA_signal_4656, new_AGEMA_signal_4655, rd_I_n2213}), .c ({state_out_s2[259], state_out_s1[259], state_out_s0[259]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1420 ( .a ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, rd_I_n2467}), .b ({new_AGEMA_signal_3702, new_AGEMA_signal_3701, rd_I_n2469}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_4656, new_AGEMA_signal_4655, rd_I_n2213}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1416 ( .a ({new_AGEMA_signal_5416, new_AGEMA_signal_5415, rd_I_n2209}), .b ({new_AGEMA_signal_3930, new_AGEMA_signal_3929, rd_I_n2208}), .c ({state_out_s2[58], state_out_s1[58], state_out_s0[58]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1415 ( .a ({new_AGEMA_signal_4658, new_AGEMA_signal_4657, rd_I_n2207}), .b ({new_AGEMA_signal_3932, new_AGEMA_signal_3931, rd_I_n2206}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_5416, new_AGEMA_signal_5415, rd_I_n2209}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1413 ( .a ({new_AGEMA_signal_3830, new_AGEMA_signal_3829, rd_I_n2204}), .b ({new_AGEMA_signal_4660, new_AGEMA_signal_4659, rd_I_n2203}), .c ({state_out_s2[35], state_out_s1[35], state_out_s0[35]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1412 ( .a ({new_AGEMA_signal_3832, new_AGEMA_signal_3831, rd_I_n2202}), .b ({new_AGEMA_signal_3828, new_AGEMA_signal_3827, rd_I_n2201}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_4660, new_AGEMA_signal_4659, rd_I_n2203}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1411 ( .a ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, rd_I_n2200}), .b ({new_AGEMA_signal_4036, new_AGEMA_signal_4035, rd_I_n2199}), .c ({state_out_s2[219], state_out_s1[219], state_out_s0[219]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1410 ( .a ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, rd_I_n2198}), .b ({new_AGEMA_signal_4034, new_AGEMA_signal_4033, rd_I_n2197}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_5420, new_AGEMA_signal_5419, rd_I_n2200}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1408 ( .a ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, rd_I_n2195}), .b ({new_AGEMA_signal_4166, new_AGEMA_signal_4165, rd_I_n2194}), .c ({state_out_s2[196], state_out_s1[196], state_out_s0[196]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1407 ( .a ({new_AGEMA_signal_4664, new_AGEMA_signal_4663, rd_I_n2193}), .b ({new_AGEMA_signal_4168, new_AGEMA_signal_4167, rd_I_n2192}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_5422, new_AGEMA_signal_5421, rd_I_n2195}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1405 ( .a ({new_AGEMA_signal_3968, new_AGEMA_signal_3967, rd_I_n2501}), .b ({new_AGEMA_signal_4666, new_AGEMA_signal_4665, rd_I_n2190}), .c ({state_out_s2[374], state_out_s1[374], state_out_s0[374]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1404 ( .a ({new_AGEMA_signal_3970, new_AGEMA_signal_3969, rd_I_n2500}), .b ({new_AGEMA_signal_3966, new_AGEMA_signal_3965, rd_I_n2503}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_4666, new_AGEMA_signal_4665, rd_I_n2190}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1403 ( .a ({new_AGEMA_signal_5426, new_AGEMA_signal_5425, rd_I_n2189}), .b ({new_AGEMA_signal_4440, new_AGEMA_signal_4439, rd_I_n2323}), .c ({state_out_s2[365], state_out_s1[365], state_out_s0[365]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1402 ( .a ({new_AGEMA_signal_4668, new_AGEMA_signal_4667, rd_I_n2188}), .b ({new_AGEMA_signal_4442, new_AGEMA_signal_4441, rd_I_n2326}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_5426, new_AGEMA_signal_5425, rd_I_n2189}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1400 ( .a ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, rd_I_n2187}), .b ({new_AGEMA_signal_3720, new_AGEMA_signal_3719, rd_I_n2380}), .c ({state_out_s2[56], state_out_s1[56], state_out_s0[56]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1399 ( .a ({new_AGEMA_signal_4670, new_AGEMA_signal_4669, rd_I_n2186}), .b ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, rd_I_n2383}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_5428, new_AGEMA_signal_5427, rd_I_n2187}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1397 ( .a ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, rd_I_n2185}), .b ({new_AGEMA_signal_3714, new_AGEMA_signal_3713, rd_I_n2526}), .c ({state_out_s2[33], state_out_s1[33], state_out_s0[33]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1396 ( .a ({new_AGEMA_signal_4672, new_AGEMA_signal_4671, rd_I_n2184}), .b ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, rd_I_n2529}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, rd_I_n2185}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1394 ( .a ({new_AGEMA_signal_4010, new_AGEMA_signal_4009, rd_I_n2183}), .b ({new_AGEMA_signal_4674, new_AGEMA_signal_4673, rd_I_n2182}), .c ({state_out_s2[217], state_out_s1[217], state_out_s0[217]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1393 ( .a ({new_AGEMA_signal_4008, new_AGEMA_signal_4007, rd_I_n2181}), .b ({new_AGEMA_signal_4012, new_AGEMA_signal_4011, rd_I_n2180}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_4674, new_AGEMA_signal_4673, rd_I_n2182}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1392 ( .a ({new_AGEMA_signal_3848, new_AGEMA_signal_3847, rd_I_n2179}), .b ({new_AGEMA_signal_4676, new_AGEMA_signal_4675, rd_I_n2178}), .c ({state_out_s2[194], state_out_s1[194], state_out_s0[194]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1391 ( .a ({new_AGEMA_signal_3846, new_AGEMA_signal_3845, rd_I_n2177}), .b ({new_AGEMA_signal_3850, new_AGEMA_signal_3849, rd_I_n2176}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_4676, new_AGEMA_signal_4675, rd_I_n2178}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1390 ( .a ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, rd_I_n2175}), .b ({new_AGEMA_signal_3822, new_AGEMA_signal_3821, rd_I_n2174}), .c ({state_out_s2[372], state_out_s1[372], state_out_s0[372]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1389 ( .a ({new_AGEMA_signal_4678, new_AGEMA_signal_4677, rd_I_n2173}), .b ({new_AGEMA_signal_3824, new_AGEMA_signal_3823, rd_I_n2172}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, rd_I_n2175}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1387 ( .a ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, rd_I_n2170}), .b ({new_AGEMA_signal_3828, new_AGEMA_signal_3827, rd_I_n2201}), .c ({state_out_s2[363], state_out_s1[363], state_out_s0[363]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1386 ( .a ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, rd_I_n2169}), .b ({new_AGEMA_signal_3830, new_AGEMA_signal_3829, rd_I_n2204}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_5438, new_AGEMA_signal_5437, rd_I_n2170}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1384 ( .a ({new_AGEMA_signal_4388, new_AGEMA_signal_4387, rd_I_n2406}), .b ({new_AGEMA_signal_4682, new_AGEMA_signal_4681, rd_I_n2168}), .c ({state_out_s2[50], state_out_s1[50], state_out_s0[50]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1383 ( .a ({new_AGEMA_signal_4390, new_AGEMA_signal_4389, rd_I_n2405}), .b ({new_AGEMA_signal_4386, new_AGEMA_signal_4385, rd_I_n2408}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_4682, new_AGEMA_signal_4681, rd_I_n2168}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1382 ( .a ({new_AGEMA_signal_4142, new_AGEMA_signal_4141, rd_I_n2167}), .b ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, rd_I_n2166}), .c ({state_out_s2[211], state_out_s1[211], state_out_s0[211]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1381 ( .a ({new_AGEMA_signal_4144, new_AGEMA_signal_4143, rd_I_n2165}), .b ({new_AGEMA_signal_4140, new_AGEMA_signal_4139, rd_I_n2164}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_4684, new_AGEMA_signal_4683, rd_I_n2166}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1380 ( .a ({new_AGEMA_signal_5444, new_AGEMA_signal_5443, rd_I_n2163}), .b ({new_AGEMA_signal_3780, new_AGEMA_signal_3779, rd_I_n2371}), .c ({state_out_s2[357], state_out_s1[357], state_out_s0[357]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1379 ( .a ({new_AGEMA_signal_4686, new_AGEMA_signal_4685, rd_I_n2162}), .b ({new_AGEMA_signal_3782, new_AGEMA_signal_3781, rd_I_n2374}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_5444, new_AGEMA_signal_5443, rd_I_n2163}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1377 ( .a ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, rd_I_n2161}), .b ({new_AGEMA_signal_4946, new_AGEMA_signal_4945, rd_I_n2160}), .c ({state_out_s2[13], state_out_s1[13], state_out_s0[13]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1376 ( .a ({new_AGEMA_signal_4688, new_AGEMA_signal_4687, rd_I_n2159}), .b ({new_AGEMA_signal_3938, new_AGEMA_signal_3937, rd_I_n2158}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_5446, new_AGEMA_signal_5445, rd_I_n2161}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1374 ( .a ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, rd_I_n2156}), .b ({new_AGEMA_signal_4090, new_AGEMA_signal_4089, rd_I_n2155}), .c ({state_out_s2[4], state_out_s1[4], state_out_s0[4]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1373 ( .a ({new_AGEMA_signal_4690, new_AGEMA_signal_4689, rd_I_n2154}), .b ({new_AGEMA_signal_4088, new_AGEMA_signal_4087, rd_I_n2153}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, rd_I_n2156}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1371 ( .a ({new_AGEMA_signal_3788, new_AGEMA_signal_3787, rd_I_n2151}), .b ({new_AGEMA_signal_4692, new_AGEMA_signal_4691, rd_I_n2150}), .c ({state_out_s2[174], state_out_s1[174], state_out_s0[174]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1370 ( .a ({new_AGEMA_signal_3790, new_AGEMA_signal_3789, rd_I_n2149}), .b ({new_AGEMA_signal_3786, new_AGEMA_signal_3785, rd_I_n2148}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_4692, new_AGEMA_signal_4691, rd_I_n2150}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1369 ( .a ({new_AGEMA_signal_3902, new_AGEMA_signal_3901, rd_I_n2274}), .b ({new_AGEMA_signal_4694, new_AGEMA_signal_4693, rd_I_n2147}), .c ({state_out_s2[165], state_out_s1[165], state_out_s0[165]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1368 ( .a ({new_AGEMA_signal_3904, new_AGEMA_signal_3903, rd_I_n2273}), .b ({new_AGEMA_signal_3900, new_AGEMA_signal_3899, rd_I_n2276}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_4694, new_AGEMA_signal_4693, rd_I_n2147}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1367 ( .a ({new_AGEMA_signal_4364, new_AGEMA_signal_4363, rd_I_n2292}), .b ({new_AGEMA_signal_4696, new_AGEMA_signal_4695, rd_I_n2146}), .c ({state_out_s2[343], state_out_s1[343], state_out_s0[343]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1366 ( .a ({new_AGEMA_signal_4366, new_AGEMA_signal_4365, rd_I_n2291}), .b ({new_AGEMA_signal_4362, new_AGEMA_signal_4361, rd_I_n2294}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_4696, new_AGEMA_signal_4695, rd_I_n2146}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1365 ( .a ({new_AGEMA_signal_5456, new_AGEMA_signal_5455, rd_I_n2145}), .b ({new_AGEMA_signal_3708, new_AGEMA_signal_3707, rd_I_n2384}), .c ({state_out_s2[320], state_out_s1[320], state_out_s0[320]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1363 ( .a ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, rd_I_n2387}), .b ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, rd_I_n2385}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_5456, new_AGEMA_signal_5455, rd_I_n2145}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1359 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, rd_I_n2140}), .b ({new_AGEMA_signal_3738, new_AGEMA_signal_3737, rd_I_n2592}), .c ({state_out_s2[54], state_out_s1[54], state_out_s0[54]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1358 ( .a ({new_AGEMA_signal_4700, new_AGEMA_signal_4699, rd_I_n2139}), .b ({new_AGEMA_signal_3740, new_AGEMA_signal_3739, rd_I_n2595}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_5458, new_AGEMA_signal_5457, rd_I_n2140}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1356 ( .a ({new_AGEMA_signal_4190, new_AGEMA_signal_4189, rd_I_n2138}), .b ({new_AGEMA_signal_4702, new_AGEMA_signal_4701, rd_I_n2137}), .c ({state_out_s2[215], state_out_s1[215], state_out_s0[215]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1355 ( .a ({new_AGEMA_signal_4188, new_AGEMA_signal_4187, rd_I_n2136}), .b ({new_AGEMA_signal_4192, new_AGEMA_signal_4191, rd_I_n2135}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_4702, new_AGEMA_signal_4701, rd_I_n2137}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1354 ( .a ({new_AGEMA_signal_3718, new_AGEMA_signal_3717, rd_I_n2527}), .b ({new_AGEMA_signal_4704, new_AGEMA_signal_4703, rd_I_n2134}), .c ({state_out_s2[361], state_out_s1[361], state_out_s0[361]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1353 ( .a ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, rd_I_n2529}), .b ({new_AGEMA_signal_3714, new_AGEMA_signal_3713, rd_I_n2526}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_4704, new_AGEMA_signal_4703, rd_I_n2134}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1349 ( .a ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, rd_I_n2131}), .b ({new_AGEMA_signal_3786, new_AGEMA_signal_3785, rd_I_n2148}), .c ({state_out_s2[45], state_out_s1[45], state_out_s0[45]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1348 ( .a ({new_AGEMA_signal_4706, new_AGEMA_signal_4705, rd_I_n2130}), .b ({new_AGEMA_signal_3788, new_AGEMA_signal_3787, rd_I_n2151}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_5464, new_AGEMA_signal_5463, rd_I_n2131}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1346 ( .a ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, rd_I_n2129}), .b ({new_AGEMA_signal_4006, new_AGEMA_signal_4005, rd_I_n2128}), .c ({state_out_s2[206], state_out_s1[206], state_out_s0[206]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1345 ( .a ({new_AGEMA_signal_4708, new_AGEMA_signal_4707, rd_I_n2127}), .b ({new_AGEMA_signal_4004, new_AGEMA_signal_4003, rd_I_n2126}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, rd_I_n2129}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1343 ( .a ({new_AGEMA_signal_3724, new_AGEMA_signal_3723, rd_I_n2381}), .b ({new_AGEMA_signal_4710, new_AGEMA_signal_4709, rd_I_n2124}), .c ({state_out_s2[352], state_out_s1[352], state_out_s0[352]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1342 ( .a ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, rd_I_n2383}), .b ({new_AGEMA_signal_3720, new_AGEMA_signal_3719, rd_I_n2380}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_4710, new_AGEMA_signal_4709, rd_I_n2124}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1338 ( .a ({new_AGEMA_signal_5470, new_AGEMA_signal_5469, rd_I_n2121}), .b ({new_AGEMA_signal_3792, new_AGEMA_signal_3791, rd_I_n2120}), .c ({state_out_s2[66], state_out_s1[66], state_out_s0[66]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1337 ( .a ({new_AGEMA_signal_4712, new_AGEMA_signal_4711, rd_I_n2119}), .b ({new_AGEMA_signal_3794, new_AGEMA_signal_3793, rd_I_n2118}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_5470, new_AGEMA_signal_5469, rd_I_n2121}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1335 ( .a ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, rd_I_n2116}), .b ({new_AGEMA_signal_4402, new_AGEMA_signal_4401, rd_I_n2115}), .c ({state_out_s2[227], state_out_s1[227], state_out_s0[227]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1334 ( .a ({new_AGEMA_signal_4714, new_AGEMA_signal_4713, rd_I_n2114}), .b ({new_AGEMA_signal_4400, new_AGEMA_signal_4399, rd_I_n2113}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, rd_I_n2116}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1332 ( .a ({new_AGEMA_signal_4004, new_AGEMA_signal_4003, rd_I_n2126}), .b ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, rd_I_n2111}), .c ({state_out_s2[277], state_out_s1[277], state_out_s0[277]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1331 ( .a ({new_AGEMA_signal_4002, new_AGEMA_signal_4001, rd_I_n2125}), .b ({new_AGEMA_signal_4006, new_AGEMA_signal_4005, rd_I_n2128}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, rd_I_n2111}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1330 ( .a ({new_AGEMA_signal_5144, new_AGEMA_signal_5143, rd_I_n2110}), .b ({new_AGEMA_signal_4718, new_AGEMA_signal_4717, rd_I_n2109}), .c ({state_out_s2[17], state_out_s1[17], state_out_s0[17]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1329 ( .a ({new_AGEMA_signal_4282, new_AGEMA_signal_4281, rd_I_n2108}), .b ({new_AGEMA_signal_4278, new_AGEMA_signal_4277, rd_I_n2107}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_4718, new_AGEMA_signal_4717, rd_I_n2109}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1328 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, rd_I_n2106}), .b ({new_AGEMA_signal_3810, new_AGEMA_signal_3809, rd_I_n2357}), .c ({state_out_s2[178], state_out_s1[178], state_out_s0[178]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1327 ( .a ({new_AGEMA_signal_4720, new_AGEMA_signal_4719, rd_I_n2105}), .b ({new_AGEMA_signal_3812, new_AGEMA_signal_3811, rd_I_n2360}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, rd_I_n2106}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1325 ( .a ({new_AGEMA_signal_3806, new_AGEMA_signal_3805, rd_I_n2339}), .b ({new_AGEMA_signal_4722, new_AGEMA_signal_4721, rd_I_n2104}), .c ({state_out_s2[324], state_out_s1[324], state_out_s0[324]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1324 ( .a ({new_AGEMA_signal_3808, new_AGEMA_signal_3807, rd_I_n2338}), .b ({new_AGEMA_signal_3804, new_AGEMA_signal_3803, rd_I_n2341}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_4722, new_AGEMA_signal_4721, rd_I_n2104}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1323 ( .a ({new_AGEMA_signal_3730, new_AGEMA_signal_3729, rd_I_n2574}), .b ({new_AGEMA_signal_4724, new_AGEMA_signal_4723, rd_I_n2103}), .c ({state_out_s2[52], state_out_s1[52], state_out_s0[52]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1322 ( .a ({new_AGEMA_signal_3728, new_AGEMA_signal_3727, rd_I_n2575}), .b ({new_AGEMA_signal_3726, new_AGEMA_signal_3725, rd_I_n2577}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_4724, new_AGEMA_signal_4723, rd_I_n2103}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1318 ( .a ({new_AGEMA_signal_3736, new_AGEMA_signal_3735, rd_I_n2569}), .b ({new_AGEMA_signal_4726, new_AGEMA_signal_4725, rd_I_n2099}), .c ({state_out_s2[43], state_out_s1[43], state_out_s0[43]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1317 ( .a ({new_AGEMA_signal_3734, new_AGEMA_signal_3733, rd_I_n2570}), .b ({new_AGEMA_signal_3732, new_AGEMA_signal_3731, rd_I_n2572}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_4726, new_AGEMA_signal_4725, rd_I_n2099}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1313 ( .a ({new_AGEMA_signal_4234, new_AGEMA_signal_4233, rd_I_n2095}), .b ({new_AGEMA_signal_4728, new_AGEMA_signal_4727, rd_I_n2094}), .c ({state_out_s2[213], state_out_s1[213], state_out_s0[213]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1312 ( .a ({new_AGEMA_signal_4230, new_AGEMA_signal_4229, rd_I_n2093}), .b ({new_AGEMA_signal_4232, new_AGEMA_signal_4231, rd_I_n2092}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_4728, new_AGEMA_signal_4727, rd_I_n2094}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1311 ( .a ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, rd_I_n2091}), .b ({new_AGEMA_signal_4180, new_AGEMA_signal_4179, rd_I_n2090}), .c ({state_out_s2[204], state_out_s1[204], state_out_s0[204]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1310 ( .a ({new_AGEMA_signal_4730, new_AGEMA_signal_4729, rd_I_n2089}), .b ({new_AGEMA_signal_4178, new_AGEMA_signal_4177, rd_I_n2088}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_5488, new_AGEMA_signal_5487, rd_I_n2091}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1308 ( .a ({new_AGEMA_signal_3742, new_AGEMA_signal_3741, rd_I_n2593}), .b ({new_AGEMA_signal_4732, new_AGEMA_signal_4731, rd_I_n2086}), .c ({state_out_s2[382], state_out_s1[382], state_out_s0[382]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1307 ( .a ({new_AGEMA_signal_3740, new_AGEMA_signal_3739, rd_I_n2595}), .b ({new_AGEMA_signal_3738, new_AGEMA_signal_3737, rd_I_n2592}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_4732, new_AGEMA_signal_4731, rd_I_n2086}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1303 ( .a ({new_AGEMA_signal_3748, new_AGEMA_signal_3747, rd_I_n2610}), .b ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, rd_I_n2085}), .c ({state_out_s2[359], state_out_s1[359], state_out_s0[359]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1302 ( .a ({new_AGEMA_signal_3746, new_AGEMA_signal_3745, rd_I_n2612}), .b ({new_AGEMA_signal_3744, new_AGEMA_signal_3743, rd_I_n2609}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, rd_I_n2085}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1298 ( .a ({new_AGEMA_signal_5494, new_AGEMA_signal_5493, rd_I_n2082}), .b ({new_AGEMA_signal_3994, new_AGEMA_signal_3993, rd_I_n2363}), .c ({state_out_s2[93], state_out_s1[93], state_out_s0[93]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1297 ( .a ({new_AGEMA_signal_4736, new_AGEMA_signal_4735, rd_I_n2081}), .b ({new_AGEMA_signal_3992, new_AGEMA_signal_3991, rd_I_n2366}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_5494, new_AGEMA_signal_5493, rd_I_n2082}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1295 ( .a ({new_AGEMA_signal_3754, new_AGEMA_signal_3753, rd_I_n2446}), .b ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, rd_I_n2080}), .c ({state_out_s2[70], state_out_s1[70], state_out_s0[70]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1294 ( .a ({new_AGEMA_signal_3752, new_AGEMA_signal_3751, rd_I_n2448}), .b ({new_AGEMA_signal_3750, new_AGEMA_signal_3749, rd_I_n2445}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_4738, new_AGEMA_signal_4737, rd_I_n2080}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1290 ( .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, rd_I_n2077}), .b ({new_AGEMA_signal_4258, new_AGEMA_signal_4257, rd_I_n2076}), .c ({state_out_s2[254], state_out_s1[254], state_out_s0[254]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1289 ( .a ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, rd_I_n2075}), .b ({new_AGEMA_signal_4256, new_AGEMA_signal_4255, rd_I_n2074}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_5498, new_AGEMA_signal_5497, rd_I_n2077}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1287 ( .a ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, rd_I_n2072}), .b ({new_AGEMA_signal_4314, new_AGEMA_signal_4313, rd_I_n2071}), .c ({state_out_s2[231], state_out_s1[231], state_out_s0[231]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1286 ( .a ({new_AGEMA_signal_4742, new_AGEMA_signal_4741, rd_I_n2070}), .b ({new_AGEMA_signal_4316, new_AGEMA_signal_4315, rd_I_n2069}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_5500, new_AGEMA_signal_5499, rd_I_n2072}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1284 ( .a ({new_AGEMA_signal_4040, new_AGEMA_signal_4039, rd_I_n2067}), .b ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, rd_I_n2066}), .c ({state_out_s2[281], state_out_s1[281], state_out_s0[281]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1283 ( .a ({new_AGEMA_signal_4038, new_AGEMA_signal_4037, rd_I_n2065}), .b ({new_AGEMA_signal_4042, new_AGEMA_signal_4041, rd_I_n2064}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_4744, new_AGEMA_signal_4743, rd_I_n2066}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1282 ( .a ({new_AGEMA_signal_4016, new_AGEMA_signal_4015, rd_I_n2437}), .b ({new_AGEMA_signal_4746, new_AGEMA_signal_4745, rd_I_n2063}), .c ({state_out_s2[272], state_out_s1[272], state_out_s0[272]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1281 ( .a ({new_AGEMA_signal_4014, new_AGEMA_signal_4013, rd_I_n2436}), .b ({new_AGEMA_signal_4018, new_AGEMA_signal_4017, rd_I_n2439}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_4746, new_AGEMA_signal_4745, rd_I_n2063}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1280 ( .a ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, rd_I_n2062}), .b ({new_AGEMA_signal_4748, new_AGEMA_signal_4747, rd_I_n2061}), .c ({state_out_s2[53], state_out_s1[53], state_out_s0[53]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1279 ( .a ({new_AGEMA_signal_3862, new_AGEMA_signal_3861, rd_I_n2060}), .b ({new_AGEMA_signal_3858, new_AGEMA_signal_3857, rd_I_n2059}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_4748, new_AGEMA_signal_4747, rd_I_n2061}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1278 ( .a ({new_AGEMA_signal_4208, new_AGEMA_signal_4207, rd_I_n2058}), .b ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, rd_I_n2057}), .c ({state_out_s2[214], state_out_s1[214], state_out_s0[214]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1277 ( .a ({new_AGEMA_signal_4206, new_AGEMA_signal_4205, rd_I_n2056}), .b ({new_AGEMA_signal_4210, new_AGEMA_signal_4209, rd_I_n2055}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_4750, new_AGEMA_signal_4749, rd_I_n2057}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1276 ( .a ({new_AGEMA_signal_5510, new_AGEMA_signal_5509, rd_I_n2054}), .b ({new_AGEMA_signal_3768, new_AGEMA_signal_3767, rd_I_n2482}), .c ({state_out_s2[360], state_out_s1[360], state_out_s0[360]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1275 ( .a ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, rd_I_n2053}), .b ({new_AGEMA_signal_3770, new_AGEMA_signal_3769, rd_I_n2485}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_5510, new_AGEMA_signal_5509, rd_I_n2054}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1273 ( .a ({new_AGEMA_signal_3824, new_AGEMA_signal_3823, rd_I_n2172}), .b ({new_AGEMA_signal_4754, new_AGEMA_signal_4753, rd_I_n2052}), .c ({state_out_s2[44], state_out_s1[44], state_out_s0[44]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1272 ( .a ({new_AGEMA_signal_3826, new_AGEMA_signal_3825, rd_I_n2171}), .b ({new_AGEMA_signal_3822, new_AGEMA_signal_3821, rd_I_n2174}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_4754, new_AGEMA_signal_4753, rd_I_n2052}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1271 ( .a ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, rd_I_n2051}), .b ({new_AGEMA_signal_4146, new_AGEMA_signal_4145, rd_I_n2050}), .c ({state_out_s2[205], state_out_s1[205], state_out_s0[205]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1270 ( .a ({new_AGEMA_signal_4756, new_AGEMA_signal_4755, rd_I_n2049}), .b ({new_AGEMA_signal_4148, new_AGEMA_signal_4147, rd_I_n2048}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, rd_I_n2051}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1268 ( .a ({new_AGEMA_signal_3974, new_AGEMA_signal_3973, rd_I_n2506}), .b ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, rd_I_n2046}), .c ({state_out_s2[383], state_out_s1[383], state_out_s0[383]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1267 ( .a ({new_AGEMA_signal_3976, new_AGEMA_signal_3975, rd_I_n2505}), .b ({new_AGEMA_signal_3972, new_AGEMA_signal_3971, rd_I_n2508}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, rd_I_n2046}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1266 ( .a ({new_AGEMA_signal_3760, new_AGEMA_signal_3759, rd_I_n2606}), .b ({new_AGEMA_signal_4760, new_AGEMA_signal_4759, rd_I_n2045}), .c ({state_out_s2[19], state_out_s1[19], state_out_s0[19]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1265 ( .a ({new_AGEMA_signal_3758, new_AGEMA_signal_3757, rd_I_n2608}), .b ({new_AGEMA_signal_3756, new_AGEMA_signal_3755, rd_I_n2605}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_4760, new_AGEMA_signal_4759, rd_I_n2045}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1260 ( .a ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, rd_I_n2041}), .b ({new_AGEMA_signal_3762, new_AGEMA_signal_3761, rd_I_n2428}), .c ({state_out_s2[180], state_out_s1[180], state_out_s0[180]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1259 ( .a ({new_AGEMA_signal_4762, new_AGEMA_signal_4761, rd_I_n2040}), .b ({new_AGEMA_signal_3764, new_AGEMA_signal_3763, rd_I_n2431}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, rd_I_n2041}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1257 ( .a ({new_AGEMA_signal_4238, new_AGEMA_signal_4237, rd_I_n2552}), .b ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, rd_I_n2039}), .c ({state_out_s2[326], state_out_s1[326], state_out_s0[326]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1256 ( .a ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, rd_I_n2551}), .b ({new_AGEMA_signal_4236, new_AGEMA_signal_4235, rd_I_n2554}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_5522, new_AGEMA_signal_5521, rd_I_n2039}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1255 ( .a ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, rd_I_n2038}), .b ({new_AGEMA_signal_4012, new_AGEMA_signal_4011, rd_I_n2180}), .c ({state_out_s2[88], state_out_s1[88], state_out_s0[88]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1254 ( .a ({new_AGEMA_signal_4764, new_AGEMA_signal_4763, rd_I_n2037}), .b ({new_AGEMA_signal_4010, new_AGEMA_signal_4009, rd_I_n2183}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_5524, new_AGEMA_signal_5523, rd_I_n2038}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1252 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, rd_I_n2036}), .b ({new_AGEMA_signal_3850, new_AGEMA_signal_3849, rd_I_n2176}), .c ({state_out_s2[65], state_out_s1[65], state_out_s0[65]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1251 ( .a ({new_AGEMA_signal_4766, new_AGEMA_signal_4765, rd_I_n2035}), .b ({new_AGEMA_signal_3848, new_AGEMA_signal_3847, rd_I_n2179}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, rd_I_n2036}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1249 ( .a ({new_AGEMA_signal_3920, new_AGEMA_signal_3919, rd_I_n2303}), .b ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, rd_I_n2034}), .c ({state_out_s2[249], state_out_s1[249], state_out_s0[249]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1248 ( .a ({new_AGEMA_signal_3922, new_AGEMA_signal_3921, rd_I_n2302}), .b ({new_AGEMA_signal_3918, new_AGEMA_signal_3917, rd_I_n2305}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_4768, new_AGEMA_signal_4767, rd_I_n2034}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1247 ( .a ({new_AGEMA_signal_3884, new_AGEMA_signal_3883, rd_I_n2246}), .b ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, rd_I_n2033}), .c ({state_out_s2[226], state_out_s1[226], state_out_s0[226]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1246 ( .a ({new_AGEMA_signal_3886, new_AGEMA_signal_3885, rd_I_n2245}), .b ({new_AGEMA_signal_3882, new_AGEMA_signal_3881, rd_I_n2248}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, rd_I_n2033}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1245 ( .a ({new_AGEMA_signal_4148, new_AGEMA_signal_4147, rd_I_n2048}), .b ({new_AGEMA_signal_4772, new_AGEMA_signal_4771, rd_I_n2032}), .c ({state_out_s2[276], state_out_s1[276], state_out_s0[276]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1244 ( .a ({new_AGEMA_signal_4150, new_AGEMA_signal_4149, rd_I_n2047}), .b ({new_AGEMA_signal_4146, new_AGEMA_signal_4145, rd_I_n2050}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_4772, new_AGEMA_signal_4771, rd_I_n2032}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1243 ( .a ({new_AGEMA_signal_4168, new_AGEMA_signal_4167, rd_I_n2192}), .b ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, rd_I_n2031}), .c ({state_out_s2[267], state_out_s1[267], state_out_s0[267]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1242 ( .a ({new_AGEMA_signal_4164, new_AGEMA_signal_4163, rd_I_n2191}), .b ({new_AGEMA_signal_4166, new_AGEMA_signal_4165, rd_I_n2194}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_4774, new_AGEMA_signal_4773, rd_I_n2031}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1241 ( .a ({new_AGEMA_signal_3766, new_AGEMA_signal_3765, rd_I_n2429}), .b ({new_AGEMA_signal_4776, new_AGEMA_signal_4775, rd_I_n2030}), .c ({state_out_s2[51], state_out_s1[51], state_out_s0[51]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1240 ( .a ({new_AGEMA_signal_3764, new_AGEMA_signal_3763, rd_I_n2431}), .b ({new_AGEMA_signal_3762, new_AGEMA_signal_3761, rd_I_n2428}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_4776, new_AGEMA_signal_4775, rd_I_n2030}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1236 ( .a ({new_AGEMA_signal_4022, new_AGEMA_signal_4021, rd_I_n2028}), .b ({new_AGEMA_signal_4778, new_AGEMA_signal_4777, rd_I_n2027}), .c ({state_out_s2[212], state_out_s1[212], state_out_s0[212]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1235 ( .a ({new_AGEMA_signal_4024, new_AGEMA_signal_4023, rd_I_n2026}), .b ({new_AGEMA_signal_4020, new_AGEMA_signal_4019, rd_I_n2025}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_4778, new_AGEMA_signal_4777, rd_I_n2027}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1234 ( .a ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, rd_I_n2024}), .b ({new_AGEMA_signal_4246, new_AGEMA_signal_4245, rd_I_n2423}), .c ({state_out_s2[358], state_out_s1[358], state_out_s0[358]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1233 ( .a ({new_AGEMA_signal_4780, new_AGEMA_signal_4779, rd_I_n2023}), .b ({new_AGEMA_signal_4244, new_AGEMA_signal_4243, rd_I_n2426}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_5540, new_AGEMA_signal_5539, rd_I_n2024}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1231 ( .a ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, rd_I_n2022}), .b ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, rd_I_n2021}), .c ({state_out_s2[0], state_out_s1[0], state_out_s0[0]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1230 ( .a ({new_AGEMA_signal_4782, new_AGEMA_signal_4781, rd_I_n2020}), .b ({new_AGEMA_signal_3866, new_AGEMA_signal_3865, rd_I_n2019}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_5542, new_AGEMA_signal_5541, rd_I_n2022}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1228 ( .a ({new_AGEMA_signal_3772, new_AGEMA_signal_3771, rd_I_n2483}), .b ({new_AGEMA_signal_4784, new_AGEMA_signal_4783, rd_I_n2017}), .c ({state_out_s2[161], state_out_s1[161], state_out_s0[161]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1227 ( .a ({new_AGEMA_signal_3770, new_AGEMA_signal_3769, rd_I_n2485}), .b ({new_AGEMA_signal_3768, new_AGEMA_signal_3767, rd_I_n2482}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_4784, new_AGEMA_signal_4783, rd_I_n2017}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1223 ( .a ({new_AGEMA_signal_5546, new_AGEMA_signal_5545, rd_I_n2014}), .b ({new_AGEMA_signal_4060, new_AGEMA_signal_4059, rd_I_n2579}), .c ({state_out_s2[339], state_out_s1[339], state_out_s0[339]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1222 ( .a ({new_AGEMA_signal_4786, new_AGEMA_signal_4785, rd_I_n2013}), .b ({new_AGEMA_signal_5042, new_AGEMA_signal_5041, rd_I_n2582}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_5546, new_AGEMA_signal_5545, rd_I_n2014}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1220 ( .a ({new_AGEMA_signal_3778, new_AGEMA_signal_3777, rd_I_n2530}), .b ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, rd_I_n2012}), .c ({state_out_s2[42], state_out_s1[42], state_out_s0[42]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1219 ( .a ({new_AGEMA_signal_3776, new_AGEMA_signal_3775, rd_I_n2531}), .b ({new_AGEMA_signal_3774, new_AGEMA_signal_3773, rd_I_n2533}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, rd_I_n2012}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1215 ( .a ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, rd_I_n2009}), .b ({new_AGEMA_signal_4198, new_AGEMA_signal_4197, rd_I_n2008}), .c ({state_out_s2[203], state_out_s1[203], state_out_s0[203]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1214 ( .a ({new_AGEMA_signal_4790, new_AGEMA_signal_4789, rd_I_n2007}), .b ({new_AGEMA_signal_4196, new_AGEMA_signal_4195, rd_I_n2006}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, rd_I_n2009}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1212 ( .a ({new_AGEMA_signal_5552, new_AGEMA_signal_5551, rd_I_n2004}), .b ({new_AGEMA_signal_3858, new_AGEMA_signal_3857, rd_I_n2059}), .c ({state_out_s2[381], state_out_s1[381], state_out_s0[381]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1211 ( .a ({new_AGEMA_signal_4792, new_AGEMA_signal_4791, rd_I_n2003}), .b ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, rd_I_n2062}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_5552, new_AGEMA_signal_5551, rd_I_n2004}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1209 ( .a ({new_AGEMA_signal_5554, new_AGEMA_signal_5553, rd_I_n2002}), .b ({new_AGEMA_signal_4374, new_AGEMA_signal_4373, rd_I_n2001}), .c ({state_out_s2[26], state_out_s1[26], state_out_s0[26]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1208 ( .a ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, rd_I_n2000}), .b ({new_AGEMA_signal_4376, new_AGEMA_signal_4375, rd_I_n1999}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_5554, new_AGEMA_signal_5553, rd_I_n2002}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1206 ( .a ({new_AGEMA_signal_3932, new_AGEMA_signal_3931, rd_I_n2206}), .b ({new_AGEMA_signal_4796, new_AGEMA_signal_4795, rd_I_n1997}), .c ({state_out_s2[187], state_out_s1[187], state_out_s0[187]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1205 ( .a ({new_AGEMA_signal_3934, new_AGEMA_signal_3933, rd_I_n2205}), .b ({new_AGEMA_signal_3930, new_AGEMA_signal_3929, rd_I_n2208}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_4796, new_AGEMA_signal_4795, rd_I_n1997}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1204 ( .a ({new_AGEMA_signal_4436, new_AGEMA_signal_4435, rd_I_n2255}), .b ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, rd_I_n1996}), .c ({state_out_s2[333], state_out_s1[333], state_out_s0[333]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1203 ( .a ({new_AGEMA_signal_4438, new_AGEMA_signal_4437, rd_I_n2254}), .b ({new_AGEMA_signal_4434, new_AGEMA_signal_4433, rd_I_n2257}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_4798, new_AGEMA_signal_4797, rd_I_n1996}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1202 ( .a ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, rd_I_n1995}), .b ({new_AGEMA_signal_4392, new_AGEMA_signal_4391, rd_I_n1994}), .c ({state_out_s2[29], state_out_s1[29], state_out_s0[29]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1201 ( .a ({new_AGEMA_signal_4800, new_AGEMA_signal_4799, rd_I_n1993}), .b ({new_AGEMA_signal_4394, new_AGEMA_signal_4393, rd_I_n1992}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_5560, new_AGEMA_signal_5559, rd_I_n1995}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1199 ( .a ({new_AGEMA_signal_3784, new_AGEMA_signal_3783, rd_I_n2372}), .b ({new_AGEMA_signal_4802, new_AGEMA_signal_4801, rd_I_n1990}), .c ({state_out_s2[190], state_out_s1[190], state_out_s0[190]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1198 ( .a ({new_AGEMA_signal_3782, new_AGEMA_signal_3781, rd_I_n2374}), .b ({new_AGEMA_signal_3780, new_AGEMA_signal_3779, rd_I_n2371}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_4802, new_AGEMA_signal_4801, rd_I_n1990}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1194 ( .a ({new_AGEMA_signal_5564, new_AGEMA_signal_5563, rd_I_n1987}), .b ({new_AGEMA_signal_4284, new_AGEMA_signal_4283, rd_I_n2617}), .c ({state_out_s2[336], state_out_s1[336], state_out_s0[336]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1193 ( .a ({new_AGEMA_signal_4804, new_AGEMA_signal_4803, rd_I_n1986}), .b ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, rd_I_n2620}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_5564, new_AGEMA_signal_5563, rd_I_n1987}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1191 ( .a ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, rd_I_n1985}), .b ({new_AGEMA_signal_3948, new_AGEMA_signal_3947, rd_I_n1984}), .c ({state_out_s2[119], state_out_s1[119], state_out_s0[119]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1190 ( .a ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, rd_I_n1983}), .b ({new_AGEMA_signal_3950, new_AGEMA_signal_3949, rd_I_n1982}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_5566, new_AGEMA_signal_5565, rd_I_n1985}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1188 ( .a ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, rd_I_n1980}), .b ({new_AGEMA_signal_4358, new_AGEMA_signal_4357, rd_I_n1979}), .c ({state_out_s2[110], state_out_s1[110], state_out_s0[110]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1187 ( .a ({new_AGEMA_signal_4360, new_AGEMA_signal_4359, rd_I_n1978}), .b ({new_AGEMA_signal_4808, new_AGEMA_signal_4807, rd_I_n1977}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, rd_I_n1980}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1185 ( .a ({new_AGEMA_signal_3836, new_AGEMA_signal_3835, rd_I_n2516}), .b ({new_AGEMA_signal_5570, new_AGEMA_signal_5569, rd_I_n1975}), .c ({state_out_s2[152], state_out_s1[152], state_out_s0[152]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1184 ( .a ({new_AGEMA_signal_3834, new_AGEMA_signal_3833, rd_I_n2515}), .b ({new_AGEMA_signal_4856, new_AGEMA_signal_4855, rd_I_n2518}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_5570, new_AGEMA_signal_5569, rd_I_n1975}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1183 ( .a ({new_AGEMA_signal_3842, new_AGEMA_signal_3841, rd_I_n2511}), .b ({new_AGEMA_signal_5572, new_AGEMA_signal_5571, rd_I_n1974}), .c ({state_out_s2[143], state_out_s1[143], state_out_s0[143]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1182 ( .a ({new_AGEMA_signal_3840, new_AGEMA_signal_3839, rd_I_n2510}), .b ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, rd_I_n2513}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_5572, new_AGEMA_signal_5571, rd_I_n1974}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1181 ( .a ({new_AGEMA_signal_4400, new_AGEMA_signal_4399, rd_I_n2113}), .b ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, rd_I_n1973}), .c ({state_out_s2[298], state_out_s1[298], state_out_s0[298]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1180 ( .a ({new_AGEMA_signal_4398, new_AGEMA_signal_4397, rd_I_n2112}), .b ({new_AGEMA_signal_4402, new_AGEMA_signal_4401, rd_I_n2115}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_4810, new_AGEMA_signal_4809, rd_I_n1973}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1179 ( .a ({new_AGEMA_signal_4418, new_AGEMA_signal_4417, rd_I_n2221}), .b ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, rd_I_n1972}), .c ({state_out_s2[289], state_out_s1[289], state_out_s0[289]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1178 ( .a ({new_AGEMA_signal_4416, new_AGEMA_signal_4415, rd_I_n2220}), .b ({new_AGEMA_signal_4420, new_AGEMA_signal_4419, rd_I_n2223}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, rd_I_n1972}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1177 ( .a ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, rd_I_n1971}), .b ({new_AGEMA_signal_3982, new_AGEMA_signal_3981, rd_I_n1970}), .c ({state_out_s2[34], state_out_s1[34], state_out_s0[34]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1176 ( .a ({new_AGEMA_signal_4814, new_AGEMA_signal_4813, rd_I_n1969}), .b ({new_AGEMA_signal_3980, new_AGEMA_signal_3979, rd_I_n1968}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_5578, new_AGEMA_signal_5577, rd_I_n1971}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1174 ( .a ({new_AGEMA_signal_3794, new_AGEMA_signal_3793, rd_I_n2118}), .b ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, rd_I_n1966}), .c ({state_out_s2[195], state_out_s1[195], state_out_s0[195]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1173 ( .a ({new_AGEMA_signal_3796, new_AGEMA_signal_3795, rd_I_n2117}), .b ({new_AGEMA_signal_3792, new_AGEMA_signal_3791, rd_I_n2120}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_4816, new_AGEMA_signal_4815, rd_I_n1966}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1172 ( .a ({new_AGEMA_signal_3790, new_AGEMA_signal_3789, rd_I_n2149}), .b ({new_AGEMA_signal_4818, new_AGEMA_signal_4817, rd_I_n1965}), .c ({state_out_s2[373], state_out_s1[373], state_out_s0[373]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1171 ( .a ({new_AGEMA_signal_3788, new_AGEMA_signal_3787, rd_I_n2151}), .b ({new_AGEMA_signal_3786, new_AGEMA_signal_3785, rd_I_n2148}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_4818, new_AGEMA_signal_4817, rd_I_n1965}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1167 ( .a ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, rd_I_n1963}), .b ({new_AGEMA_signal_4162, new_AGEMA_signal_4161, rd_I_n1962}), .c ({state_out_s2[87], state_out_s1[87], state_out_s0[87]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1166 ( .a ({new_AGEMA_signal_4820, new_AGEMA_signal_4819, rd_I_n1961}), .b ({new_AGEMA_signal_4160, new_AGEMA_signal_4159, rd_I_n1960}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_5584, new_AGEMA_signal_5583, rd_I_n1963}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1164 ( .a ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, rd_I_n1958}), .b ({new_AGEMA_signal_3898, new_AGEMA_signal_3897, rd_I_n2473}), .c ({state_out_s2[64], state_out_s1[64], state_out_s0[64]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1163 ( .a ({new_AGEMA_signal_4822, new_AGEMA_signal_4821, rd_I_n1957}), .b ({new_AGEMA_signal_3896, new_AGEMA_signal_3895, rd_I_n2476}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, rd_I_n1958}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1161 ( .a ({new_AGEMA_signal_3950, new_AGEMA_signal_3949, rd_I_n1982}), .b ({new_AGEMA_signal_4824, new_AGEMA_signal_4823, rd_I_n1956}), .c ({state_out_s2[248], state_out_s1[248], state_out_s0[248]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1160 ( .a ({new_AGEMA_signal_3952, new_AGEMA_signal_3951, rd_I_n1981}), .b ({new_AGEMA_signal_3948, new_AGEMA_signal_3947, rd_I_n1984}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_4824, new_AGEMA_signal_4823, rd_I_n1956}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1159 ( .a ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, rd_I_n1955}), .b ({new_AGEMA_signal_3798, new_AGEMA_signal_3797, rd_I_n2537}), .c ({state_out_s2[225], state_out_s1[225], state_out_s0[225]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1158 ( .a ({new_AGEMA_signal_4826, new_AGEMA_signal_4825, rd_I_n1954}), .b ({new_AGEMA_signal_3800, new_AGEMA_signal_3799, rd_I_n2540}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, rd_I_n1955}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1156 ( .a ({new_AGEMA_signal_4178, new_AGEMA_signal_4177, rd_I_n2088}), .b ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, rd_I_n1953}), .c ({state_out_s2[275], state_out_s1[275], state_out_s0[275]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1155 ( .a ({new_AGEMA_signal_4176, new_AGEMA_signal_4175, rd_I_n2087}), .b ({new_AGEMA_signal_4180, new_AGEMA_signal_4179, rd_I_n2090}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({new_AGEMA_signal_4828, new_AGEMA_signal_4827, rd_I_n1953}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1154 ( .a ({new_AGEMA_signal_3796, new_AGEMA_signal_3795, rd_I_n2117}), .b ({new_AGEMA_signal_4830, new_AGEMA_signal_4829, rd_I_n1952}), .c ({state_out_s2[266], state_out_s1[266], state_out_s0[266]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1153 ( .a ({new_AGEMA_signal_3794, new_AGEMA_signal_3793, rd_I_n2118}), .b ({new_AGEMA_signal_3792, new_AGEMA_signal_3791, rd_I_n2120}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_4830, new_AGEMA_signal_4829, rd_I_n1952}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1149 ( .a ({new_AGEMA_signal_3802, new_AGEMA_signal_3801, rd_I_n2538}), .b ({new_AGEMA_signal_4832, new_AGEMA_signal_4831, rd_I_n1949}), .c ({state_out_s2[96], state_out_s1[96], state_out_s0[96]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1148 ( .a ({new_AGEMA_signal_3800, new_AGEMA_signal_3799, rd_I_n2540}), .b ({new_AGEMA_signal_3798, new_AGEMA_signal_3797, rd_I_n2537}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({new_AGEMA_signal_4832, new_AGEMA_signal_4831, rd_I_n1949}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1144 ( .a ({new_AGEMA_signal_3866, new_AGEMA_signal_3865, rd_I_n2019}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, rd_I_n1945}), .c ({state_out_s2[129], state_out_s1[129], state_out_s0[129]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1143 ( .a ({new_AGEMA_signal_3868, new_AGEMA_signal_3867, rd_I_n2018}), .b ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, rd_I_n2021}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, rd_I_n1945}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1142 ( .a ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, rd_I_n1944}), .b ({new_AGEMA_signal_4182, new_AGEMA_signal_4181, rd_I_n1943}), .c ({state_out_s2[307], state_out_s1[307], state_out_s0[307]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1141 ( .a ({new_AGEMA_signal_4834, new_AGEMA_signal_4833, rd_I_n1942}), .b ({new_AGEMA_signal_4184, new_AGEMA_signal_4183, rd_I_n1941}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({new_AGEMA_signal_5600, new_AGEMA_signal_5599, rd_I_n1944}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1139 ( .a ({new_AGEMA_signal_3808, new_AGEMA_signal_3807, rd_I_n2338}), .b ({new_AGEMA_signal_4836, new_AGEMA_signal_4835, rd_I_n1939}), .c ({state_out_s2[28], state_out_s1[28], state_out_s0[28]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1138 ( .a ({new_AGEMA_signal_3806, new_AGEMA_signal_3805, rd_I_n2339}), .b ({new_AGEMA_signal_3804, new_AGEMA_signal_3803, rd_I_n2341}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_4836, new_AGEMA_signal_4835, rd_I_n1939}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1133 ( .a ({new_AGEMA_signal_3818, new_AGEMA_signal_3817, rd_I_n2328}), .b ({new_AGEMA_signal_4838, new_AGEMA_signal_4837, rd_I_n1934}), .c ({state_out_s2[189], state_out_s1[189], state_out_s0[189]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1132 ( .a ({new_AGEMA_signal_3820, new_AGEMA_signal_3819, rd_I_n2327}), .b ({new_AGEMA_signal_3816, new_AGEMA_signal_3815, rd_I_n2330}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({new_AGEMA_signal_4838, new_AGEMA_signal_4837, rd_I_n1934}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1131 ( .a ({new_AGEMA_signal_4106, new_AGEMA_signal_4105, rd_I_n2395}), .b ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, rd_I_n1933}), .c ({state_out_s2[335], state_out_s1[335], state_out_s0[335]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1130 ( .a ({new_AGEMA_signal_4108, new_AGEMA_signal_4107, rd_I_n2394}), .b ({new_AGEMA_signal_4104, new_AGEMA_signal_4103, rd_I_n2397}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_4840, new_AGEMA_signal_4839, rd_I_n1933}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1129 ( .a ({new_AGEMA_signal_3814, new_AGEMA_signal_3813, rd_I_n2358}), .b ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, rd_I_n1932}), .c ({state_out_s2[49], state_out_s1[49], state_out_s0[49]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1128 ( .a ({new_AGEMA_signal_3812, new_AGEMA_signal_3811, rd_I_n2360}), .b ({new_AGEMA_signal_3810, new_AGEMA_signal_3809, rd_I_n2357}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, rd_I_n1932}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1124 ( .a ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, rd_I_n1930}), .b ({new_AGEMA_signal_4042, new_AGEMA_signal_4041, rd_I_n2064}), .c ({state_out_s2[210], state_out_s1[210], state_out_s0[210]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1123 ( .a ({new_AGEMA_signal_4844, new_AGEMA_signal_4843, rd_I_n1929}), .b ({new_AGEMA_signal_4040, new_AGEMA_signal_4039, rd_I_n2067}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, rd_I_n1930}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1121 ( .a ({new_AGEMA_signal_3820, new_AGEMA_signal_3819, rd_I_n2327}), .b ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, rd_I_n1928}), .c ({state_out_s2[356], state_out_s1[356], state_out_s0[356]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1120 ( .a ({new_AGEMA_signal_3818, new_AGEMA_signal_3817, rd_I_n2328}), .b ({new_AGEMA_signal_3816, new_AGEMA_signal_3815, rd_I_n2330}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({new_AGEMA_signal_4846, new_AGEMA_signal_4845, rd_I_n1928}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1116 ( .a ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, rd_I_n2521}), .b ({new_AGEMA_signal_4848, new_AGEMA_signal_4847, rd_I_n1926}), .c ({state_out_s2[12], state_out_s1[12], state_out_s0[12]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1115 ( .a ({new_AGEMA_signal_3942, new_AGEMA_signal_3941, rd_I_n2520}), .b ({new_AGEMA_signal_3946, new_AGEMA_signal_3945, rd_I_n2523}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_4848, new_AGEMA_signal_4847, rd_I_n1926}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1114 ( .a ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, rd_I_n2376}), .b ({new_AGEMA_signal_4850, new_AGEMA_signal_4849, rd_I_n1925}), .c ({state_out_s2[3], state_out_s1[3], state_out_s0[3]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1113 ( .a ({new_AGEMA_signal_4354, new_AGEMA_signal_4353, rd_I_n2375}), .b ({new_AGEMA_signal_4350, new_AGEMA_signal_4349, rd_I_n2378}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({new_AGEMA_signal_4850, new_AGEMA_signal_4849, rd_I_n1925}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1112 ( .a ({new_AGEMA_signal_3826, new_AGEMA_signal_3825, rd_I_n2171}), .b ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, rd_I_n1924}), .c ({state_out_s2[173], state_out_s1[173], state_out_s0[173]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1111 ( .a ({new_AGEMA_signal_3824, new_AGEMA_signal_3823, rd_I_n2172}), .b ({new_AGEMA_signal_3822, new_AGEMA_signal_3821, rd_I_n2174}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_4852, new_AGEMA_signal_4851, rd_I_n1924}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1107 ( .a ({new_AGEMA_signal_3832, new_AGEMA_signal_3831, rd_I_n2202}), .b ({new_AGEMA_signal_4854, new_AGEMA_signal_4853, rd_I_n1921}), .c ({state_out_s2[164], state_out_s1[164], state_out_s0[164]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1106 ( .a ({new_AGEMA_signal_3830, new_AGEMA_signal_3829, rd_I_n2204}), .b ({new_AGEMA_signal_3828, new_AGEMA_signal_3827, rd_I_n2201}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({new_AGEMA_signal_4854, new_AGEMA_signal_4853, rd_I_n1921}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1102 ( .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, rd_I_n1918}), .b ({new_AGEMA_signal_3834, new_AGEMA_signal_3833, rd_I_n2515}), .c ({state_out_s2[351], state_out_s1[351], state_out_s0[351]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1100 ( .a ({new_AGEMA_signal_4856, new_AGEMA_signal_4855, rd_I_n2518}), .b ({new_AGEMA_signal_3836, new_AGEMA_signal_3835, rd_I_n2516}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, rd_I_n1918}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1096 ( .a ({new_AGEMA_signal_5624, new_AGEMA_signal_5623, rd_I_n1914}), .b ({new_AGEMA_signal_3840, new_AGEMA_signal_3839, rd_I_n2510}), .c ({state_out_s2[342], state_out_s1[342], state_out_s0[342]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1094 ( .a ({new_AGEMA_signal_4858, new_AGEMA_signal_4857, rd_I_n2513}), .b ({new_AGEMA_signal_3842, new_AGEMA_signal_3841, rd_I_n2511}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({new_AGEMA_signal_5624, new_AGEMA_signal_5623, rd_I_n1914}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1090 ( .a ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, rd_I_n1910}), .b ({new_AGEMA_signal_3928, new_AGEMA_signal_3927, rd_I_n2432}), .c ({state_out_s2[95], state_out_s1[95], state_out_s0[95]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1089 ( .a ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, rd_I_n1909}), .b ({new_AGEMA_signal_3926, new_AGEMA_signal_3925, rd_I_n2435}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, rd_I_n1910}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1087 ( .a ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, rd_I_n1908}), .b ({new_AGEMA_signal_4192, new_AGEMA_signal_4191, rd_I_n2135}), .c ({state_out_s2[86], state_out_s1[86], state_out_s0[86]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1086 ( .a ({new_AGEMA_signal_4862, new_AGEMA_signal_4861, rd_I_n1907}), .b ({new_AGEMA_signal_4190, new_AGEMA_signal_4189, rd_I_n2138}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, rd_I_n1908}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1084 ( .a ({new_AGEMA_signal_4064, new_AGEMA_signal_4063, rd_I_n1906}), .b ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, rd_I_n1905}), .c ({state_out_s2[247], state_out_s1[247], state_out_s0[247]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1083 ( .a ({new_AGEMA_signal_4062, new_AGEMA_signal_4061, rd_I_n1904}), .b ({new_AGEMA_signal_4066, new_AGEMA_signal_4065, rd_I_n1903}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_4864, new_AGEMA_signal_4863, rd_I_n1905}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1082 ( .a ({new_AGEMA_signal_4070, new_AGEMA_signal_4069, rd_I_n1902}), .b ({new_AGEMA_signal_4866, new_AGEMA_signal_4865, rd_I_n1901}), .c ({state_out_s2[224], state_out_s1[224], state_out_s0[224]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1081 ( .a ({new_AGEMA_signal_4072, new_AGEMA_signal_4071, rd_I_n1900}), .b ({new_AGEMA_signal_4068, new_AGEMA_signal_4067, rd_I_n1899}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({new_AGEMA_signal_4866, new_AGEMA_signal_4865, rd_I_n1901}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1080 ( .a ({new_AGEMA_signal_4196, new_AGEMA_signal_4195, rd_I_n2006}), .b ({new_AGEMA_signal_4868, new_AGEMA_signal_4867, rd_I_n1898}), .c ({state_out_s2[274], state_out_s1[274], state_out_s0[274]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1079 ( .a ({new_AGEMA_signal_4194, new_AGEMA_signal_4193, rd_I_n2005}), .b ({new_AGEMA_signal_4198, new_AGEMA_signal_4197, rd_I_n2008}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_4868, new_AGEMA_signal_4867, rd_I_n1898}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1078 ( .a ({new_AGEMA_signal_4870, new_AGEMA_signal_4869, rd_I_n1897}), .b ({new_AGEMA_signal_3846, new_AGEMA_signal_3845, rd_I_n2177}), .c ({state_out_s2[265], state_out_s1[265], state_out_s0[265]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1076 ( .a ({new_AGEMA_signal_3850, new_AGEMA_signal_3849, rd_I_n2176}), .b ({new_AGEMA_signal_3848, new_AGEMA_signal_3847, rd_I_n2179}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({new_AGEMA_signal_4870, new_AGEMA_signal_4869, rd_I_n1897}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1072 ( .a ({new_AGEMA_signal_3856, new_AGEMA_signal_3855, rd_I_n2546}), .b ({new_AGEMA_signal_4872, new_AGEMA_signal_4871, rd_I_n1892}), .c ({state_out_s2[21], state_out_s1[21], state_out_s0[21]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1071 ( .a ({new_AGEMA_signal_3854, new_AGEMA_signal_3853, rd_I_n2547}), .b ({new_AGEMA_signal_3852, new_AGEMA_signal_3851, rd_I_n2549}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_4872, new_AGEMA_signal_4871, rd_I_n1892}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1066 ( .a ({new_AGEMA_signal_3862, new_AGEMA_signal_3861, rd_I_n2060}), .b ({new_AGEMA_signal_4874, new_AGEMA_signal_4873, rd_I_n1889}), .c ({state_out_s2[182], state_out_s1[182], state_out_s0[182]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1065 ( .a ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, rd_I_n2062}), .b ({new_AGEMA_signal_3858, new_AGEMA_signal_3857, rd_I_n2059}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({new_AGEMA_signal_4874, new_AGEMA_signal_4873, rd_I_n1889}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1061 ( .a ({new_AGEMA_signal_3868, new_AGEMA_signal_3867, rd_I_n2018}), .b ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, rd_I_n1888}), .c ({state_out_s2[328], state_out_s1[328], state_out_s0[328]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1060 ( .a ({new_AGEMA_signal_3866, new_AGEMA_signal_3865, rd_I_n2019}), .b ({new_AGEMA_signal_4876, new_AGEMA_signal_4875, rd_I_n2021}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_5642, new_AGEMA_signal_5641, rd_I_n1888}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1054 ( .a ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, rd_I_n1884}), .b ({new_AGEMA_signal_4068, new_AGEMA_signal_4067, rd_I_n1899}), .c ({state_out_s2[127], state_out_s1[127], state_out_s0[127]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1053 ( .a ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, rd_I_n1883}), .b ({new_AGEMA_signal_4070, new_AGEMA_signal_4069, rd_I_n1902}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, rd_I_n1884}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1051 ( .a ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, rd_I_n1882}), .b ({new_AGEMA_signal_4066, new_AGEMA_signal_4065, rd_I_n1903}), .c ({state_out_s2[118], state_out_s1[118], state_out_s0[118]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1050 ( .a ({new_AGEMA_signal_4880, new_AGEMA_signal_4879, rd_I_n1881}), .b ({new_AGEMA_signal_4064, new_AGEMA_signal_4063, rd_I_n1906}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, rd_I_n1882}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1048 ( .a ({new_AGEMA_signal_3874, new_AGEMA_signal_3873, rd_I_n2597}), .b ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, rd_I_n1880}), .c ({state_out_s2[151], state_out_s1[151], state_out_s0[151]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1047 ( .a ({new_AGEMA_signal_4882, new_AGEMA_signal_4881, rd_I_n2599}), .b ({new_AGEMA_signal_3870, new_AGEMA_signal_3869, rd_I_n2596}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({new_AGEMA_signal_5648, new_AGEMA_signal_5647, rd_I_n1880}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1041 ( .a ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, rd_I_n1875}), .b ({new_AGEMA_signal_3876, new_AGEMA_signal_3875, rd_I_n2622}), .c ({state_out_s2[128], state_out_s1[128], state_out_s0[128]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1039 ( .a ({new_AGEMA_signal_3880, new_AGEMA_signal_3879, rd_I_n2621}), .b ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, rd_I_n2624}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, rd_I_n1875}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1035 ( .a ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, rd_I_n1872}), .b ({new_AGEMA_signal_4204, new_AGEMA_signal_4203, rd_I_n1871}), .c ({state_out_s2[306], state_out_s1[306], state_out_s0[306]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1034 ( .a ({new_AGEMA_signal_4886, new_AGEMA_signal_4885, rd_I_n1870}), .b ({new_AGEMA_signal_4202, new_AGEMA_signal_4201, rd_I_n1869}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, rd_I_n1872}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1032 ( .a ({new_AGEMA_signal_3886, new_AGEMA_signal_3885, rd_I_n2245}), .b ({new_AGEMA_signal_4888, new_AGEMA_signal_4887, rd_I_n1867}), .c ({state_out_s2[297], state_out_s1[297], state_out_s0[297]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1031 ( .a ({new_AGEMA_signal_3884, new_AGEMA_signal_3883, rd_I_n2246}), .b ({new_AGEMA_signal_3882, new_AGEMA_signal_3881, rd_I_n2248}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_4888, new_AGEMA_signal_4887, rd_I_n1867}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1027 ( .a ({new_AGEMA_signal_5656, new_AGEMA_signal_5655, rd_I_n1866}), .b ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, rd_I_n1865}), .c ({state_out_s2[27], state_out_s1[27], state_out_s0[27]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1026 ( .a ({new_AGEMA_signal_4890, new_AGEMA_signal_4889, rd_I_n1864}), .b ({new_AGEMA_signal_4094, new_AGEMA_signal_4093, rd_I_n1863}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({new_AGEMA_signal_5656, new_AGEMA_signal_5655, rd_I_n1866}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1024 ( .a ({new_AGEMA_signal_3908, new_AGEMA_signal_3907, rd_I_n2279}), .b ({new_AGEMA_signal_4892, new_AGEMA_signal_4891, rd_I_n1861}), .c ({state_out_s2[188], state_out_s1[188], state_out_s0[188]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1023 ( .a ({new_AGEMA_signal_3910, new_AGEMA_signal_3909, rd_I_n2278}), .b ({new_AGEMA_signal_3906, new_AGEMA_signal_3905, rd_I_n2281}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_4892, new_AGEMA_signal_4891, rd_I_n1861}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1022 ( .a ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, rd_I_n1860}), .b ({new_AGEMA_signal_4324, new_AGEMA_signal_4323, rd_I_n1859}), .c ({state_out_s2[334], state_out_s1[334], state_out_s0[334]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1021 ( .a ({new_AGEMA_signal_4894, new_AGEMA_signal_4893, rd_I_n1858}), .b ({new_AGEMA_signal_5160, new_AGEMA_signal_5159, rd_I_n1857}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({new_AGEMA_signal_5660, new_AGEMA_signal_5659, rd_I_n1860}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1019 ( .a ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, rd_I_n1855}), .b ({new_AGEMA_signal_3960, new_AGEMA_signal_3959, rd_I_n2415}), .c ({state_out_s2[94], state_out_s1[94], state_out_s0[94]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1018 ( .a ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, rd_I_n1854}), .b ({new_AGEMA_signal_3962, new_AGEMA_signal_3961, rd_I_n2418}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, rd_I_n1855}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1016 ( .a ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, rd_I_n1853}), .b ({new_AGEMA_signal_4210, new_AGEMA_signal_4209, rd_I_n2055}), .c ({state_out_s2[85], state_out_s1[85], state_out_s0[85]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1015 ( .a ({new_AGEMA_signal_4898, new_AGEMA_signal_4897, rd_I_n1852}), .b ({new_AGEMA_signal_4208, new_AGEMA_signal_4207, rd_I_n2058}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, rd_I_n1853}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1013 ( .a ({new_AGEMA_signal_3892, new_AGEMA_signal_3891, rd_I_n2562}), .b ({new_AGEMA_signal_4900, new_AGEMA_signal_4899, rd_I_n1851}), .c ({state_out_s2[255], state_out_s1[255], state_out_s0[255]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1012 ( .a ({new_AGEMA_signal_3890, new_AGEMA_signal_3889, rd_I_n2564}), .b ({new_AGEMA_signal_3888, new_AGEMA_signal_3887, rd_I_n2561}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_4900, new_AGEMA_signal_4899, rd_I_n1851}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1008 ( .a ({new_AGEMA_signal_4124, new_AGEMA_signal_4123, rd_I_n2557}), .b ({new_AGEMA_signal_4902, new_AGEMA_signal_4901, rd_I_n1848}), .c ({state_out_s2[246], state_out_s1[246], state_out_s0[246]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1007 ( .a ({new_AGEMA_signal_4122, new_AGEMA_signal_4121, rd_I_n2556}), .b ({new_AGEMA_signal_4126, new_AGEMA_signal_4125, rd_I_n2559}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({new_AGEMA_signal_4902, new_AGEMA_signal_4901, rd_I_n1848}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1006 ( .a ({new_AGEMA_signal_4222, new_AGEMA_signal_4221, rd_I_n2478}), .b ({new_AGEMA_signal_4904, new_AGEMA_signal_4903, rd_I_n1847}), .c ({state_out_s2[273], state_out_s1[273], state_out_s0[273]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1005 ( .a ({new_AGEMA_signal_4218, new_AGEMA_signal_4217, rd_I_n2477}), .b ({new_AGEMA_signal_4220, new_AGEMA_signal_4219, rd_I_n2480}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_4904, new_AGEMA_signal_4903, rd_I_n1847}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1004 ( .a ({new_AGEMA_signal_4906, new_AGEMA_signal_4905, rd_I_n1846}), .b ({new_AGEMA_signal_3894, new_AGEMA_signal_3893, rd_I_n2474}), .c ({state_out_s2[264], state_out_s1[264], state_out_s0[264]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U1002 ( .a ({new_AGEMA_signal_3898, new_AGEMA_signal_3897, rd_I_n2473}), .b ({new_AGEMA_signal_3896, new_AGEMA_signal_3895, rd_I_n2476}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({new_AGEMA_signal_4906, new_AGEMA_signal_4905, rd_I_n1846}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U998 ( .a ({new_AGEMA_signal_4076, new_AGEMA_signal_4075, rd_I_n1842}), .b ({new_AGEMA_signal_4908, new_AGEMA_signal_4907, rd_I_n1841}), .c ({state_out_s2[57], state_out_s1[57], state_out_s0[57]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U997 ( .a ({new_AGEMA_signal_4078, new_AGEMA_signal_4077, rd_I_n1840}), .b ({new_AGEMA_signal_4074, new_AGEMA_signal_4073, rd_I_n1839}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_4908, new_AGEMA_signal_4907, rd_I_n1841}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U996 ( .a ({new_AGEMA_signal_4082, new_AGEMA_signal_4081, rd_I_n2310}), .b ({new_AGEMA_signal_4910, new_AGEMA_signal_4909, rd_I_n1838}), .c ({state_out_s2[48], state_out_s1[48], state_out_s0[48]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U995 ( .a ({new_AGEMA_signal_4084, new_AGEMA_signal_4083, rd_I_n2309}), .b ({new_AGEMA_signal_4080, new_AGEMA_signal_4079, rd_I_n2312}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({new_AGEMA_signal_4910, new_AGEMA_signal_4909, rd_I_n1838}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U994 ( .a ({new_AGEMA_signal_4100, new_AGEMA_signal_4099, rd_I_n2231}), .b ({new_AGEMA_signal_4912, new_AGEMA_signal_4911, rd_I_n1837}), .c ({state_out_s2[218], state_out_s1[218], state_out_s0[218]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U993 ( .a ({new_AGEMA_signal_4098, new_AGEMA_signal_4097, rd_I_n2230}), .b ({new_AGEMA_signal_4102, new_AGEMA_signal_4101, rd_I_n2233}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_4912, new_AGEMA_signal_4911, rd_I_n1837}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U992 ( .a ({new_AGEMA_signal_4268, new_AGEMA_signal_4267, rd_I_n2226}), .b ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, rd_I_n1836}), .c ({state_out_s2[209], state_out_s1[209], state_out_s0[209]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U991 ( .a ({new_AGEMA_signal_4266, new_AGEMA_signal_4265, rd_I_n2225}), .b ({new_AGEMA_signal_4270, new_AGEMA_signal_4269, rd_I_n2228}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, rd_I_n1836}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U990 ( .a ({new_AGEMA_signal_3904, new_AGEMA_signal_3903, rd_I_n2273}), .b ({new_AGEMA_signal_4916, new_AGEMA_signal_4915, rd_I_n1835}), .c ({state_out_s2[364], state_out_s1[364], state_out_s0[364]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U989 ( .a ({new_AGEMA_signal_3902, new_AGEMA_signal_3901, rd_I_n2274}), .b ({new_AGEMA_signal_3900, new_AGEMA_signal_3899, rd_I_n2276}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_4916, new_AGEMA_signal_4915, rd_I_n1835}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U985 ( .a ({new_AGEMA_signal_3910, new_AGEMA_signal_3909, rd_I_n2278}), .b ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, rd_I_n1832}), .c ({state_out_s2[355], state_out_s1[355], state_out_s0[355]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U984 ( .a ({new_AGEMA_signal_3908, new_AGEMA_signal_3907, rd_I_n2279}), .b ({new_AGEMA_signal_3906, new_AGEMA_signal_3905, rd_I_n2281}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({new_AGEMA_signal_4918, new_AGEMA_signal_4917, rd_I_n1832}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U980 ( .a ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, rd_I_n1829}), .b ({new_AGEMA_signal_4252, new_AGEMA_signal_4251, rd_I_n1828}), .c ({state_out_s2[9], state_out_s1[9], state_out_s0[9]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U979 ( .a ({new_AGEMA_signal_4250, new_AGEMA_signal_4249, rd_I_n1827}), .b ({new_AGEMA_signal_4920, new_AGEMA_signal_4919, rd_I_n1826}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, rd_I_n1829}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U977 ( .a ({new_AGEMA_signal_3916, new_AGEMA_signal_3915, rd_I_n2487}), .b ({new_AGEMA_signal_4922, new_AGEMA_signal_4921, rd_I_n1824}), .c ({state_out_s2[170], state_out_s1[170], state_out_s0[170]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U976 ( .a ({new_AGEMA_signal_3914, new_AGEMA_signal_3913, rd_I_n2489}), .b ({new_AGEMA_signal_3912, new_AGEMA_signal_3911, rd_I_n2486}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({new_AGEMA_signal_4922, new_AGEMA_signal_4921, rd_I_n1824}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U972 ( .a ({new_AGEMA_signal_5690, new_AGEMA_signal_5689, rd_I_n1821}), .b ({new_AGEMA_signal_4050, new_AGEMA_signal_4049, rd_I_n2583}), .c ({state_out_s2[348], state_out_s1[348], state_out_s0[348]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U971 ( .a ({new_AGEMA_signal_4924, new_AGEMA_signal_4923, rd_I_n1820}), .b ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, rd_I_n2586}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_5690, new_AGEMA_signal_5689, rd_I_n1821}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U969 ( .a ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, rd_I_n1819}), .b ({new_AGEMA_signal_4414, new_AGEMA_signal_4413, rd_I_n1818}), .c ({state_out_s2[109], state_out_s1[109], state_out_s0[109]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U968 ( .a ({new_AGEMA_signal_4926, new_AGEMA_signal_4925, rd_I_n1817}), .b ({new_AGEMA_signal_4412, new_AGEMA_signal_4411, rd_I_n1816}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, rd_I_n1819}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U966 ( .a ({new_AGEMA_signal_3938, new_AGEMA_signal_3937, rd_I_n2158}), .b ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, rd_I_n1814}), .c ({state_out_s2[142], state_out_s1[142], state_out_s0[142]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U965 ( .a ({new_AGEMA_signal_3940, new_AGEMA_signal_3939, rd_I_n2157}), .b ({new_AGEMA_signal_4946, new_AGEMA_signal_4945, rd_I_n2160}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, rd_I_n1814}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U964 ( .a ({new_AGEMA_signal_3922, new_AGEMA_signal_3921, rd_I_n2302}), .b ({new_AGEMA_signal_4928, new_AGEMA_signal_4927, rd_I_n1813}), .c ({state_out_s2[288], state_out_s1[288], state_out_s0[288]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U963 ( .a ({new_AGEMA_signal_3920, new_AGEMA_signal_3919, rd_I_n2303}), .b ({new_AGEMA_signal_3918, new_AGEMA_signal_3917, rd_I_n2305}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({new_AGEMA_signal_4928, new_AGEMA_signal_4927, rd_I_n1813}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U959 ( .a ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, rd_I_n1810}), .b ({new_AGEMA_signal_4232, new_AGEMA_signal_4231, rd_I_n2092}), .c ({state_out_s2[84], state_out_s1[84], state_out_s0[84]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U958 ( .a ({new_AGEMA_signal_4930, new_AGEMA_signal_4929, rd_I_n1809}), .b ({new_AGEMA_signal_4234, new_AGEMA_signal_4233, rd_I_n2095}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, rd_I_n1810}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U956 ( .a ({new_AGEMA_signal_4214, new_AGEMA_signal_4213, rd_I_n1808}), .b ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, rd_I_n1807}), .c ({state_out_s2[245], state_out_s1[245], state_out_s0[245]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U955 ( .a ({new_AGEMA_signal_4212, new_AGEMA_signal_4211, rd_I_n1806}), .b ({new_AGEMA_signal_4216, new_AGEMA_signal_4215, rd_I_n1805}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, rd_I_n1807}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U954 ( .a ({new_AGEMA_signal_4934, new_AGEMA_signal_4933, rd_I_n1804}), .b ({new_AGEMA_signal_3924, new_AGEMA_signal_3923, rd_I_n2433}), .c ({state_out_s2[263], state_out_s1[263], state_out_s0[263]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U952 ( .a ({new_AGEMA_signal_3928, new_AGEMA_signal_3927, rd_I_n2432}), .b ({new_AGEMA_signal_3926, new_AGEMA_signal_3925, rd_I_n2435}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_4934, new_AGEMA_signal_4933, rd_I_n1804}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U948 ( .a ({new_AGEMA_signal_4370, new_AGEMA_signal_4369, rd_I_n2267}), .b ({new_AGEMA_signal_4936, new_AGEMA_signal_4935, rd_I_n1799}), .c ({state_out_s2[47], state_out_s1[47], state_out_s0[47]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U947 ( .a ({new_AGEMA_signal_4372, new_AGEMA_signal_4371, rd_I_n2266}), .b ({new_AGEMA_signal_4368, new_AGEMA_signal_4367, rd_I_n2269}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({new_AGEMA_signal_4936, new_AGEMA_signal_4935, rd_I_n1799}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U946 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, rd_I_n1798}), .b ({new_AGEMA_signal_3954, new_AGEMA_signal_3953, rd_I_n2449}), .c ({state_out_s2[208], state_out_s1[208], state_out_s0[208]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U945 ( .a ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, rd_I_n1797}), .b ({new_AGEMA_signal_3956, new_AGEMA_signal_3955, rd_I_n2452}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, rd_I_n1798}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U943 ( .a ({new_AGEMA_signal_3934, new_AGEMA_signal_3933, rd_I_n2205}), .b ({new_AGEMA_signal_4940, new_AGEMA_signal_4939, rd_I_n1796}), .c ({state_out_s2[354], state_out_s1[354], state_out_s0[354]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U942 ( .a ({new_AGEMA_signal_3932, new_AGEMA_signal_3931, rd_I_n2206}), .b ({new_AGEMA_signal_3930, new_AGEMA_signal_3929, rd_I_n2208}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({new_AGEMA_signal_4940, new_AGEMA_signal_4939, rd_I_n1796}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U938 ( .a ({new_AGEMA_signal_4406, new_AGEMA_signal_4405, rd_I_n2496}), .b ({new_AGEMA_signal_4942, new_AGEMA_signal_4941, rd_I_n1792}), .c ({state_out_s2[2], state_out_s1[2], state_out_s0[2]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U937 ( .a ({new_AGEMA_signal_4408, new_AGEMA_signal_4407, rd_I_n2495}), .b ({new_AGEMA_signal_4404, new_AGEMA_signal_4403, rd_I_n2498}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_4942, new_AGEMA_signal_4941, rd_I_n1792}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U936 ( .a ({new_AGEMA_signal_3980, new_AGEMA_signal_3979, rd_I_n1968}), .b ({new_AGEMA_signal_4944, new_AGEMA_signal_4943, rd_I_n1791}), .c ({state_out_s2[163], state_out_s1[163], state_out_s0[163]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U935 ( .a ({new_AGEMA_signal_3978, new_AGEMA_signal_3977, rd_I_n1967}), .b ({new_AGEMA_signal_3982, new_AGEMA_signal_3981, rd_I_n1970}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({new_AGEMA_signal_4944, new_AGEMA_signal_4943, rd_I_n1791}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U934 ( .a ({new_AGEMA_signal_3940, new_AGEMA_signal_3939, rd_I_n2157}), .b ({new_AGEMA_signal_5714, new_AGEMA_signal_5713, rd_I_n1790}), .c ({state_out_s2[341], state_out_s1[341], state_out_s0[341]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U933 ( .a ({new_AGEMA_signal_3938, new_AGEMA_signal_3937, rd_I_n2158}), .b ({new_AGEMA_signal_4946, new_AGEMA_signal_4945, rd_I_n2160}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_5714, new_AGEMA_signal_5713, rd_I_n1790}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U925 ( .a ({new_AGEMA_signal_5716, new_AGEMA_signal_5715, rd_I_n1785}), .b ({new_AGEMA_signal_4312, new_AGEMA_signal_4311, rd_I_n2457}), .c ({state_out_s2[123], state_out_s1[123], state_out_s0[123]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U924 ( .a ({new_AGEMA_signal_4948, new_AGEMA_signal_4947, rd_I_n1784}), .b ({new_AGEMA_signal_4310, new_AGEMA_signal_4309, rd_I_n2460}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({new_AGEMA_signal_5716, new_AGEMA_signal_5715, rd_I_n1785}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U922 ( .a ({new_AGEMA_signal_3986, new_AGEMA_signal_3985, rd_I_n2390}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, rd_I_n1783}), .c ({state_out_s2[114], state_out_s1[114], state_out_s0[114]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U921 ( .a ({new_AGEMA_signal_3988, new_AGEMA_signal_3987, rd_I_n2389}), .b ({new_AGEMA_signal_3984, new_AGEMA_signal_3983, rd_I_n2392}), .clk (clk), .r ({Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, rd_I_n1783}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U920 ( .a ({new_AGEMA_signal_4094, new_AGEMA_signal_4093, rd_I_n1863}), .b ({new_AGEMA_signal_5720, new_AGEMA_signal_5719, rd_I_n1782}), .c ({state_out_s2[156], state_out_s1[156], state_out_s0[156]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U919 ( .a ({new_AGEMA_signal_4092, new_AGEMA_signal_4091, rd_I_n1862}), .b ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, rd_I_n1865}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771]}), .c ({new_AGEMA_signal_5720, new_AGEMA_signal_5719, rd_I_n1782}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U918 ( .a ({new_AGEMA_signal_5722, new_AGEMA_signal_5721, rd_I_n1781}), .b ({new_AGEMA_signal_4384, new_AGEMA_signal_4383, rd_I_n1780}), .c ({state_out_s2[147], state_out_s1[147], state_out_s0[147]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U917 ( .a ({new_AGEMA_signal_4952, new_AGEMA_signal_4951, rd_I_n1779}), .b ({new_AGEMA_signal_4382, new_AGEMA_signal_4381, rd_I_n1778}), .clk (clk), .r ({Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_5722, new_AGEMA_signal_5721, rd_I_n1781}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U915 ( .a ({new_AGEMA_signal_4316, new_AGEMA_signal_4315, rd_I_n2069}), .b ({new_AGEMA_signal_4954, new_AGEMA_signal_4953, rd_I_n1776}), .c ({state_out_s2[302], state_out_s1[302], state_out_s0[302]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U914 ( .a ({new_AGEMA_signal_4318, new_AGEMA_signal_4317, rd_I_n2068}), .b ({new_AGEMA_signal_4314, new_AGEMA_signal_4313, rd_I_n2071}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777]}), .c ({new_AGEMA_signal_4954, new_AGEMA_signal_4953, rd_I_n1776}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U913 ( .a ({new_AGEMA_signal_4256, new_AGEMA_signal_4255, rd_I_n2074}), .b ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, rd_I_n1775}), .c ({state_out_s2[293], state_out_s1[293], state_out_s0[293]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U912 ( .a ({new_AGEMA_signal_4254, new_AGEMA_signal_4253, rd_I_n2073}), .b ({new_AGEMA_signal_4258, new_AGEMA_signal_4257, rd_I_n2076}), .clk (clk), .r ({Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, rd_I_n1775}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U911 ( .a ({new_AGEMA_signal_4154, new_AGEMA_signal_4153, rd_I_n2236}), .b ({new_AGEMA_signal_4958, new_AGEMA_signal_4957, rd_I_n1774}), .c ({state_out_s2[108], state_out_s1[108], state_out_s0[108]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U910 ( .a ({new_AGEMA_signal_4152, new_AGEMA_signal_4151, rd_I_n2235}), .b ({new_AGEMA_signal_4156, new_AGEMA_signal_4155, rd_I_n2238}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783]}), .c ({new_AGEMA_signal_4958, new_AGEMA_signal_4957, rd_I_n1774}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U909 ( .a ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, rd_I_n1773}), .b ({new_AGEMA_signal_3942, new_AGEMA_signal_3941, rd_I_n2520}), .c ({state_out_s2[141], state_out_s1[141], state_out_s0[141]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U907 ( .a ({new_AGEMA_signal_3946, new_AGEMA_signal_3945, rd_I_n2523}), .b ({new_AGEMA_signal_4960, new_AGEMA_signal_4959, rd_I_n2521}), .clk (clk), .r ({Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, rd_I_n1773}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U899 ( .a ({new_AGEMA_signal_3952, new_AGEMA_signal_3951, rd_I_n1981}), .b ({new_AGEMA_signal_4962, new_AGEMA_signal_4961, rd_I_n1766}), .c ({state_out_s2[319], state_out_s1[319], state_out_s0[319]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U898 ( .a ({new_AGEMA_signal_3950, new_AGEMA_signal_3949, rd_I_n1982}), .b ({new_AGEMA_signal_3948, new_AGEMA_signal_3947, rd_I_n1984}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789]}), .c ({new_AGEMA_signal_4962, new_AGEMA_signal_4961, rd_I_n1766}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U894 ( .a ({new_AGEMA_signal_3958, new_AGEMA_signal_3957, rd_I_n2450}), .b ({new_AGEMA_signal_4964, new_AGEMA_signal_4963, rd_I_n1765}), .c ({state_out_s2[79], state_out_s1[79], state_out_s0[79]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U893 ( .a ({new_AGEMA_signal_3956, new_AGEMA_signal_3955, rd_I_n2452}), .b ({new_AGEMA_signal_3954, new_AGEMA_signal_3953, rd_I_n2449}), .clk (clk), .r ({Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_4964, new_AGEMA_signal_4963, rd_I_n1765}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U889 ( .a ({new_AGEMA_signal_3998, new_AGEMA_signal_3997, rd_I_n2298}), .b ({new_AGEMA_signal_4966, new_AGEMA_signal_4965, rd_I_n1763}), .c ({state_out_s2[240], state_out_s1[240], state_out_s0[240]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U888 ( .a ({new_AGEMA_signal_4000, new_AGEMA_signal_3999, rd_I_n2297}), .b ({new_AGEMA_signal_3996, new_AGEMA_signal_3995, rd_I_n2300}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795]}), .c ({new_AGEMA_signal_4966, new_AGEMA_signal_4965, rd_I_n1763}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U887 ( .a ({new_AGEMA_signal_4034, new_AGEMA_signal_4033, rd_I_n2197}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, rd_I_n1762}), .c ({state_out_s2[258], state_out_s1[258], state_out_s0[258]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U886 ( .a ({new_AGEMA_signal_4032, new_AGEMA_signal_4031, rd_I_n2196}), .b ({new_AGEMA_signal_4036, new_AGEMA_signal_4035, rd_I_n2199}), .clk (clk), .r ({Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, rd_I_n1762}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U885 ( .a ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, rd_I_n1761}), .b ({new_AGEMA_signal_4044, new_AGEMA_signal_4043, rd_I_n2319}), .c ({state_out_s2[92], state_out_s1[92], state_out_s0[92]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U884 ( .a ({new_AGEMA_signal_4970, new_AGEMA_signal_4969, rd_I_n1760}), .b ({new_AGEMA_signal_4046, new_AGEMA_signal_4045, rd_I_n2322}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801]}), .c ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, rd_I_n1761}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U882 ( .a ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, rd_I_n1759}), .b ({new_AGEMA_signal_4020, new_AGEMA_signal_4019, rd_I_n2025}), .c ({state_out_s2[83], state_out_s1[83], state_out_s0[83]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U881 ( .a ({new_AGEMA_signal_4972, new_AGEMA_signal_4971, rd_I_n1758}), .b ({new_AGEMA_signal_4022, new_AGEMA_signal_4021, rd_I_n2028}), .clk (clk), .r ({Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, rd_I_n1759}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U879 ( .a ({new_AGEMA_signal_4298, new_AGEMA_signal_4297, rd_I_n2349}), .b ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, rd_I_n1757}), .c ({state_out_s2[253], state_out_s1[253], state_out_s0[253]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U878 ( .a ({new_AGEMA_signal_4296, new_AGEMA_signal_4295, rd_I_n2348}), .b ({new_AGEMA_signal_4300, new_AGEMA_signal_4299, rd_I_n2351}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807]}), .c ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, rd_I_n1757}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U877 ( .a ({new_AGEMA_signal_4292, new_AGEMA_signal_4291, rd_I_n2344}), .b ({new_AGEMA_signal_4976, new_AGEMA_signal_4975, rd_I_n1756}), .c ({state_out_s2[244], state_out_s1[244], state_out_s0[244]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U876 ( .a ({new_AGEMA_signal_4290, new_AGEMA_signal_4289, rd_I_n2343}), .b ({new_AGEMA_signal_4294, new_AGEMA_signal_4293, rd_I_n2346}), .clk (clk), .r ({Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_4976, new_AGEMA_signal_4975, rd_I_n1756}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U875 ( .a ({new_AGEMA_signal_4130, new_AGEMA_signal_4129, rd_I_n2411}), .b ({new_AGEMA_signal_4978, new_AGEMA_signal_4977, rd_I_n1755}), .c ({state_out_s2[271], state_out_s1[271], state_out_s0[271]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U874 ( .a ({new_AGEMA_signal_4132, new_AGEMA_signal_4131, rd_I_n2410}), .b ({new_AGEMA_signal_4128, new_AGEMA_signal_4127, rd_I_n2413}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813]}), .c ({new_AGEMA_signal_4978, new_AGEMA_signal_4977, rd_I_n1755}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U873 ( .a ({new_AGEMA_signal_3964, new_AGEMA_signal_3963, rd_I_n2416}), .b ({new_AGEMA_signal_4980, new_AGEMA_signal_4979, rd_I_n1754}), .c ({state_out_s2[262], state_out_s1[262], state_out_s0[262]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U872 ( .a ({new_AGEMA_signal_3962, new_AGEMA_signal_3961, rd_I_n2418}), .b ({new_AGEMA_signal_3960, new_AGEMA_signal_3959, rd_I_n2415}), .clk (clk), .r ({Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_4980, new_AGEMA_signal_4979, rd_I_n1754}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U868 ( .a ({new_AGEMA_signal_3970, new_AGEMA_signal_3969, rd_I_n2500}), .b ({new_AGEMA_signal_4982, new_AGEMA_signal_4981, rd_I_n1752}), .c ({state_out_s2[46], state_out_s1[46], state_out_s0[46]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U867 ( .a ({new_AGEMA_signal_3968, new_AGEMA_signal_3967, rd_I_n2501}), .b ({new_AGEMA_signal_3966, new_AGEMA_signal_3965, rd_I_n2503}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819]}), .c ({new_AGEMA_signal_4982, new_AGEMA_signal_4981, rd_I_n1752}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U863 ( .a ({new_AGEMA_signal_4172, new_AGEMA_signal_4171, rd_I_n1750}), .b ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, rd_I_n1749}), .c ({state_out_s2[207], state_out_s1[207], state_out_s0[207]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U862 ( .a ({new_AGEMA_signal_4170, new_AGEMA_signal_4169, rd_I_n1748}), .b ({new_AGEMA_signal_4174, new_AGEMA_signal_4173, rd_I_n1747}), .clk (clk), .r ({Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_4984, new_AGEMA_signal_4983, rd_I_n1749}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U861 ( .a ({new_AGEMA_signal_5756, new_AGEMA_signal_5755, rd_I_n1746}), .b ({new_AGEMA_signal_4074, new_AGEMA_signal_4073, rd_I_n1839}), .c ({state_out_s2[353], state_out_s1[353], state_out_s0[353]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U860 ( .a ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, rd_I_n1745}), .b ({new_AGEMA_signal_4076, new_AGEMA_signal_4075, rd_I_n1842}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825]}), .c ({new_AGEMA_signal_5756, new_AGEMA_signal_5755, rd_I_n1746}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U858 ( .a ({new_AGEMA_signal_3976, new_AGEMA_signal_3975, rd_I_n2505}), .b ({new_AGEMA_signal_4988, new_AGEMA_signal_4987, rd_I_n1744}), .c ({state_out_s2[55], state_out_s1[55], state_out_s0[55]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U857 ( .a ({new_AGEMA_signal_3974, new_AGEMA_signal_3973, rd_I_n2506}), .b ({new_AGEMA_signal_3972, new_AGEMA_signal_3971, rd_I_n2508}), .clk (clk), .r ({Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_4988, new_AGEMA_signal_4987, rd_I_n1744}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U853 ( .a ({new_AGEMA_signal_4160, new_AGEMA_signal_4159, rd_I_n1960}), .b ({new_AGEMA_signal_4990, new_AGEMA_signal_4989, rd_I_n1742}), .c ({state_out_s2[216], state_out_s1[216], state_out_s0[216]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U852 ( .a ({new_AGEMA_signal_4158, new_AGEMA_signal_4157, rd_I_n1959}), .b ({new_AGEMA_signal_4162, new_AGEMA_signal_4161, rd_I_n1962}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831]}), .c ({new_AGEMA_signal_4990, new_AGEMA_signal_4989, rd_I_n1742}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U851 ( .a ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, rd_I_n1741}), .b ({new_AGEMA_signal_3978, new_AGEMA_signal_3977, rd_I_n1967}), .c ({state_out_s2[362], state_out_s1[362], state_out_s0[362]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U849 ( .a ({new_AGEMA_signal_3982, new_AGEMA_signal_3981, rd_I_n1970}), .b ({new_AGEMA_signal_3980, new_AGEMA_signal_3979, rd_I_n1968}), .clk (clk), .r ({Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, rd_I_n1741}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U845 ( .a ({new_AGEMA_signal_5764, new_AGEMA_signal_5763, rd_I_n1738}), .b ({new_AGEMA_signal_4140, new_AGEMA_signal_4139, rd_I_n2164}), .c ({state_out_s2[82], state_out_s1[82], state_out_s0[82]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U844 ( .a ({new_AGEMA_signal_4994, new_AGEMA_signal_4993, rd_I_n1737}), .b ({new_AGEMA_signal_4142, new_AGEMA_signal_4141, rd_I_n2167}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837]}), .c ({new_AGEMA_signal_5764, new_AGEMA_signal_5763, rd_I_n1738}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U842 ( .a ({new_AGEMA_signal_3988, new_AGEMA_signal_3987, rd_I_n2389}), .b ({new_AGEMA_signal_4996, new_AGEMA_signal_4995, rd_I_n1736}), .c ({state_out_s2[243], state_out_s1[243], state_out_s0[243]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U841 ( .a ({new_AGEMA_signal_3986, new_AGEMA_signal_3985, rd_I_n2390}), .b ({new_AGEMA_signal_3984, new_AGEMA_signal_3983, rd_I_n2392}), .clk (clk), .r ({Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_4996, new_AGEMA_signal_4995, rd_I_n1736}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U837 ( .a ({new_AGEMA_signal_4998, new_AGEMA_signal_4997, rd_I_n1732}), .b ({new_AGEMA_signal_3990, new_AGEMA_signal_3989, rd_I_n2364}), .c ({state_out_s2[261], state_out_s1[261], state_out_s0[261]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U835 ( .a ({new_AGEMA_signal_3994, new_AGEMA_signal_3993, rd_I_n2363}), .b ({new_AGEMA_signal_3992, new_AGEMA_signal_3991, rd_I_n2366}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843]}), .c ({new_AGEMA_signal_4998, new_AGEMA_signal_4997, rd_I_n1732}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U831 ( .a ({new_AGEMA_signal_5770, new_AGEMA_signal_5769, rd_I_n1728}), .b ({new_AGEMA_signal_4430, new_AGEMA_signal_4429, rd_I_n2453}), .c ({state_out_s2[100], state_out_s1[100], state_out_s0[100]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U830 ( .a ({new_AGEMA_signal_4432, new_AGEMA_signal_4431, rd_I_n2456}), .b ({new_AGEMA_signal_5000, new_AGEMA_signal_4999, rd_I_n1727}), .clk (clk), .r ({Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_5770, new_AGEMA_signal_5769, rd_I_n1728}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U828 ( .a ({new_AGEMA_signal_4088, new_AGEMA_signal_4087, rd_I_n2153}), .b ({new_AGEMA_signal_5002, new_AGEMA_signal_5001, rd_I_n1726}), .c ({state_out_s2[133], state_out_s1[133], state_out_s0[133]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U827 ( .a ({new_AGEMA_signal_4086, new_AGEMA_signal_4085, rd_I_n2152}), .b ({new_AGEMA_signal_4090, new_AGEMA_signal_4089, rd_I_n2155}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849]}), .c ({new_AGEMA_signal_5002, new_AGEMA_signal_5001, rd_I_n1726}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U826 ( .a ({new_AGEMA_signal_4000, new_AGEMA_signal_3999, rd_I_n2297}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, rd_I_n1725}), .c ({state_out_s2[311], state_out_s1[311], state_out_s0[311]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U825 ( .a ({new_AGEMA_signal_3998, new_AGEMA_signal_3997, rd_I_n2298}), .b ({new_AGEMA_signal_3996, new_AGEMA_signal_3995, rd_I_n2300}), .clk (clk), .r ({Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, rd_I_n1725}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U821 ( .a ({new_AGEMA_signal_5006, new_AGEMA_signal_5005, rd_I_n1722}), .b ({new_AGEMA_signal_4002, new_AGEMA_signal_4001, rd_I_n2125}), .c ({state_out_s2[77], state_out_s1[77], state_out_s0[77]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U819 ( .a ({new_AGEMA_signal_4006, new_AGEMA_signal_4005, rd_I_n2128}), .b ({new_AGEMA_signal_4004, new_AGEMA_signal_4003, rd_I_n2126}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855]}), .c ({new_AGEMA_signal_5006, new_AGEMA_signal_5005, rd_I_n1722}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U815 ( .a ({new_AGEMA_signal_4412, new_AGEMA_signal_4411, rd_I_n1816}), .b ({new_AGEMA_signal_5008, new_AGEMA_signal_5007, rd_I_n1718}), .c ({state_out_s2[238], state_out_s1[238], state_out_s0[238]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U814 ( .a ({new_AGEMA_signal_4410, new_AGEMA_signal_4409, rd_I_n1815}), .b ({new_AGEMA_signal_4414, new_AGEMA_signal_4413, rd_I_n1818}), .clk (clk), .r ({Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_5008, new_AGEMA_signal_5007, rd_I_n1718}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U813 ( .a ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, rd_I_n1717}), .b ({new_AGEMA_signal_4008, new_AGEMA_signal_4007, rd_I_n2181}), .c ({state_out_s2[256], state_out_s1[256], state_out_s0[256]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U811 ( .a ({new_AGEMA_signal_4012, new_AGEMA_signal_4011, rd_I_n2180}), .b ({new_AGEMA_signal_4010, new_AGEMA_signal_4009, rd_I_n2183}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861]}), .c ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, rd_I_n1717}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U805 ( .a ({new_AGEMA_signal_5012, new_AGEMA_signal_5011, rd_I_n1714}), .b ({new_AGEMA_signal_4014, new_AGEMA_signal_4013, rd_I_n2436}), .c ({state_out_s2[72], state_out_s1[72], state_out_s0[72]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U803 ( .a ({new_AGEMA_signal_4018, new_AGEMA_signal_4017, rd_I_n2439}), .b ({new_AGEMA_signal_4016, new_AGEMA_signal_4015, rd_I_n2437}), .clk (clk), .r ({Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_5012, new_AGEMA_signal_5011, rd_I_n1714}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U797 ( .a ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, rd_I_n1710}), .b ({new_AGEMA_signal_4276, new_AGEMA_signal_4275, rd_I_n1709}), .c ({state_out_s2[233], state_out_s1[233], state_out_s0[233]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U796 ( .a ({new_AGEMA_signal_5014, new_AGEMA_signal_5013, rd_I_n1708}), .b ({new_AGEMA_signal_4274, new_AGEMA_signal_4273, rd_I_n1707}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867]}), .c ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, rd_I_n1710}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U794 ( .a ({new_AGEMA_signal_4024, new_AGEMA_signal_4023, rd_I_n2026}), .b ({new_AGEMA_signal_5016, new_AGEMA_signal_5015, rd_I_n1705}), .c ({state_out_s2[283], state_out_s1[283], state_out_s0[283]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U793 ( .a ({new_AGEMA_signal_4022, new_AGEMA_signal_4021, rd_I_n2028}), .b ({new_AGEMA_signal_4020, new_AGEMA_signal_4019, rd_I_n2025}), .clk (clk), .r ({Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_5016, new_AGEMA_signal_5015, rd_I_n1705}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U789 ( .a ({new_AGEMA_signal_5160, new_AGEMA_signal_5159, rd_I_n1857}), .b ({new_AGEMA_signal_5018, new_AGEMA_signal_5017, rd_I_n1704}), .c ({state_out_s2[6], state_out_s1[6], state_out_s0[6]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U788 ( .a ({new_AGEMA_signal_4320, new_AGEMA_signal_4319, rd_I_n1856}), .b ({new_AGEMA_signal_4324, new_AGEMA_signal_4323, rd_I_n1859}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873]}), .c ({new_AGEMA_signal_5018, new_AGEMA_signal_5017, rd_I_n1704}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U787 ( .a ({new_AGEMA_signal_5020, new_AGEMA_signal_5019, rd_I_n1703}), .b ({new_AGEMA_signal_4026, new_AGEMA_signal_4025, rd_I_n2368}), .c ({state_out_s2[167], state_out_s1[167], state_out_s0[167]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U785 ( .a ({new_AGEMA_signal_4030, new_AGEMA_signal_4029, rd_I_n2367}), .b ({new_AGEMA_signal_4028, new_AGEMA_signal_4027, rd_I_n2370}), .clk (clk), .r ({Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_5020, new_AGEMA_signal_5019, rd_I_n1703}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U778 ( .a ({new_AGEMA_signal_5792, new_AGEMA_signal_5791, rd_I_n1697}), .b ({new_AGEMA_signal_4278, new_AGEMA_signal_4277, rd_I_n2107}), .c ({state_out_s2[345], state_out_s1[345], state_out_s0[345]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U777 ( .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, rd_I_n1696}), .b ({new_AGEMA_signal_5144, new_AGEMA_signal_5143, rd_I_n2110}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879]}), .c ({new_AGEMA_signal_5792, new_AGEMA_signal_5791, rd_I_n1697}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U775 ( .a ({new_AGEMA_signal_5024, new_AGEMA_signal_5023, rd_I_n1695}), .b ({new_AGEMA_signal_4032, new_AGEMA_signal_4031, rd_I_n2196}), .c ({state_out_s2[90], state_out_s1[90], state_out_s0[90]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U773 ( .a ({new_AGEMA_signal_4036, new_AGEMA_signal_4035, rd_I_n2199}), .b ({new_AGEMA_signal_4034, new_AGEMA_signal_4033, rd_I_n2197}), .clk (clk), .r ({Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_5024, new_AGEMA_signal_5023, rd_I_n1695}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U769 ( .a ({new_AGEMA_signal_5026, new_AGEMA_signal_5025, rd_I_n1691}), .b ({new_AGEMA_signal_4038, new_AGEMA_signal_4037, rd_I_n2065}), .c ({state_out_s2[81], state_out_s1[81], state_out_s0[81]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U767 ( .a ({new_AGEMA_signal_4042, new_AGEMA_signal_4041, rd_I_n2064}), .b ({new_AGEMA_signal_4040, new_AGEMA_signal_4039, rd_I_n2067}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885]}), .c ({new_AGEMA_signal_5026, new_AGEMA_signal_5025, rd_I_n1691}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U761 ( .a ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, rd_I_n1687}), .b ({new_AGEMA_signal_4336, new_AGEMA_signal_4335, rd_I_n2283}), .c ({state_out_s2[251], state_out_s1[251], state_out_s0[251]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U760 ( .a ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, rd_I_n1686}), .b ({new_AGEMA_signal_4334, new_AGEMA_signal_4333, rd_I_n2286}), .clk (clk), .r ({Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_5798, new_AGEMA_signal_5797, rd_I_n1687}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U758 ( .a ({new_AGEMA_signal_4328, new_AGEMA_signal_4327, rd_I_n1685}), .b ({new_AGEMA_signal_5030, new_AGEMA_signal_5029, rd_I_n1684}), .c ({state_out_s2[242], state_out_s1[242], state_out_s0[242]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U757 ( .a ({new_AGEMA_signal_4326, new_AGEMA_signal_4325, rd_I_n1683}), .b ({new_AGEMA_signal_4330, new_AGEMA_signal_4329, rd_I_n1682}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891]}), .c ({new_AGEMA_signal_5030, new_AGEMA_signal_5029, rd_I_n1684}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U756 ( .a ({new_AGEMA_signal_4262, new_AGEMA_signal_4261, rd_I_n2315}), .b ({new_AGEMA_signal_5032, new_AGEMA_signal_5031, rd_I_n1681}), .c ({state_out_s2[269], state_out_s1[269], state_out_s0[269]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U755 ( .a ({new_AGEMA_signal_4264, new_AGEMA_signal_4263, rd_I_n2314}), .b ({new_AGEMA_signal_4260, new_AGEMA_signal_4259, rd_I_n2317}), .clk (clk), .r ({Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_5032, new_AGEMA_signal_5031, rd_I_n1681}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U754 ( .a ({new_AGEMA_signal_4048, new_AGEMA_signal_4047, rd_I_n2320}), .b ({new_AGEMA_signal_5034, new_AGEMA_signal_5033, rd_I_n1680}), .c ({state_out_s2[260], state_out_s1[260], state_out_s0[260]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U753 ( .a ({new_AGEMA_signal_4046, new_AGEMA_signal_4045, rd_I_n2322}), .b ({new_AGEMA_signal_4044, new_AGEMA_signal_4043, rd_I_n2319}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897]}), .c ({new_AGEMA_signal_5034, new_AGEMA_signal_5033, rd_I_n1680}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U749 ( .a ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, rd_I_n1678}), .b ({new_AGEMA_signal_4216, new_AGEMA_signal_4215, rd_I_n1805}), .c ({state_out_s2[116], state_out_s1[116], state_out_s0[116]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U748 ( .a ({new_AGEMA_signal_5036, new_AGEMA_signal_5035, rd_I_n1677}), .b ({new_AGEMA_signal_4214, new_AGEMA_signal_4213, rd_I_n1808}), .clk (clk), .r ({Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_5806, new_AGEMA_signal_5805, rd_I_n1678}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U746 ( .a ({new_AGEMA_signal_4184, new_AGEMA_signal_4183, rd_I_n1941}), .b ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, rd_I_n1676}), .c ({state_out_s2[107], state_out_s1[107], state_out_s0[107]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U745 ( .a ({new_AGEMA_signal_4186, new_AGEMA_signal_4185, rd_I_n1940}), .b ({new_AGEMA_signal_4182, new_AGEMA_signal_4181, rd_I_n1943}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903]}), .c ({new_AGEMA_signal_5038, new_AGEMA_signal_5037, rd_I_n1676}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U744 ( .a ({new_AGEMA_signal_4054, new_AGEMA_signal_4053, rd_I_n2584}), .b ({new_AGEMA_signal_5810, new_AGEMA_signal_5809, rd_I_n1675}), .c ({state_out_s2[149], state_out_s1[149], state_out_s0[149]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U743 ( .a ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, rd_I_n2586}), .b ({new_AGEMA_signal_4050, new_AGEMA_signal_4049, rd_I_n2583}), .clk (clk), .r ({Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_5810, new_AGEMA_signal_5809, rd_I_n1675}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U737 ( .a ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, rd_I_n1670}), .b ({new_AGEMA_signal_4056, new_AGEMA_signal_4055, rd_I_n2580}), .c ({state_out_s2[140], state_out_s1[140], state_out_s0[140]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U735 ( .a ({new_AGEMA_signal_4060, new_AGEMA_signal_4059, rd_I_n2579}), .b ({new_AGEMA_signal_5042, new_AGEMA_signal_5041, rd_I_n2582}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909]}), .c ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, rd_I_n1670}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U727 ( .a ({new_AGEMA_signal_5044, new_AGEMA_signal_5043, rd_I_n1663}), .b ({new_AGEMA_signal_4062, new_AGEMA_signal_4061, rd_I_n1904}), .c ({state_out_s2[318], state_out_s1[318], state_out_s0[318]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U725 ( .a ({new_AGEMA_signal_4066, new_AGEMA_signal_4065, rd_I_n1903}), .b ({new_AGEMA_signal_4064, new_AGEMA_signal_4063, rd_I_n1906}), .clk (clk), .r ({Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_5044, new_AGEMA_signal_5043, rd_I_n1663}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U721 ( .a ({new_AGEMA_signal_4072, new_AGEMA_signal_4071, rd_I_n1900}), .b ({new_AGEMA_signal_5046, new_AGEMA_signal_5045, rd_I_n1660}), .c ({state_out_s2[295], state_out_s1[295], state_out_s0[295]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U720 ( .a ({new_AGEMA_signal_4070, new_AGEMA_signal_4069, rd_I_n1902}), .b ({new_AGEMA_signal_4068, new_AGEMA_signal_4067, rd_I_n1899}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915]}), .c ({new_AGEMA_signal_5046, new_AGEMA_signal_5045, rd_I_n1660}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U716 ( .a ({new_AGEMA_signal_4424, new_AGEMA_signal_4423, rd_I_n2491}), .b ({new_AGEMA_signal_5048, new_AGEMA_signal_5047, rd_I_n1659}), .c ({state_out_s2[25], state_out_s1[25], state_out_s0[25]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U715 ( .a ({new_AGEMA_signal_4426, new_AGEMA_signal_4425, rd_I_n2490}), .b ({new_AGEMA_signal_4422, new_AGEMA_signal_4421, rd_I_n2493}), .clk (clk), .r ({Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_5048, new_AGEMA_signal_5047, rd_I_n1659}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U714 ( .a ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, rd_I_n1658}), .b ({new_AGEMA_signal_4446, new_AGEMA_signal_4445, rd_I_n1657}), .c ({state_out_s2[16], state_out_s1[16], state_out_s0[16]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U713 ( .a ({new_AGEMA_signal_5050, new_AGEMA_signal_5049, rd_I_n1656}), .b ({new_AGEMA_signal_4448, new_AGEMA_signal_4447, rd_I_n1655}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921]}), .c ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, rd_I_n1658}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U711 ( .a ({new_AGEMA_signal_4078, new_AGEMA_signal_4077, rd_I_n1840}), .b ({new_AGEMA_signal_5052, new_AGEMA_signal_5051, rd_I_n1653}), .c ({state_out_s2[186], state_out_s1[186], state_out_s0[186]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U710 ( .a ({new_AGEMA_signal_4076, new_AGEMA_signal_4075, rd_I_n1842}), .b ({new_AGEMA_signal_4074, new_AGEMA_signal_4073, rd_I_n1839}), .clk (clk), .r ({Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_5052, new_AGEMA_signal_5051, rd_I_n1653}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U706 ( .a ({new_AGEMA_signal_4084, new_AGEMA_signal_4083, rd_I_n2309}), .b ({new_AGEMA_signal_5054, new_AGEMA_signal_5053, rd_I_n1651}), .c ({state_out_s2[177], state_out_s1[177], state_out_s0[177]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U705 ( .a ({new_AGEMA_signal_4082, new_AGEMA_signal_4081, rd_I_n2310}), .b ({new_AGEMA_signal_4080, new_AGEMA_signal_4079, rd_I_n2312}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927]}), .c ({new_AGEMA_signal_5054, new_AGEMA_signal_5053, rd_I_n1651}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U701 ( .a ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, rd_I_n1648}), .b ({new_AGEMA_signal_4086, new_AGEMA_signal_4085, rd_I_n2152}), .c ({state_out_s2[332], state_out_s1[332], state_out_s0[332]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U699 ( .a ({new_AGEMA_signal_4090, new_AGEMA_signal_4089, rd_I_n2155}), .b ({new_AGEMA_signal_4088, new_AGEMA_signal_4087, rd_I_n2153}), .clk (clk), .r ({Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_5056, new_AGEMA_signal_5055, rd_I_n1648}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U695 ( .a ({new_AGEMA_signal_5828, new_AGEMA_signal_5827, rd_I_n1646}), .b ({new_AGEMA_signal_4092, new_AGEMA_signal_4091, rd_I_n1862}), .c ({state_out_s2[323], state_out_s1[323], state_out_s0[323]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U693 ( .a ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, rd_I_n1865}), .b ({new_AGEMA_signal_4094, new_AGEMA_signal_4093, rd_I_n1863}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933]}), .c ({new_AGEMA_signal_5828, new_AGEMA_signal_5827, rd_I_n1646}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U689 ( .a ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, rd_I_n1643}), .b ({new_AGEMA_signal_4174, new_AGEMA_signal_4173, rd_I_n1747}), .c ({state_out_s2[78], state_out_s1[78], state_out_s0[78]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U688 ( .a ({new_AGEMA_signal_5060, new_AGEMA_signal_5059, rd_I_n1642}), .b ({new_AGEMA_signal_4172, new_AGEMA_signal_4171, rd_I_n1750}), .clk (clk), .r ({Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, rd_I_n1643}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U686 ( .a ({new_AGEMA_signal_4360, new_AGEMA_signal_4359, rd_I_n1978}), .b ({new_AGEMA_signal_5062, new_AGEMA_signal_5061, rd_I_n1641}), .c ({state_out_s2[239], state_out_s1[239], state_out_s0[239]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U685 ( .a ({new_AGEMA_signal_4356, new_AGEMA_signal_4355, rd_I_n1976}), .b ({new_AGEMA_signal_4358, new_AGEMA_signal_4357, rd_I_n1979}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939]}), .c ({new_AGEMA_signal_5062, new_AGEMA_signal_5061, rd_I_n1641}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U684 ( .a ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, rd_I_n1640}), .b ({new_AGEMA_signal_4098, new_AGEMA_signal_4097, rd_I_n2230}), .c ({state_out_s2[257], state_out_s1[257], state_out_s0[257]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U682 ( .a ({new_AGEMA_signal_4102, new_AGEMA_signal_4101, rd_I_n2233}), .b ({new_AGEMA_signal_4100, new_AGEMA_signal_4099, rd_I_n2231}), .clk (clk), .r ({Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, rd_I_n1640}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U676 ( .a ({new_AGEMA_signal_4108, new_AGEMA_signal_4107, rd_I_n2394}), .b ({new_AGEMA_signal_5066, new_AGEMA_signal_5065, rd_I_n1636}), .c ({state_out_s2[7], state_out_s1[7], state_out_s0[7]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U675 ( .a ({new_AGEMA_signal_4106, new_AGEMA_signal_4105, rd_I_n2395}), .b ({new_AGEMA_signal_4104, new_AGEMA_signal_4103, rd_I_n2397}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945]}), .c ({new_AGEMA_signal_5066, new_AGEMA_signal_5065, rd_I_n1636}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U669 ( .a ({new_AGEMA_signal_5068, new_AGEMA_signal_5067, rd_I_n1631}), .b ({new_AGEMA_signal_4110, new_AGEMA_signal_4109, rd_I_n2420}), .c ({state_out_s2[168], state_out_s1[168], state_out_s0[168]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U667 ( .a ({new_AGEMA_signal_4114, new_AGEMA_signal_4113, rd_I_n2419}), .b ({new_AGEMA_signal_4112, new_AGEMA_signal_4111, rd_I_n2422}), .clk (clk), .r ({Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_5068, new_AGEMA_signal_5067, rd_I_n1631}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U663 ( .a ({new_AGEMA_signal_4382, new_AGEMA_signal_4381, rd_I_n1778}), .b ({new_AGEMA_signal_5070, new_AGEMA_signal_5069, rd_I_n1627}), .c ({state_out_s2[346], state_out_s1[346], state_out_s0[346]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U662 ( .a ({new_AGEMA_signal_4380, new_AGEMA_signal_4379, rd_I_n1777}), .b ({new_AGEMA_signal_4384, new_AGEMA_signal_4383, rd_I_n1780}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951]}), .c ({new_AGEMA_signal_5070, new_AGEMA_signal_5069, rd_I_n1627}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U661 ( .a ({new_AGEMA_signal_4202, new_AGEMA_signal_4201, rd_I_n1869}), .b ({new_AGEMA_signal_5072, new_AGEMA_signal_5071, rd_I_n1626}), .c ({state_out_s2[106], state_out_s1[106], state_out_s0[106]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U660 ( .a ({new_AGEMA_signal_4200, new_AGEMA_signal_4199, rd_I_n1868}), .b ({new_AGEMA_signal_4204, new_AGEMA_signal_4203, rd_I_n1871}), .clk (clk), .r ({Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_5072, new_AGEMA_signal_5071, rd_I_n1626}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U659 ( .a ({new_AGEMA_signal_4120, new_AGEMA_signal_4119, rd_I_n2600}), .b ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, rd_I_n1625}), .c ({state_out_s2[139], state_out_s1[139], state_out_s0[139]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U658 ( .a ({new_AGEMA_signal_5074, new_AGEMA_signal_5073, rd_I_n2601}), .b ({new_AGEMA_signal_4116, new_AGEMA_signal_4115, rd_I_n2603}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957]}), .c ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, rd_I_n1625}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U647 ( .a ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, rd_I_n1618}), .b ({new_AGEMA_signal_4122, new_AGEMA_signal_4121, rd_I_n2556}), .c ({state_out_s2[317], state_out_s1[317], state_out_s0[317]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U645 ( .a ({new_AGEMA_signal_4126, new_AGEMA_signal_4125, rd_I_n2559}), .b ({new_AGEMA_signal_4124, new_AGEMA_signal_4123, rd_I_n2557}), .clk (clk), .r ({Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, rd_I_n1618}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U641 ( .a ({new_AGEMA_signal_4132, new_AGEMA_signal_4131, rd_I_n2410}), .b ({new_AGEMA_signal_5078, new_AGEMA_signal_5077, rd_I_n1615}), .c ({state_out_s2[71], state_out_s1[71], state_out_s0[71]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U640 ( .a ({new_AGEMA_signal_4130, new_AGEMA_signal_4129, rd_I_n2411}), .b ({new_AGEMA_signal_4128, new_AGEMA_signal_4127, rd_I_n2413}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963]}), .c ({new_AGEMA_signal_5078, new_AGEMA_signal_5077, rd_I_n1615}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U636 ( .a ({new_AGEMA_signal_5080, new_AGEMA_signal_5079, rd_I_n1613}), .b ({new_AGEMA_signal_4134, new_AGEMA_signal_4133, rd_I_n2400}), .c ({state_out_s2[232], state_out_s1[232], state_out_s0[232]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U634 ( .a ({new_AGEMA_signal_4138, new_AGEMA_signal_4137, rd_I_n2399}), .b ({new_AGEMA_signal_4136, new_AGEMA_signal_4135, rd_I_n2402}), .clk (clk), .r ({Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_5080, new_AGEMA_signal_5079, rd_I_n1613}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U630 ( .a ({new_AGEMA_signal_4144, new_AGEMA_signal_4143, rd_I_n2165}), .b ({new_AGEMA_signal_5082, new_AGEMA_signal_5081, rd_I_n1610}), .c ({state_out_s2[282], state_out_s1[282], state_out_s0[282]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U629 ( .a ({new_AGEMA_signal_4142, new_AGEMA_signal_4141, rd_I_n2167}), .b ({new_AGEMA_signal_4140, new_AGEMA_signal_4139, rd_I_n2164}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969]}), .c ({new_AGEMA_signal_5082, new_AGEMA_signal_5081, rd_I_n1610}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U623 ( .a ({new_AGEMA_signal_4150, new_AGEMA_signal_4149, rd_I_n2047}), .b ({new_AGEMA_signal_5084, new_AGEMA_signal_5083, rd_I_n1605}), .c ({state_out_s2[76], state_out_s1[76], state_out_s0[76]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U622 ( .a ({new_AGEMA_signal_4148, new_AGEMA_signal_4147, rd_I_n2048}), .b ({new_AGEMA_signal_4146, new_AGEMA_signal_4145, rd_I_n2050}), .clk (clk), .r ({Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_5084, new_AGEMA_signal_5083, rd_I_n1605}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U616 ( .a ({new_AGEMA_signal_5086, new_AGEMA_signal_5085, rd_I_n1599}), .b ({new_AGEMA_signal_4152, new_AGEMA_signal_4151, rd_I_n2235}), .c ({state_out_s2[237], state_out_s1[237], state_out_s0[237]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U614 ( .a ({new_AGEMA_signal_4156, new_AGEMA_signal_4155, rd_I_n2238}), .b ({new_AGEMA_signal_4154, new_AGEMA_signal_4153, rd_I_n2236}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975]}), .c ({new_AGEMA_signal_5086, new_AGEMA_signal_5085, rd_I_n1599}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U607 ( .a ({new_AGEMA_signal_5088, new_AGEMA_signal_5087, rd_I_n1594}), .b ({new_AGEMA_signal_4158, new_AGEMA_signal_4157, rd_I_n1959}), .c ({state_out_s2[287], state_out_s1[287], state_out_s0[287]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U604 ( .a ({new_AGEMA_signal_4162, new_AGEMA_signal_4161, rd_I_n1962}), .b ({new_AGEMA_signal_4160, new_AGEMA_signal_4159, rd_I_n1960}), .clk (clk), .r ({Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_5088, new_AGEMA_signal_5087, rd_I_n1594}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U597 ( .a ({new_AGEMA_signal_5090, new_AGEMA_signal_5089, rd_I_n1587}), .b ({new_AGEMA_signal_4164, new_AGEMA_signal_4163, rd_I_n2191}), .c ({state_out_s2[67], state_out_s1[67], state_out_s0[67]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U595 ( .a ({new_AGEMA_signal_4168, new_AGEMA_signal_4167, rd_I_n2192}), .b ({new_AGEMA_signal_4166, new_AGEMA_signal_4165, rd_I_n2194}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981]}), .c ({new_AGEMA_signal_5090, new_AGEMA_signal_5089, rd_I_n1587}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U584 ( .a ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, rd_I_n1581}), .b ({new_AGEMA_signal_4348, new_AGEMA_signal_4347, rd_I_n2287}), .c ({state_out_s2[228], state_out_s1[228], state_out_s0[228]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U583 ( .a ({new_AGEMA_signal_5092, new_AGEMA_signal_5091, rd_I_n1580}), .b ({new_AGEMA_signal_4346, new_AGEMA_signal_4345, rd_I_n2290}), .clk (clk), .r ({Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, rd_I_n1581}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U581 ( .a ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, rd_I_n1579}), .b ({new_AGEMA_signal_4170, new_AGEMA_signal_4169, rd_I_n1748}), .c ({state_out_s2[278], state_out_s1[278], state_out_s0[278]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U579 ( .a ({new_AGEMA_signal_4174, new_AGEMA_signal_4173, rd_I_n1747}), .b ({new_AGEMA_signal_4172, new_AGEMA_signal_4171, rd_I_n1750}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987]}), .c ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, rd_I_n1579}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U573 ( .a ({new_AGEMA_signal_5096, new_AGEMA_signal_5095, rd_I_n1576}), .b ({new_AGEMA_signal_4176, new_AGEMA_signal_4175, rd_I_n2087}), .c ({state_out_s2[75], state_out_s1[75], state_out_s0[75]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U571 ( .a ({new_AGEMA_signal_4180, new_AGEMA_signal_4179, rd_I_n2090}), .b ({new_AGEMA_signal_4178, new_AGEMA_signal_4177, rd_I_n2088}), .clk (clk), .r ({Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_5096, new_AGEMA_signal_5095, rd_I_n1576}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U562 ( .a ({new_AGEMA_signal_4186, new_AGEMA_signal_4185, rd_I_n1940}), .b ({new_AGEMA_signal_5098, new_AGEMA_signal_5097, rd_I_n1570}), .c ({state_out_s2[236], state_out_s1[236], state_out_s0[236]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U561 ( .a ({new_AGEMA_signal_4184, new_AGEMA_signal_4183, rd_I_n1941}), .b ({new_AGEMA_signal_4182, new_AGEMA_signal_4181, rd_I_n1943}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993]}), .c ({new_AGEMA_signal_5098, new_AGEMA_signal_5097, rd_I_n1570}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U555 ( .a ({new_AGEMA_signal_5100, new_AGEMA_signal_5099, rd_I_n1565}), .b ({new_AGEMA_signal_4188, new_AGEMA_signal_4187, rd_I_n2136}), .c ({state_out_s2[286], state_out_s1[286], state_out_s0[286]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U552 ( .a ({new_AGEMA_signal_4192, new_AGEMA_signal_4191, rd_I_n2135}), .b ({new_AGEMA_signal_4190, new_AGEMA_signal_4189, rd_I_n2138}), .clk (clk), .r ({Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_5100, new_AGEMA_signal_5099, rd_I_n1565}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U543 ( .a ({new_AGEMA_signal_5102, new_AGEMA_signal_5101, rd_I_n1558}), .b ({new_AGEMA_signal_4194, new_AGEMA_signal_4193, rd_I_n2005}), .c ({state_out_s2[74], state_out_s1[74], state_out_s0[74]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U541 ( .a ({new_AGEMA_signal_4198, new_AGEMA_signal_4197, rd_I_n2008}), .b ({new_AGEMA_signal_4196, new_AGEMA_signal_4195, rd_I_n2006}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999]}), .c ({new_AGEMA_signal_5102, new_AGEMA_signal_5101, rd_I_n1558}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U532 ( .a ({new_AGEMA_signal_5104, new_AGEMA_signal_5103, rd_I_n1552}), .b ({new_AGEMA_signal_4200, new_AGEMA_signal_4199, rd_I_n1868}), .c ({state_out_s2[235], state_out_s1[235], state_out_s0[235]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U530 ( .a ({new_AGEMA_signal_4204, new_AGEMA_signal_4203, rd_I_n1871}), .b ({new_AGEMA_signal_4202, new_AGEMA_signal_4201, rd_I_n1869}), .clk (clk), .r ({Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_5104, new_AGEMA_signal_5103, rd_I_n1552}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U521 ( .a ({new_AGEMA_signal_5106, new_AGEMA_signal_5105, rd_I_n1547}), .b ({new_AGEMA_signal_4206, new_AGEMA_signal_4205, rd_I_n2056}), .c ({state_out_s2[285], state_out_s1[285], state_out_s0[285]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U516 ( .a ({new_AGEMA_signal_4210, new_AGEMA_signal_4209, rd_I_n2055}), .b ({new_AGEMA_signal_4208, new_AGEMA_signal_4207, rd_I_n2058}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005]}), .c ({new_AGEMA_signal_5106, new_AGEMA_signal_5105, rd_I_n1547}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U507 ( .a ({new_AGEMA_signal_4226, new_AGEMA_signal_4225, rd_I_n2542}), .b ({new_AGEMA_signal_5108, new_AGEMA_signal_5107, rd_I_n1540}), .c ({state_out_s2[105], state_out_s1[105], state_out_s0[105]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U506 ( .a ({new_AGEMA_signal_4228, new_AGEMA_signal_4227, rd_I_n2541}), .b ({new_AGEMA_signal_4224, new_AGEMA_signal_4223, rd_I_n2544}), .clk (clk), .r ({Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_5108, new_AGEMA_signal_5107, rd_I_n1540}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U505 ( .a ({new_AGEMA_signal_4250, new_AGEMA_signal_4249, rd_I_n1827}), .b ({new_AGEMA_signal_5110, new_AGEMA_signal_5109, rd_I_n1539}), .c ({state_out_s2[138], state_out_s1[138], state_out_s0[138]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U504 ( .a ({new_AGEMA_signal_4248, new_AGEMA_signal_4247, rd_I_n1825}), .b ({new_AGEMA_signal_4252, new_AGEMA_signal_4251, rd_I_n1828}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011]}), .c ({new_AGEMA_signal_5110, new_AGEMA_signal_5109, rd_I_n1539}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U503 ( .a ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, rd_I_n1538}), .b ({new_AGEMA_signal_4212, new_AGEMA_signal_4211, rd_I_n1806}), .c ({state_out_s2[316], state_out_s1[316], state_out_s0[316]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U501 ( .a ({new_AGEMA_signal_4216, new_AGEMA_signal_4215, rd_I_n1805}), .b ({new_AGEMA_signal_4214, new_AGEMA_signal_4213, rd_I_n1808}), .clk (clk), .r ({Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, rd_I_n1538}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U495 ( .a ({new_AGEMA_signal_5114, new_AGEMA_signal_5113, rd_I_n1534}), .b ({new_AGEMA_signal_4218, new_AGEMA_signal_4217, rd_I_n2477}), .c ({state_out_s2[73], state_out_s1[73], state_out_s0[73]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U493 ( .a ({new_AGEMA_signal_4222, new_AGEMA_signal_4221, rd_I_n2478}), .b ({new_AGEMA_signal_4220, new_AGEMA_signal_4219, rd_I_n2480}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017]}), .c ({new_AGEMA_signal_5114, new_AGEMA_signal_5113, rd_I_n1534}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U482 ( .a ({new_AGEMA_signal_4228, new_AGEMA_signal_4227, rd_I_n2541}), .b ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, rd_I_n1528}), .c ({state_out_s2[234], state_out_s1[234], state_out_s0[234]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U481 ( .a ({new_AGEMA_signal_4226, new_AGEMA_signal_4225, rd_I_n2542}), .b ({new_AGEMA_signal_4224, new_AGEMA_signal_4223, rd_I_n2544}), .clk (clk), .r ({Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_5116, new_AGEMA_signal_5115, rd_I_n1528}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U477 ( .a ({new_AGEMA_signal_5118, new_AGEMA_signal_5117, rd_I_n1527}), .b ({new_AGEMA_signal_4230, new_AGEMA_signal_4229, rd_I_n2093}), .c ({state_out_s2[284], state_out_s1[284], state_out_s0[284]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U470 ( .a ({new_AGEMA_signal_4234, new_AGEMA_signal_4233, rd_I_n2095}), .b ({new_AGEMA_signal_4232, new_AGEMA_signal_4231, rd_I_n2092}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023]}), .c ({new_AGEMA_signal_5118, new_AGEMA_signal_5117, rd_I_n1527}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U459 ( .a ({new_AGEMA_signal_5122, new_AGEMA_signal_5121, rd_I_n2551}), .b ({new_AGEMA_signal_5120, new_AGEMA_signal_5119, rd_I_n1520}), .c ({state_out_s2[30], state_out_s1[30], state_out_s0[30]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U458 ( .a ({new_AGEMA_signal_4238, new_AGEMA_signal_4237, rd_I_n2552}), .b ({new_AGEMA_signal_4236, new_AGEMA_signal_4235, rd_I_n2554}), .clk (clk), .r ({Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_5120, new_AGEMA_signal_5119, rd_I_n1520}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U443 ( .a ({new_AGEMA_signal_5124, new_AGEMA_signal_5123, rd_I_n1513}), .b ({new_AGEMA_signal_4242, new_AGEMA_signal_4241, rd_I_n2424}), .c ({state_out_s2[191], state_out_s1[191], state_out_s0[191]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U441 ( .a ({new_AGEMA_signal_4246, new_AGEMA_signal_4245, rd_I_n2423}), .b ({new_AGEMA_signal_4244, new_AGEMA_signal_4243, rd_I_n2426}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029]}), .c ({new_AGEMA_signal_5124, new_AGEMA_signal_5123, rd_I_n1513}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U430 ( .a ({new_AGEMA_signal_5126, new_AGEMA_signal_5125, rd_I_n1508}), .b ({new_AGEMA_signal_4248, new_AGEMA_signal_4247, rd_I_n1825}), .c ({state_out_s2[337], state_out_s1[337], state_out_s0[337]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U425 ( .a ({new_AGEMA_signal_4252, new_AGEMA_signal_4251, rd_I_n1828}), .b ({new_AGEMA_signal_4250, new_AGEMA_signal_4249, rd_I_n1827}), .clk (clk), .r ({Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_5126, new_AGEMA_signal_5125, rd_I_n1508}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U415 ( .a ({new_AGEMA_signal_5128, new_AGEMA_signal_5127, rd_I_n1500}), .b ({new_AGEMA_signal_4254, new_AGEMA_signal_4253, rd_I_n2073}), .c ({state_out_s2[125], state_out_s1[125], state_out_s0[125]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U413 ( .a ({new_AGEMA_signal_4258, new_AGEMA_signal_4257, rd_I_n2076}), .b ({new_AGEMA_signal_4256, new_AGEMA_signal_4255, rd_I_n2074}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035]}), .c ({new_AGEMA_signal_5128, new_AGEMA_signal_5127, rd_I_n1500}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U407 ( .a ({new_AGEMA_signal_4394, new_AGEMA_signal_4393, rd_I_n1992}), .b ({new_AGEMA_signal_5130, new_AGEMA_signal_5129, rd_I_n1496}), .c ({state_out_s2[158], state_out_s1[158], state_out_s0[158]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U406 ( .a ({new_AGEMA_signal_4396, new_AGEMA_signal_4395, rd_I_n1991}), .b ({new_AGEMA_signal_4392, new_AGEMA_signal_4391, rd_I_n1994}), .clk (clk), .r ({Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_5130, new_AGEMA_signal_5129, rd_I_n1496}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U405 ( .a ({new_AGEMA_signal_4274, new_AGEMA_signal_4273, rd_I_n1707}), .b ({new_AGEMA_signal_5132, new_AGEMA_signal_5131, rd_I_n1495}), .c ({state_out_s2[304], state_out_s1[304], state_out_s0[304]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U404 ( .a ({new_AGEMA_signal_4272, new_AGEMA_signal_4271, rd_I_n1706}), .b ({new_AGEMA_signal_4276, new_AGEMA_signal_4275, rd_I_n1709}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041]}), .c ({new_AGEMA_signal_5132, new_AGEMA_signal_5131, rd_I_n1495}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U403 ( .a ({new_AGEMA_signal_4264, new_AGEMA_signal_4263, rd_I_n2314}), .b ({new_AGEMA_signal_5134, new_AGEMA_signal_5133, rd_I_n1494}), .c ({state_out_s2[69], state_out_s1[69], state_out_s0[69]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U402 ( .a ({new_AGEMA_signal_4262, new_AGEMA_signal_4261, rd_I_n2315}), .b ({new_AGEMA_signal_4260, new_AGEMA_signal_4259, rd_I_n2317}), .clk (clk), .r ({Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_5134, new_AGEMA_signal_5133, rd_I_n1494}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U398 ( .a ({new_AGEMA_signal_4340, new_AGEMA_signal_4339, rd_I_n2260}), .b ({new_AGEMA_signal_5136, new_AGEMA_signal_5135, rd_I_n1492}), .c ({state_out_s2[230], state_out_s1[230], state_out_s0[230]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U397 ( .a ({new_AGEMA_signal_4338, new_AGEMA_signal_4337, rd_I_n2259}), .b ({new_AGEMA_signal_4342, new_AGEMA_signal_4341, rd_I_n2262}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047]}), .c ({new_AGEMA_signal_5136, new_AGEMA_signal_5135, rd_I_n1492}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U396 ( .a ({new_AGEMA_signal_5138, new_AGEMA_signal_5137, rd_I_n1491}), .b ({new_AGEMA_signal_4266, new_AGEMA_signal_4265, rd_I_n2225}), .c ({state_out_s2[280], state_out_s1[280], state_out_s0[280]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U394 ( .a ({new_AGEMA_signal_4270, new_AGEMA_signal_4269, rd_I_n2228}), .b ({new_AGEMA_signal_4268, new_AGEMA_signal_4267, rd_I_n2226}), .clk (clk), .r ({Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_5138, new_AGEMA_signal_5137, rd_I_n1491}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U388 ( .a ({new_AGEMA_signal_5908, new_AGEMA_signal_5907, rd_I_n1488}), .b ({new_AGEMA_signal_4330, new_AGEMA_signal_4329, rd_I_n1682}), .c ({state_out_s2[113], state_out_s1[113], state_out_s0[113]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U387 ( .a ({new_AGEMA_signal_5140, new_AGEMA_signal_5139, rd_I_n1487}), .b ({new_AGEMA_signal_4328, new_AGEMA_signal_4327, rd_I_n1685}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053]}), .c ({new_AGEMA_signal_5908, new_AGEMA_signal_5907, rd_I_n1488}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U385 ( .a ({new_AGEMA_signal_5142, new_AGEMA_signal_5141, rd_I_n1486}), .b ({new_AGEMA_signal_4272, new_AGEMA_signal_4271, rd_I_n1706}), .c ({state_out_s2[104], state_out_s1[104], state_out_s0[104]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U383 ( .a ({new_AGEMA_signal_4276, new_AGEMA_signal_4275, rd_I_n1709}), .b ({new_AGEMA_signal_4274, new_AGEMA_signal_4273, rd_I_n1707}), .clk (clk), .r ({Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_5142, new_AGEMA_signal_5141, rd_I_n1486}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U377 ( .a ({new_AGEMA_signal_4282, new_AGEMA_signal_4281, rd_I_n2108}), .b ({new_AGEMA_signal_5912, new_AGEMA_signal_5911, rd_I_n1482}), .c ({state_out_s2[146], state_out_s1[146], state_out_s0[146]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U376 ( .a ({new_AGEMA_signal_5144, new_AGEMA_signal_5143, rd_I_n2110}), .b ({new_AGEMA_signal_4278, new_AGEMA_signal_4277, rd_I_n2107}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059]}), .c ({new_AGEMA_signal_5912, new_AGEMA_signal_5911, rd_I_n1482}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U370 ( .a ({new_AGEMA_signal_4288, new_AGEMA_signal_4287, rd_I_n2618}), .b ({new_AGEMA_signal_5914, new_AGEMA_signal_5913, rd_I_n1477}), .c ({state_out_s2[137], state_out_s1[137], state_out_s0[137]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U369 ( .a ({new_AGEMA_signal_5146, new_AGEMA_signal_5145, rd_I_n2620}), .b ({new_AGEMA_signal_4284, new_AGEMA_signal_4283, rd_I_n2617}), .clk (clk), .r ({Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_5914, new_AGEMA_signal_5913, rd_I_n1477}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U359 ( .a ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, rd_I_n1473}), .b ({new_AGEMA_signal_4290, new_AGEMA_signal_4289, rd_I_n2343}), .c ({state_out_s2[315], state_out_s1[315], state_out_s0[315]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U354 ( .a ({new_AGEMA_signal_4294, new_AGEMA_signal_4293, rd_I_n2346}), .b ({new_AGEMA_signal_4292, new_AGEMA_signal_4291, rd_I_n2344}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065]}), .c ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, rd_I_n1473}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U345 ( .a ({new_AGEMA_signal_5150, new_AGEMA_signal_5149, rd_I_n1466}), .b ({new_AGEMA_signal_4296, new_AGEMA_signal_4295, rd_I_n2348}), .c ({state_out_s2[292], state_out_s1[292], state_out_s0[292]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U343 ( .a ({new_AGEMA_signal_4300, new_AGEMA_signal_4299, rd_I_n2351}), .b ({new_AGEMA_signal_4298, new_AGEMA_signal_4297, rd_I_n2349}), .clk (clk), .r ({Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_5150, new_AGEMA_signal_5149, rd_I_n1466}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U334 ( .a ({new_AGEMA_signal_5152, new_AGEMA_signal_5151, rd_I_n1461}), .b ({new_AGEMA_signal_4302, new_AGEMA_signal_4301, rd_I_n2251}), .c ({state_out_s2[112], state_out_s1[112], state_out_s0[112]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U332 ( .a ({new_AGEMA_signal_4306, new_AGEMA_signal_4305, rd_I_n2250}), .b ({new_AGEMA_signal_4304, new_AGEMA_signal_4303, rd_I_n2253}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071]}), .c ({new_AGEMA_signal_5152, new_AGEMA_signal_5151, rd_I_n1461}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U326 ( .a ({new_AGEMA_signal_4448, new_AGEMA_signal_4447, rd_I_n1655}), .b ({new_AGEMA_signal_5154, new_AGEMA_signal_5153, rd_I_n1456}), .c ({state_out_s2[145], state_out_s1[145], state_out_s0[145]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U325 ( .a ({new_AGEMA_signal_4450, new_AGEMA_signal_4449, rd_I_n1654}), .b ({new_AGEMA_signal_4446, new_AGEMA_signal_4445, rd_I_n1657}), .clk (clk), .r ({Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_5154, new_AGEMA_signal_5153, rd_I_n1456}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U324 ( .a ({new_AGEMA_signal_5156, new_AGEMA_signal_5155, rd_I_n1455}), .b ({new_AGEMA_signal_4308, new_AGEMA_signal_4307, rd_I_n2458}), .c ({state_out_s2[291], state_out_s1[291], state_out_s0[291]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U322 ( .a ({new_AGEMA_signal_4312, new_AGEMA_signal_4311, rd_I_n2457}), .b ({new_AGEMA_signal_4310, new_AGEMA_signal_4309, rd_I_n2460}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077]}), .c ({new_AGEMA_signal_5156, new_AGEMA_signal_5155, rd_I_n1455}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U316 ( .a ({new_AGEMA_signal_4318, new_AGEMA_signal_4317, rd_I_n2068}), .b ({new_AGEMA_signal_5158, new_AGEMA_signal_5157, rd_I_n1452}), .c ({state_out_s2[102], state_out_s1[102], state_out_s0[102]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U315 ( .a ({new_AGEMA_signal_4316, new_AGEMA_signal_4315, rd_I_n2069}), .b ({new_AGEMA_signal_4314, new_AGEMA_signal_4313, rd_I_n2071}), .clk (clk), .r ({Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_5158, new_AGEMA_signal_5157, rd_I_n1452}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U305 ( .a ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, rd_I_n1446}), .b ({new_AGEMA_signal_4320, new_AGEMA_signal_4319, rd_I_n1856}), .c ({state_out_s2[135], state_out_s1[135], state_out_s0[135]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U303 ( .a ({new_AGEMA_signal_4324, new_AGEMA_signal_4323, rd_I_n1859}), .b ({new_AGEMA_signal_5160, new_AGEMA_signal_5159, rd_I_n1857}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083]}), .c ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, rd_I_n1446}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U297 ( .a ({new_AGEMA_signal_5162, new_AGEMA_signal_5161, rd_I_n1440}), .b ({new_AGEMA_signal_4326, new_AGEMA_signal_4325, rd_I_n1683}), .c ({state_out_s2[313], state_out_s1[313], state_out_s0[313]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U294 ( .a ({new_AGEMA_signal_4330, new_AGEMA_signal_4329, rd_I_n1682}), .b ({new_AGEMA_signal_4328, new_AGEMA_signal_4327, rd_I_n1685}), .clk (clk), .r ({Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_5162, new_AGEMA_signal_5161, rd_I_n1440}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U285 ( .a ({new_AGEMA_signal_5164, new_AGEMA_signal_5163, rd_I_n1433}), .b ({new_AGEMA_signal_4332, new_AGEMA_signal_4331, rd_I_n2284}), .c ({state_out_s2[122], state_out_s1[122], state_out_s0[122]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U283 ( .a ({new_AGEMA_signal_4336, new_AGEMA_signal_4335, rd_I_n2283}), .b ({new_AGEMA_signal_4334, new_AGEMA_signal_4333, rd_I_n2286}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089]}), .c ({new_AGEMA_signal_5164, new_AGEMA_signal_5163, rd_I_n1433}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U277 ( .a ({new_AGEMA_signal_4376, new_AGEMA_signal_4375, rd_I_n1999}), .b ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, rd_I_n1429}), .c ({state_out_s2[155], state_out_s1[155], state_out_s0[155]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U276 ( .a ({new_AGEMA_signal_4378, new_AGEMA_signal_4377, rd_I_n1998}), .b ({new_AGEMA_signal_4374, new_AGEMA_signal_4373, rd_I_n2001}), .clk (clk), .r ({Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, rd_I_n1429}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U275 ( .a ({new_AGEMA_signal_5168, new_AGEMA_signal_5167, rd_I_n1428}), .b ({new_AGEMA_signal_4338, new_AGEMA_signal_4337, rd_I_n2259}), .c ({state_out_s2[301], state_out_s1[301], state_out_s0[301]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U273 ( .a ({new_AGEMA_signal_4342, new_AGEMA_signal_4341, rd_I_n2262}), .b ({new_AGEMA_signal_4340, new_AGEMA_signal_4339, rd_I_n2260}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095]}), .c ({new_AGEMA_signal_5168, new_AGEMA_signal_5167, rd_I_n1428}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U267 ( .a ({new_AGEMA_signal_5170, new_AGEMA_signal_5169, rd_I_n1425}), .b ({new_AGEMA_signal_4344, new_AGEMA_signal_4343, rd_I_n2288}), .c ({state_out_s2[99], state_out_s1[99], state_out_s0[99]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U265 ( .a ({new_AGEMA_signal_4348, new_AGEMA_signal_4347, rd_I_n2287}), .b ({new_AGEMA_signal_4346, new_AGEMA_signal_4345, rd_I_n2290}), .clk (clk), .r ({Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_5170, new_AGEMA_signal_5169, rd_I_n1425}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U254 ( .a ({new_AGEMA_signal_4354, new_AGEMA_signal_4353, rd_I_n2375}), .b ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, rd_I_n1419}), .c ({state_out_s2[132], state_out_s1[132], state_out_s0[132]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U253 ( .a ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, rd_I_n2376}), .b ({new_AGEMA_signal_4350, new_AGEMA_signal_4349, rd_I_n2378}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101]}), .c ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, rd_I_n1419}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U242 ( .a ({new_AGEMA_signal_5174, new_AGEMA_signal_5173, rd_I_n1413}), .b ({new_AGEMA_signal_4356, new_AGEMA_signal_4355, rd_I_n1976}), .c ({state_out_s2[310], state_out_s1[310], state_out_s0[310]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U237 ( .a ({new_AGEMA_signal_4360, new_AGEMA_signal_4359, rd_I_n1978}), .b ({new_AGEMA_signal_4358, new_AGEMA_signal_4357, rd_I_n1979}), .clk (clk), .r ({Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_5174, new_AGEMA_signal_5173, rd_I_n1413}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U229 ( .a ({new_AGEMA_signal_4366, new_AGEMA_signal_4365, rd_I_n2291}), .b ({new_AGEMA_signal_5176, new_AGEMA_signal_5175, rd_I_n1408}), .c ({state_out_s2[15], state_out_s1[15], state_out_s0[15]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U228 ( .a ({new_AGEMA_signal_4364, new_AGEMA_signal_4363, rd_I_n2292}), .b ({new_AGEMA_signal_4362, new_AGEMA_signal_4361, rd_I_n2294}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107]}), .c ({new_AGEMA_signal_5176, new_AGEMA_signal_5175, rd_I_n1408}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U213 ( .a ({new_AGEMA_signal_4372, new_AGEMA_signal_4371, rd_I_n2266}), .b ({new_AGEMA_signal_5178, new_AGEMA_signal_5177, rd_I_n1401}), .c ({state_out_s2[176], state_out_s1[176], state_out_s0[176]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U212 ( .a ({new_AGEMA_signal_4370, new_AGEMA_signal_4369, rd_I_n2267}), .b ({new_AGEMA_signal_4368, new_AGEMA_signal_4367, rd_I_n2269}), .clk (clk), .r ({Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_5178, new_AGEMA_signal_5177, rd_I_n1401}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U198 ( .a ({new_AGEMA_signal_4378, new_AGEMA_signal_4377, rd_I_n1998}), .b ({new_AGEMA_signal_5180, new_AGEMA_signal_5179, rd_I_n1396}), .c ({state_out_s2[322], state_out_s1[322], state_out_s0[322]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U197 ( .a ({new_AGEMA_signal_4376, new_AGEMA_signal_4375, rd_I_n1999}), .b ({new_AGEMA_signal_4374, new_AGEMA_signal_4373, rd_I_n2001}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113]}), .c ({new_AGEMA_signal_5180, new_AGEMA_signal_5179, rd_I_n1396}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U182 ( .a ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, rd_I_n1390}), .b ({new_AGEMA_signal_4380, new_AGEMA_signal_4379, rd_I_n1777}), .c ({state_out_s2[18], state_out_s1[18], state_out_s0[18]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U179 ( .a ({new_AGEMA_signal_4384, new_AGEMA_signal_4383, rd_I_n1780}), .b ({new_AGEMA_signal_4382, new_AGEMA_signal_4381, rd_I_n1778}), .clk (clk), .r ({Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_5182, new_AGEMA_signal_5181, rd_I_n1390}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U168 ( .a ({new_AGEMA_signal_4390, new_AGEMA_signal_4389, rd_I_n2405}), .b ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, rd_I_n1383}), .c ({state_out_s2[179], state_out_s1[179], state_out_s0[179]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U167 ( .a ({new_AGEMA_signal_4388, new_AGEMA_signal_4387, rd_I_n2406}), .b ({new_AGEMA_signal_4386, new_AGEMA_signal_4385, rd_I_n2408}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119]}), .c ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, rd_I_n1383}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U153 ( .a ({new_AGEMA_signal_4396, new_AGEMA_signal_4395, rd_I_n1991}), .b ({new_AGEMA_signal_5186, new_AGEMA_signal_5185, rd_I_n1378}), .c ({state_out_s2[325], state_out_s1[325], state_out_s0[325]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U152 ( .a ({new_AGEMA_signal_4394, new_AGEMA_signal_4393, rd_I_n1992}), .b ({new_AGEMA_signal_4392, new_AGEMA_signal_4391, rd_I_n1994}), .clk (clk), .r ({Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_5186, new_AGEMA_signal_5185, rd_I_n1378}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U132 ( .a ({new_AGEMA_signal_5188, new_AGEMA_signal_5187, rd_I_n1370}), .b ({new_AGEMA_signal_4398, new_AGEMA_signal_4397, rd_I_n2112}), .c ({state_out_s2[98], state_out_s1[98], state_out_s0[98]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U130 ( .a ({new_AGEMA_signal_4402, new_AGEMA_signal_4401, rd_I_n2115}), .b ({new_AGEMA_signal_4400, new_AGEMA_signal_4399, rd_I_n2113}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125]}), .c ({new_AGEMA_signal_5188, new_AGEMA_signal_5187, rd_I_n1370}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U121 ( .a ({new_AGEMA_signal_4408, new_AGEMA_signal_4407, rd_I_n2495}), .b ({new_AGEMA_signal_5190, new_AGEMA_signal_5189, rd_I_n1364}), .c ({state_out_s2[131], state_out_s1[131], state_out_s0[131]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U120 ( .a ({new_AGEMA_signal_4406, new_AGEMA_signal_4405, rd_I_n2496}), .b ({new_AGEMA_signal_4404, new_AGEMA_signal_4403, rd_I_n2498}), .clk (clk), .r ({Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_5190, new_AGEMA_signal_5189, rd_I_n1364}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U109 ( .a ({new_AGEMA_signal_5192, new_AGEMA_signal_5191, rd_I_n1358}), .b ({new_AGEMA_signal_4410, new_AGEMA_signal_4409, rd_I_n1815}), .c ({state_out_s2[309], state_out_s1[309], state_out_s0[309]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U104 ( .a ({new_AGEMA_signal_4414, new_AGEMA_signal_4413, rd_I_n1818}), .b ({new_AGEMA_signal_4412, new_AGEMA_signal_4411, rd_I_n1816}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131]}), .c ({new_AGEMA_signal_5192, new_AGEMA_signal_5191, rd_I_n1358}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U95 ( .a ({new_AGEMA_signal_5194, new_AGEMA_signal_5193, rd_I_n1351}), .b ({new_AGEMA_signal_4416, new_AGEMA_signal_4415, rd_I_n2220}), .c ({state_out_s2[121], state_out_s1[121], state_out_s0[121]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U93 ( .a ({new_AGEMA_signal_4420, new_AGEMA_signal_4419, rd_I_n2223}), .b ({new_AGEMA_signal_4418, new_AGEMA_signal_4417, rd_I_n2221}), .clk (clk), .r ({Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_5194, new_AGEMA_signal_5193, rd_I_n1351}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U82 ( .a ({new_AGEMA_signal_4426, new_AGEMA_signal_4425, rd_I_n2490}), .b ({new_AGEMA_signal_5196, new_AGEMA_signal_5195, rd_I_n1345}), .c ({state_out_s2[154], state_out_s1[154], state_out_s0[154]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U81 ( .a ({new_AGEMA_signal_4424, new_AGEMA_signal_4423, rd_I_n2491}), .b ({new_AGEMA_signal_4422, new_AGEMA_signal_4421, rd_I_n2493}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137]}), .c ({new_AGEMA_signal_5196, new_AGEMA_signal_5195, rd_I_n1345}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U70 ( .a ({new_AGEMA_signal_5198, new_AGEMA_signal_5197, rd_I_n1339}), .b ({new_AGEMA_signal_4428, new_AGEMA_signal_4427, rd_I_n2454}), .c ({state_out_s2[300], state_out_s1[300], state_out_s0[300]}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U65 ( .a ({new_AGEMA_signal_4432, new_AGEMA_signal_4431, rd_I_n2456}), .b ({new_AGEMA_signal_4430, new_AGEMA_signal_4429, rd_I_n2453}), .clk (clk), .r ({Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_5198, new_AGEMA_signal_5197, rd_I_n1339}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U52 ( .a ({new_AGEMA_signal_4438, new_AGEMA_signal_4437, rd_I_n2254}), .b ({new_AGEMA_signal_5200, new_AGEMA_signal_5199, rd_I_n1332}), .c ({state_out_s2[5], state_out_s1[5], state_out_s0[5]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U51 ( .a ({new_AGEMA_signal_4436, new_AGEMA_signal_4435, rd_I_n2255}), .b ({new_AGEMA_signal_4434, new_AGEMA_signal_4433, rd_I_n2257}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143]}), .c ({new_AGEMA_signal_5200, new_AGEMA_signal_5199, rd_I_n1332}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U36 ( .a ({new_AGEMA_signal_4444, new_AGEMA_signal_4443, rd_I_n2324}), .b ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, rd_I_n1325}), .c ({state_out_s2[166], state_out_s1[166], state_out_s0[166]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U35 ( .a ({new_AGEMA_signal_4442, new_AGEMA_signal_4441, rd_I_n2326}), .b ({new_AGEMA_signal_4440, new_AGEMA_signal_4439, rd_I_n2323}), .clk (clk), .r ({Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, rd_I_n1325}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U21 ( .a ({new_AGEMA_signal_4450, new_AGEMA_signal_4449, rd_I_n1654}), .b ({new_AGEMA_signal_5204, new_AGEMA_signal_5203, rd_I_n1320}), .c ({state_out_s2[344], state_out_s1[344], state_out_s0[344]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) rd_I_U20 ( .a ({new_AGEMA_signal_4448, new_AGEMA_signal_4447, rd_I_n1655}), .b ({new_AGEMA_signal_4446, new_AGEMA_signal_4445, rd_I_n1657}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149]}), .c ({new_AGEMA_signal_5204, new_AGEMA_signal_5203, rd_I_n1320}) ) ;

endmodule
