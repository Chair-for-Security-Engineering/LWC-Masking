/* modified netlist. Source: module elephant_perm in file ./test/elephant_perm.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module elephant_perm_HPC2_ClockGating_d3 (input0_s0, lfsr, rev_lfsr, clk, input0_s1, input0_s2, input0_s3, Fresh, /*rst,*/ output0_s0, output0_s1, output0_s2, output0_s3/*, Synch*/);
    input [159:0] input0_s0 ;
    input [6:0] lfsr ;
    input [6:0] rev_lfsr ;
    input clk ;
    input [159:0] input0_s1 ;
    input [159:0] input0_s2 ;
    input [159:0] input0_s3 ;
    //input rst ;
    input [1679:0] Fresh ;
    output [159:0] output0_s0 ;
    output [159:0] output0_s1 ;
    output [159:0] output0_s2 ;
    output [159:0] output0_s3 ;
    //output Synch ;
    wire input_array_6 ;
    wire input_array_5 ;
    wire input_array_4 ;
    wire input_array_3 ;
    wire input_array_2 ;
    wire input_array_1 ;
    wire input_array_0 ;
    wire sbox_inst_39_n20 ;
    wire sbox_inst_39_n19 ;
    wire sbox_inst_39_n18 ;
    wire sbox_inst_39_n17 ;
    wire sbox_inst_39_n16 ;
    wire sbox_inst_39_n15 ;
    wire sbox_inst_39_n14 ;
    wire sbox_inst_39_n13 ;
    wire sbox_inst_39_n12 ;
    wire sbox_inst_39_n11 ;
    wire sbox_inst_39_T6 ;
    wire sbox_inst_39_L0 ;
    wire sbox_inst_39_T5 ;
    wire sbox_inst_39_T4 ;
    wire sbox_inst_39_T3 ;
    wire sbox_inst_39_T2 ;
    wire sbox_inst_39_T1 ;
    wire sbox_inst_39_T0 ;
    wire sbox_inst_38_n20 ;
    wire sbox_inst_38_n19 ;
    wire sbox_inst_38_n18 ;
    wire sbox_inst_38_n17 ;
    wire sbox_inst_38_n16 ;
    wire sbox_inst_38_n15 ;
    wire sbox_inst_38_n14 ;
    wire sbox_inst_38_n13 ;
    wire sbox_inst_38_n12 ;
    wire sbox_inst_38_n11 ;
    wire sbox_inst_38_T6 ;
    wire sbox_inst_38_L0 ;
    wire sbox_inst_38_T5 ;
    wire sbox_inst_38_T4 ;
    wire sbox_inst_38_T3 ;
    wire sbox_inst_38_T2 ;
    wire sbox_inst_38_T1 ;
    wire sbox_inst_38_T0 ;
    wire sbox_inst_37_n20 ;
    wire sbox_inst_37_n19 ;
    wire sbox_inst_37_n18 ;
    wire sbox_inst_37_n17 ;
    wire sbox_inst_37_n16 ;
    wire sbox_inst_37_n15 ;
    wire sbox_inst_37_n14 ;
    wire sbox_inst_37_n13 ;
    wire sbox_inst_37_n12 ;
    wire sbox_inst_37_n11 ;
    wire sbox_inst_37_T6 ;
    wire sbox_inst_37_L0 ;
    wire sbox_inst_37_T5 ;
    wire sbox_inst_37_T4 ;
    wire sbox_inst_37_T3 ;
    wire sbox_inst_37_T2 ;
    wire sbox_inst_37_T1 ;
    wire sbox_inst_37_T0 ;
    wire sbox_inst_36_n20 ;
    wire sbox_inst_36_n19 ;
    wire sbox_inst_36_n18 ;
    wire sbox_inst_36_n17 ;
    wire sbox_inst_36_n16 ;
    wire sbox_inst_36_n15 ;
    wire sbox_inst_36_n14 ;
    wire sbox_inst_36_n13 ;
    wire sbox_inst_36_n12 ;
    wire sbox_inst_36_n11 ;
    wire sbox_inst_36_T6 ;
    wire sbox_inst_36_L0 ;
    wire sbox_inst_36_T5 ;
    wire sbox_inst_36_T4 ;
    wire sbox_inst_36_T3 ;
    wire sbox_inst_36_T2 ;
    wire sbox_inst_36_T1 ;
    wire sbox_inst_36_T0 ;
    wire sbox_inst_35_n20 ;
    wire sbox_inst_35_n19 ;
    wire sbox_inst_35_n18 ;
    wire sbox_inst_35_n17 ;
    wire sbox_inst_35_n16 ;
    wire sbox_inst_35_n15 ;
    wire sbox_inst_35_n14 ;
    wire sbox_inst_35_n13 ;
    wire sbox_inst_35_n12 ;
    wire sbox_inst_35_n11 ;
    wire sbox_inst_35_T6 ;
    wire sbox_inst_35_L0 ;
    wire sbox_inst_35_T5 ;
    wire sbox_inst_35_T4 ;
    wire sbox_inst_35_T3 ;
    wire sbox_inst_35_T2 ;
    wire sbox_inst_35_T1 ;
    wire sbox_inst_35_T0 ;
    wire sbox_inst_34_n20 ;
    wire sbox_inst_34_n19 ;
    wire sbox_inst_34_n18 ;
    wire sbox_inst_34_n17 ;
    wire sbox_inst_34_n16 ;
    wire sbox_inst_34_n15 ;
    wire sbox_inst_34_n14 ;
    wire sbox_inst_34_n13 ;
    wire sbox_inst_34_n12 ;
    wire sbox_inst_34_n11 ;
    wire sbox_inst_34_T6 ;
    wire sbox_inst_34_L0 ;
    wire sbox_inst_34_T5 ;
    wire sbox_inst_34_T4 ;
    wire sbox_inst_34_T3 ;
    wire sbox_inst_34_T2 ;
    wire sbox_inst_34_T1 ;
    wire sbox_inst_34_T0 ;
    wire sbox_inst_33_n20 ;
    wire sbox_inst_33_n19 ;
    wire sbox_inst_33_n18 ;
    wire sbox_inst_33_n17 ;
    wire sbox_inst_33_n16 ;
    wire sbox_inst_33_n15 ;
    wire sbox_inst_33_n14 ;
    wire sbox_inst_33_n13 ;
    wire sbox_inst_33_n12 ;
    wire sbox_inst_33_n11 ;
    wire sbox_inst_33_T6 ;
    wire sbox_inst_33_L0 ;
    wire sbox_inst_33_T5 ;
    wire sbox_inst_33_T4 ;
    wire sbox_inst_33_T3 ;
    wire sbox_inst_33_T2 ;
    wire sbox_inst_33_T1 ;
    wire sbox_inst_33_T0 ;
    wire sbox_inst_32_n20 ;
    wire sbox_inst_32_n19 ;
    wire sbox_inst_32_n18 ;
    wire sbox_inst_32_n17 ;
    wire sbox_inst_32_n16 ;
    wire sbox_inst_32_n15 ;
    wire sbox_inst_32_n14 ;
    wire sbox_inst_32_n13 ;
    wire sbox_inst_32_n12 ;
    wire sbox_inst_32_n11 ;
    wire sbox_inst_32_T6 ;
    wire sbox_inst_32_L0 ;
    wire sbox_inst_32_T5 ;
    wire sbox_inst_32_T4 ;
    wire sbox_inst_32_T3 ;
    wire sbox_inst_32_T2 ;
    wire sbox_inst_32_T1 ;
    wire sbox_inst_32_T0 ;
    wire sbox_inst_31_n20 ;
    wire sbox_inst_31_n19 ;
    wire sbox_inst_31_n18 ;
    wire sbox_inst_31_n17 ;
    wire sbox_inst_31_n16 ;
    wire sbox_inst_31_n15 ;
    wire sbox_inst_31_n14 ;
    wire sbox_inst_31_n13 ;
    wire sbox_inst_31_n12 ;
    wire sbox_inst_31_n11 ;
    wire sbox_inst_31_T6 ;
    wire sbox_inst_31_L0 ;
    wire sbox_inst_31_T5 ;
    wire sbox_inst_31_T4 ;
    wire sbox_inst_31_T3 ;
    wire sbox_inst_31_T2 ;
    wire sbox_inst_31_T1 ;
    wire sbox_inst_31_T0 ;
    wire sbox_inst_30_n20 ;
    wire sbox_inst_30_n19 ;
    wire sbox_inst_30_n18 ;
    wire sbox_inst_30_n17 ;
    wire sbox_inst_30_n16 ;
    wire sbox_inst_30_n15 ;
    wire sbox_inst_30_n14 ;
    wire sbox_inst_30_n13 ;
    wire sbox_inst_30_n12 ;
    wire sbox_inst_30_n11 ;
    wire sbox_inst_30_T6 ;
    wire sbox_inst_30_L0 ;
    wire sbox_inst_30_T5 ;
    wire sbox_inst_30_T4 ;
    wire sbox_inst_30_T3 ;
    wire sbox_inst_30_T2 ;
    wire sbox_inst_30_T1 ;
    wire sbox_inst_30_T0 ;
    wire sbox_inst_29_n20 ;
    wire sbox_inst_29_n19 ;
    wire sbox_inst_29_n18 ;
    wire sbox_inst_29_n17 ;
    wire sbox_inst_29_n16 ;
    wire sbox_inst_29_n15 ;
    wire sbox_inst_29_n14 ;
    wire sbox_inst_29_n13 ;
    wire sbox_inst_29_n12 ;
    wire sbox_inst_29_n11 ;
    wire sbox_inst_29_T6 ;
    wire sbox_inst_29_L0 ;
    wire sbox_inst_29_T5 ;
    wire sbox_inst_29_T4 ;
    wire sbox_inst_29_T3 ;
    wire sbox_inst_29_T2 ;
    wire sbox_inst_29_T1 ;
    wire sbox_inst_29_T0 ;
    wire sbox_inst_28_n20 ;
    wire sbox_inst_28_n19 ;
    wire sbox_inst_28_n18 ;
    wire sbox_inst_28_n17 ;
    wire sbox_inst_28_n16 ;
    wire sbox_inst_28_n15 ;
    wire sbox_inst_28_n14 ;
    wire sbox_inst_28_n13 ;
    wire sbox_inst_28_n12 ;
    wire sbox_inst_28_n11 ;
    wire sbox_inst_28_T6 ;
    wire sbox_inst_28_L0 ;
    wire sbox_inst_28_T5 ;
    wire sbox_inst_28_T4 ;
    wire sbox_inst_28_T3 ;
    wire sbox_inst_28_T2 ;
    wire sbox_inst_28_T1 ;
    wire sbox_inst_28_T0 ;
    wire sbox_inst_27_n20 ;
    wire sbox_inst_27_n19 ;
    wire sbox_inst_27_n18 ;
    wire sbox_inst_27_n17 ;
    wire sbox_inst_27_n16 ;
    wire sbox_inst_27_n15 ;
    wire sbox_inst_27_n14 ;
    wire sbox_inst_27_n13 ;
    wire sbox_inst_27_n12 ;
    wire sbox_inst_27_n11 ;
    wire sbox_inst_27_T6 ;
    wire sbox_inst_27_L0 ;
    wire sbox_inst_27_T5 ;
    wire sbox_inst_27_T4 ;
    wire sbox_inst_27_T3 ;
    wire sbox_inst_27_T2 ;
    wire sbox_inst_27_T1 ;
    wire sbox_inst_27_T0 ;
    wire sbox_inst_26_n20 ;
    wire sbox_inst_26_n19 ;
    wire sbox_inst_26_n18 ;
    wire sbox_inst_26_n17 ;
    wire sbox_inst_26_n16 ;
    wire sbox_inst_26_n15 ;
    wire sbox_inst_26_n14 ;
    wire sbox_inst_26_n13 ;
    wire sbox_inst_26_n12 ;
    wire sbox_inst_26_n11 ;
    wire sbox_inst_26_T6 ;
    wire sbox_inst_26_L0 ;
    wire sbox_inst_26_T5 ;
    wire sbox_inst_26_T4 ;
    wire sbox_inst_26_T3 ;
    wire sbox_inst_26_T2 ;
    wire sbox_inst_26_T1 ;
    wire sbox_inst_26_T0 ;
    wire sbox_inst_25_n20 ;
    wire sbox_inst_25_n19 ;
    wire sbox_inst_25_n18 ;
    wire sbox_inst_25_n17 ;
    wire sbox_inst_25_n16 ;
    wire sbox_inst_25_n15 ;
    wire sbox_inst_25_n14 ;
    wire sbox_inst_25_n13 ;
    wire sbox_inst_25_n12 ;
    wire sbox_inst_25_n11 ;
    wire sbox_inst_25_T6 ;
    wire sbox_inst_25_L0 ;
    wire sbox_inst_25_T5 ;
    wire sbox_inst_25_T4 ;
    wire sbox_inst_25_T3 ;
    wire sbox_inst_25_T2 ;
    wire sbox_inst_25_T1 ;
    wire sbox_inst_25_T0 ;
    wire sbox_inst_24_n20 ;
    wire sbox_inst_24_n19 ;
    wire sbox_inst_24_n18 ;
    wire sbox_inst_24_n17 ;
    wire sbox_inst_24_n16 ;
    wire sbox_inst_24_n15 ;
    wire sbox_inst_24_n14 ;
    wire sbox_inst_24_n13 ;
    wire sbox_inst_24_n12 ;
    wire sbox_inst_24_n11 ;
    wire sbox_inst_24_T6 ;
    wire sbox_inst_24_L0 ;
    wire sbox_inst_24_T5 ;
    wire sbox_inst_24_T4 ;
    wire sbox_inst_24_T3 ;
    wire sbox_inst_24_T2 ;
    wire sbox_inst_24_T1 ;
    wire sbox_inst_24_T0 ;
    wire sbox_inst_23_n20 ;
    wire sbox_inst_23_n19 ;
    wire sbox_inst_23_n18 ;
    wire sbox_inst_23_n17 ;
    wire sbox_inst_23_n16 ;
    wire sbox_inst_23_n15 ;
    wire sbox_inst_23_n14 ;
    wire sbox_inst_23_n13 ;
    wire sbox_inst_23_n12 ;
    wire sbox_inst_23_n11 ;
    wire sbox_inst_23_T6 ;
    wire sbox_inst_23_L0 ;
    wire sbox_inst_23_T5 ;
    wire sbox_inst_23_T4 ;
    wire sbox_inst_23_T3 ;
    wire sbox_inst_23_T2 ;
    wire sbox_inst_23_T1 ;
    wire sbox_inst_23_T0 ;
    wire sbox_inst_22_n20 ;
    wire sbox_inst_22_n19 ;
    wire sbox_inst_22_n18 ;
    wire sbox_inst_22_n17 ;
    wire sbox_inst_22_n16 ;
    wire sbox_inst_22_n15 ;
    wire sbox_inst_22_n14 ;
    wire sbox_inst_22_n13 ;
    wire sbox_inst_22_n12 ;
    wire sbox_inst_22_n11 ;
    wire sbox_inst_22_T6 ;
    wire sbox_inst_22_L0 ;
    wire sbox_inst_22_T5 ;
    wire sbox_inst_22_T4 ;
    wire sbox_inst_22_T3 ;
    wire sbox_inst_22_T2 ;
    wire sbox_inst_22_T1 ;
    wire sbox_inst_22_T0 ;
    wire sbox_inst_21_n20 ;
    wire sbox_inst_21_n19 ;
    wire sbox_inst_21_n18 ;
    wire sbox_inst_21_n17 ;
    wire sbox_inst_21_n16 ;
    wire sbox_inst_21_n15 ;
    wire sbox_inst_21_n14 ;
    wire sbox_inst_21_n13 ;
    wire sbox_inst_21_n12 ;
    wire sbox_inst_21_n11 ;
    wire sbox_inst_21_T6 ;
    wire sbox_inst_21_L0 ;
    wire sbox_inst_21_T5 ;
    wire sbox_inst_21_T4 ;
    wire sbox_inst_21_T3 ;
    wire sbox_inst_21_T2 ;
    wire sbox_inst_21_T1 ;
    wire sbox_inst_21_T0 ;
    wire sbox_inst_20_n20 ;
    wire sbox_inst_20_n19 ;
    wire sbox_inst_20_n18 ;
    wire sbox_inst_20_n17 ;
    wire sbox_inst_20_n16 ;
    wire sbox_inst_20_n15 ;
    wire sbox_inst_20_n14 ;
    wire sbox_inst_20_n13 ;
    wire sbox_inst_20_n12 ;
    wire sbox_inst_20_n11 ;
    wire sbox_inst_20_T6 ;
    wire sbox_inst_20_L0 ;
    wire sbox_inst_20_T5 ;
    wire sbox_inst_20_T4 ;
    wire sbox_inst_20_T3 ;
    wire sbox_inst_20_T2 ;
    wire sbox_inst_20_T1 ;
    wire sbox_inst_20_T0 ;
    wire sbox_inst_19_n20 ;
    wire sbox_inst_19_n19 ;
    wire sbox_inst_19_n18 ;
    wire sbox_inst_19_n17 ;
    wire sbox_inst_19_n16 ;
    wire sbox_inst_19_n15 ;
    wire sbox_inst_19_n14 ;
    wire sbox_inst_19_n13 ;
    wire sbox_inst_19_n12 ;
    wire sbox_inst_19_n11 ;
    wire sbox_inst_19_T6 ;
    wire sbox_inst_19_L0 ;
    wire sbox_inst_19_T5 ;
    wire sbox_inst_19_T4 ;
    wire sbox_inst_19_T3 ;
    wire sbox_inst_19_T2 ;
    wire sbox_inst_19_T1 ;
    wire sbox_inst_19_T0 ;
    wire sbox_inst_18_n20 ;
    wire sbox_inst_18_n19 ;
    wire sbox_inst_18_n18 ;
    wire sbox_inst_18_n17 ;
    wire sbox_inst_18_n16 ;
    wire sbox_inst_18_n15 ;
    wire sbox_inst_18_n14 ;
    wire sbox_inst_18_n13 ;
    wire sbox_inst_18_n12 ;
    wire sbox_inst_18_n11 ;
    wire sbox_inst_18_T6 ;
    wire sbox_inst_18_L0 ;
    wire sbox_inst_18_T5 ;
    wire sbox_inst_18_T4 ;
    wire sbox_inst_18_T3 ;
    wire sbox_inst_18_T2 ;
    wire sbox_inst_18_T1 ;
    wire sbox_inst_18_T0 ;
    wire sbox_inst_17_n20 ;
    wire sbox_inst_17_n19 ;
    wire sbox_inst_17_n18 ;
    wire sbox_inst_17_n17 ;
    wire sbox_inst_17_n16 ;
    wire sbox_inst_17_n15 ;
    wire sbox_inst_17_n14 ;
    wire sbox_inst_17_n13 ;
    wire sbox_inst_17_n12 ;
    wire sbox_inst_17_n11 ;
    wire sbox_inst_17_T6 ;
    wire sbox_inst_17_L0 ;
    wire sbox_inst_17_T5 ;
    wire sbox_inst_17_T4 ;
    wire sbox_inst_17_T3 ;
    wire sbox_inst_17_T2 ;
    wire sbox_inst_17_T1 ;
    wire sbox_inst_17_T0 ;
    wire sbox_inst_16_n20 ;
    wire sbox_inst_16_n19 ;
    wire sbox_inst_16_n18 ;
    wire sbox_inst_16_n17 ;
    wire sbox_inst_16_n16 ;
    wire sbox_inst_16_n15 ;
    wire sbox_inst_16_n14 ;
    wire sbox_inst_16_n13 ;
    wire sbox_inst_16_n12 ;
    wire sbox_inst_16_n11 ;
    wire sbox_inst_16_T6 ;
    wire sbox_inst_16_L0 ;
    wire sbox_inst_16_T5 ;
    wire sbox_inst_16_T4 ;
    wire sbox_inst_16_T3 ;
    wire sbox_inst_16_T2 ;
    wire sbox_inst_16_T1 ;
    wire sbox_inst_16_T0 ;
    wire sbox_inst_15_n20 ;
    wire sbox_inst_15_n19 ;
    wire sbox_inst_15_n18 ;
    wire sbox_inst_15_n17 ;
    wire sbox_inst_15_n16 ;
    wire sbox_inst_15_n15 ;
    wire sbox_inst_15_n14 ;
    wire sbox_inst_15_n13 ;
    wire sbox_inst_15_n12 ;
    wire sbox_inst_15_n11 ;
    wire sbox_inst_15_T6 ;
    wire sbox_inst_15_L0 ;
    wire sbox_inst_15_T5 ;
    wire sbox_inst_15_T4 ;
    wire sbox_inst_15_T3 ;
    wire sbox_inst_15_T2 ;
    wire sbox_inst_15_T1 ;
    wire sbox_inst_15_T0 ;
    wire sbox_inst_14_n20 ;
    wire sbox_inst_14_n19 ;
    wire sbox_inst_14_n18 ;
    wire sbox_inst_14_n17 ;
    wire sbox_inst_14_n16 ;
    wire sbox_inst_14_n15 ;
    wire sbox_inst_14_n14 ;
    wire sbox_inst_14_n13 ;
    wire sbox_inst_14_n12 ;
    wire sbox_inst_14_n11 ;
    wire sbox_inst_14_T6 ;
    wire sbox_inst_14_L0 ;
    wire sbox_inst_14_T5 ;
    wire sbox_inst_14_T4 ;
    wire sbox_inst_14_T3 ;
    wire sbox_inst_14_T2 ;
    wire sbox_inst_14_T1 ;
    wire sbox_inst_14_T0 ;
    wire sbox_inst_13_n20 ;
    wire sbox_inst_13_n19 ;
    wire sbox_inst_13_n18 ;
    wire sbox_inst_13_n17 ;
    wire sbox_inst_13_n16 ;
    wire sbox_inst_13_n15 ;
    wire sbox_inst_13_n14 ;
    wire sbox_inst_13_n13 ;
    wire sbox_inst_13_n12 ;
    wire sbox_inst_13_n11 ;
    wire sbox_inst_13_T6 ;
    wire sbox_inst_13_L0 ;
    wire sbox_inst_13_T5 ;
    wire sbox_inst_13_T4 ;
    wire sbox_inst_13_T3 ;
    wire sbox_inst_13_T2 ;
    wire sbox_inst_13_T1 ;
    wire sbox_inst_13_T0 ;
    wire sbox_inst_12_n20 ;
    wire sbox_inst_12_n19 ;
    wire sbox_inst_12_n18 ;
    wire sbox_inst_12_n17 ;
    wire sbox_inst_12_n16 ;
    wire sbox_inst_12_n15 ;
    wire sbox_inst_12_n14 ;
    wire sbox_inst_12_n13 ;
    wire sbox_inst_12_n12 ;
    wire sbox_inst_12_n11 ;
    wire sbox_inst_12_T6 ;
    wire sbox_inst_12_L0 ;
    wire sbox_inst_12_T5 ;
    wire sbox_inst_12_T4 ;
    wire sbox_inst_12_T3 ;
    wire sbox_inst_12_T2 ;
    wire sbox_inst_12_T1 ;
    wire sbox_inst_12_T0 ;
    wire sbox_inst_11_n20 ;
    wire sbox_inst_11_n19 ;
    wire sbox_inst_11_n18 ;
    wire sbox_inst_11_n17 ;
    wire sbox_inst_11_n16 ;
    wire sbox_inst_11_n15 ;
    wire sbox_inst_11_n14 ;
    wire sbox_inst_11_n13 ;
    wire sbox_inst_11_n12 ;
    wire sbox_inst_11_n11 ;
    wire sbox_inst_11_T6 ;
    wire sbox_inst_11_L0 ;
    wire sbox_inst_11_T5 ;
    wire sbox_inst_11_T4 ;
    wire sbox_inst_11_T3 ;
    wire sbox_inst_11_T2 ;
    wire sbox_inst_11_T1 ;
    wire sbox_inst_11_T0 ;
    wire sbox_inst_10_n20 ;
    wire sbox_inst_10_n19 ;
    wire sbox_inst_10_n18 ;
    wire sbox_inst_10_n17 ;
    wire sbox_inst_10_n16 ;
    wire sbox_inst_10_n15 ;
    wire sbox_inst_10_n14 ;
    wire sbox_inst_10_n13 ;
    wire sbox_inst_10_n12 ;
    wire sbox_inst_10_n11 ;
    wire sbox_inst_10_T6 ;
    wire sbox_inst_10_L0 ;
    wire sbox_inst_10_T5 ;
    wire sbox_inst_10_T4 ;
    wire sbox_inst_10_T3 ;
    wire sbox_inst_10_T2 ;
    wire sbox_inst_10_T1 ;
    wire sbox_inst_10_T0 ;
    wire sbox_inst_9_n20 ;
    wire sbox_inst_9_n19 ;
    wire sbox_inst_9_n18 ;
    wire sbox_inst_9_n17 ;
    wire sbox_inst_9_n16 ;
    wire sbox_inst_9_n15 ;
    wire sbox_inst_9_n14 ;
    wire sbox_inst_9_n13 ;
    wire sbox_inst_9_n12 ;
    wire sbox_inst_9_n11 ;
    wire sbox_inst_9_T6 ;
    wire sbox_inst_9_L0 ;
    wire sbox_inst_9_T5 ;
    wire sbox_inst_9_T4 ;
    wire sbox_inst_9_T3 ;
    wire sbox_inst_9_T2 ;
    wire sbox_inst_9_T1 ;
    wire sbox_inst_9_T0 ;
    wire sbox_inst_8_n20 ;
    wire sbox_inst_8_n19 ;
    wire sbox_inst_8_n18 ;
    wire sbox_inst_8_n17 ;
    wire sbox_inst_8_n16 ;
    wire sbox_inst_8_n15 ;
    wire sbox_inst_8_n14 ;
    wire sbox_inst_8_n13 ;
    wire sbox_inst_8_n12 ;
    wire sbox_inst_8_n11 ;
    wire sbox_inst_8_T6 ;
    wire sbox_inst_8_L0 ;
    wire sbox_inst_8_T5 ;
    wire sbox_inst_8_T4 ;
    wire sbox_inst_8_T3 ;
    wire sbox_inst_8_T2 ;
    wire sbox_inst_8_T1 ;
    wire sbox_inst_8_T0 ;
    wire sbox_inst_7_n20 ;
    wire sbox_inst_7_n19 ;
    wire sbox_inst_7_n18 ;
    wire sbox_inst_7_n17 ;
    wire sbox_inst_7_n16 ;
    wire sbox_inst_7_n15 ;
    wire sbox_inst_7_n14 ;
    wire sbox_inst_7_n13 ;
    wire sbox_inst_7_n12 ;
    wire sbox_inst_7_n11 ;
    wire sbox_inst_7_T6 ;
    wire sbox_inst_7_L0 ;
    wire sbox_inst_7_T5 ;
    wire sbox_inst_7_T4 ;
    wire sbox_inst_7_T3 ;
    wire sbox_inst_7_T2 ;
    wire sbox_inst_7_T1 ;
    wire sbox_inst_7_T0 ;
    wire sbox_inst_6_n20 ;
    wire sbox_inst_6_n19 ;
    wire sbox_inst_6_n18 ;
    wire sbox_inst_6_n17 ;
    wire sbox_inst_6_n16 ;
    wire sbox_inst_6_n15 ;
    wire sbox_inst_6_n14 ;
    wire sbox_inst_6_n13 ;
    wire sbox_inst_6_n12 ;
    wire sbox_inst_6_n11 ;
    wire sbox_inst_6_T6 ;
    wire sbox_inst_6_L0 ;
    wire sbox_inst_6_T5 ;
    wire sbox_inst_6_T4 ;
    wire sbox_inst_6_T3 ;
    wire sbox_inst_6_T2 ;
    wire sbox_inst_6_T1 ;
    wire sbox_inst_6_T0 ;
    wire sbox_inst_5_n20 ;
    wire sbox_inst_5_n19 ;
    wire sbox_inst_5_n18 ;
    wire sbox_inst_5_n17 ;
    wire sbox_inst_5_n16 ;
    wire sbox_inst_5_n15 ;
    wire sbox_inst_5_n14 ;
    wire sbox_inst_5_n13 ;
    wire sbox_inst_5_n12 ;
    wire sbox_inst_5_n11 ;
    wire sbox_inst_5_T6 ;
    wire sbox_inst_5_L0 ;
    wire sbox_inst_5_T5 ;
    wire sbox_inst_5_T4 ;
    wire sbox_inst_5_T3 ;
    wire sbox_inst_5_T2 ;
    wire sbox_inst_5_T1 ;
    wire sbox_inst_5_T0 ;
    wire sbox_inst_4_n20 ;
    wire sbox_inst_4_n19 ;
    wire sbox_inst_4_n18 ;
    wire sbox_inst_4_n17 ;
    wire sbox_inst_4_n16 ;
    wire sbox_inst_4_n15 ;
    wire sbox_inst_4_n14 ;
    wire sbox_inst_4_n13 ;
    wire sbox_inst_4_n12 ;
    wire sbox_inst_4_n11 ;
    wire sbox_inst_4_T6 ;
    wire sbox_inst_4_L0 ;
    wire sbox_inst_4_T5 ;
    wire sbox_inst_4_T4 ;
    wire sbox_inst_4_T3 ;
    wire sbox_inst_4_T2 ;
    wire sbox_inst_4_T1 ;
    wire sbox_inst_4_T0 ;
    wire sbox_inst_3_n20 ;
    wire sbox_inst_3_n19 ;
    wire sbox_inst_3_n18 ;
    wire sbox_inst_3_n17 ;
    wire sbox_inst_3_n16 ;
    wire sbox_inst_3_n15 ;
    wire sbox_inst_3_n14 ;
    wire sbox_inst_3_n13 ;
    wire sbox_inst_3_n12 ;
    wire sbox_inst_3_n11 ;
    wire sbox_inst_3_T6 ;
    wire sbox_inst_3_L0 ;
    wire sbox_inst_3_T5 ;
    wire sbox_inst_3_T4 ;
    wire sbox_inst_3_T3 ;
    wire sbox_inst_3_T2 ;
    wire sbox_inst_3_T1 ;
    wire sbox_inst_3_T0 ;
    wire sbox_inst_2_n20 ;
    wire sbox_inst_2_n19 ;
    wire sbox_inst_2_n18 ;
    wire sbox_inst_2_n17 ;
    wire sbox_inst_2_n16 ;
    wire sbox_inst_2_n15 ;
    wire sbox_inst_2_n14 ;
    wire sbox_inst_2_n13 ;
    wire sbox_inst_2_n12 ;
    wire sbox_inst_2_n11 ;
    wire sbox_inst_2_T6 ;
    wire sbox_inst_2_L0 ;
    wire sbox_inst_2_T5 ;
    wire sbox_inst_2_T4 ;
    wire sbox_inst_2_T3 ;
    wire sbox_inst_2_T2 ;
    wire sbox_inst_2_T1 ;
    wire sbox_inst_2_T0 ;
    wire sbox_inst_1_n20 ;
    wire sbox_inst_1_n19 ;
    wire sbox_inst_1_n18 ;
    wire sbox_inst_1_n17 ;
    wire sbox_inst_1_n16 ;
    wire sbox_inst_1_n15 ;
    wire sbox_inst_1_n14 ;
    wire sbox_inst_1_n13 ;
    wire sbox_inst_1_n12 ;
    wire sbox_inst_1_n11 ;
    wire sbox_inst_1_T6 ;
    wire sbox_inst_1_L0 ;
    wire sbox_inst_1_T5 ;
    wire sbox_inst_1_T4 ;
    wire sbox_inst_1_T3 ;
    wire sbox_inst_1_T2 ;
    wire sbox_inst_1_T1 ;
    wire sbox_inst_1_T0 ;
    wire sbox_inst_0_n20 ;
    wire sbox_inst_0_n19 ;
    wire sbox_inst_0_n18 ;
    wire sbox_inst_0_n17 ;
    wire sbox_inst_0_n16 ;
    wire sbox_inst_0_n15 ;
    wire sbox_inst_0_n14 ;
    wire sbox_inst_0_n13 ;
    wire sbox_inst_0_n12 ;
    wire sbox_inst_0_n11 ;
    wire sbox_inst_0_T6 ;
    wire sbox_inst_0_L0 ;
    wire sbox_inst_0_T5 ;
    wire sbox_inst_0_T4 ;
    wire sbox_inst_0_T3 ;
    wire sbox_inst_0_T2 ;
    wire sbox_inst_0_T1 ;
    wire sbox_inst_0_T0 ;
    wire [159:153] input_array ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) U29 ( .a ({input0_s3[1], input0_s2[1], input0_s1[1], input0_s0[1]}), .b ({1'b0, 1'b0, 1'b0, lfsr[1]}), .c ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, input_array_1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U30 ( .a ({input0_s3[157], input0_s2[157], input0_s1[157], input0_s0[157]}), .b ({1'b0, 1'b0, 1'b0, rev_lfsr[4]}), .c ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, input_array[157]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U31 ( .a ({input0_s3[153], input0_s2[153], input0_s1[153], input0_s0[153]}), .b ({1'b0, 1'b0, 1'b0, rev_lfsr[0]}), .c ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, input_array[153]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U32 ( .a ({input0_s3[5], input0_s2[5], input0_s1[5], input0_s0[5]}), .b ({1'b0, 1'b0, 1'b0, lfsr[5]}), .c ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, input_array_5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U33 ( .a ({input0_s3[6], input0_s2[6], input0_s1[6], input0_s0[6]}), .b ({1'b0, 1'b0, 1'b0, lfsr[6]}), .c ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, input_array_6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U34 ( .a ({input0_s3[4], input0_s2[4], input0_s1[4], input0_s0[4]}), .b ({1'b0, 1'b0, 1'b0, lfsr[4]}), .c ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, new_AGEMA_signal_1108, input_array_4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U35 ( .a ({input0_s3[3], input0_s2[3], input0_s1[3], input0_s0[3]}), .b ({1'b0, 1'b0, 1'b0, lfsr[3]}), .c ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, new_AGEMA_signal_1114, input_array_3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U36 ( .a ({input0_s3[2], input0_s2[2], input0_s1[2], input0_s0[2]}), .b ({1'b0, 1'b0, 1'b0, lfsr[2]}), .c ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, new_AGEMA_signal_1120, input_array_2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U37 ( .a ({input0_s3[0], input0_s2[0], input0_s1[0], input0_s0[0]}), .b ({1'b0, 1'b0, 1'b0, lfsr[0]}), .c ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, input_array_0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U38 ( .a ({input0_s3[159], input0_s2[159], input0_s1[159], input0_s0[159]}), .b ({1'b0, 1'b0, 1'b0, rev_lfsr[6]}), .c ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, new_AGEMA_signal_1132, input_array[159]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U39 ( .a ({input0_s3[158], input0_s2[158], input0_s1[158], input0_s0[158]}), .b ({1'b0, 1'b0, 1'b0, rev_lfsr[5]}), .c ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, input_array[158]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U40 ( .a ({input0_s3[156], input0_s2[156], input0_s1[156], input0_s0[156]}), .b ({1'b0, 1'b0, 1'b0, rev_lfsr[3]}), .c ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, new_AGEMA_signal_1144, input_array[156]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U41 ( .a ({input0_s3[155], input0_s2[155], input0_s1[155], input0_s0[155]}), .b ({1'b0, 1'b0, 1'b0, rev_lfsr[2]}), .c ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, input_array[155]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U42 ( .a ({input0_s3[154], input0_s2[154], input0_s1[154], input0_s0[154]}), .b ({1'b0, 1'b0, 1'b0, rev_lfsr[1]}), .c ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, input_array[154]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U1 ( .a ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, input_array[158]}), .b ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, input_array[157]}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, new_AGEMA_signal_2239, sbox_inst_39_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U1 ( .a ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, input_array[154]}), .b ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, input_array[153]}), .c ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, new_AGEMA_signal_2257, sbox_inst_38_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U1 ( .a ({input0_s3[150], input0_s2[150], input0_s1[150], input0_s0[150]}), .b ({input0_s3[149], input0_s2[149], input0_s1[149], input0_s0[149]}), .c ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, new_AGEMA_signal_1165, sbox_inst_37_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U1 ( .a ({input0_s3[146], input0_s2[146], input0_s1[146], input0_s0[146]}), .b ({input0_s3[145], input0_s2[145], input0_s1[145], input0_s0[145]}), .c ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, sbox_inst_36_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U1 ( .a ({input0_s3[142], input0_s2[142], input0_s1[142], input0_s0[142]}), .b ({input0_s3[141], input0_s2[141], input0_s1[141], input0_s0[141]}), .c ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, new_AGEMA_signal_1225, sbox_inst_35_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U1 ( .a ({input0_s3[138], input0_s2[138], input0_s1[138], input0_s0[138]}), .b ({input0_s3[137], input0_s2[137], input0_s1[137], input0_s0[137]}), .c ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, new_AGEMA_signal_1255, sbox_inst_34_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U1 ( .a ({input0_s3[134], input0_s2[134], input0_s1[134], input0_s0[134]}), .b ({input0_s3[133], input0_s2[133], input0_s1[133], input0_s0[133]}), .c ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, new_AGEMA_signal_1285, sbox_inst_33_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U1 ( .a ({input0_s3[130], input0_s2[130], input0_s1[130], input0_s0[130]}), .b ({input0_s3[129], input0_s2[129], input0_s1[129], input0_s0[129]}), .c ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, sbox_inst_32_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U1 ( .a ({input0_s3[126], input0_s2[126], input0_s1[126], input0_s0[126]}), .b ({input0_s3[125], input0_s2[125], input0_s1[125], input0_s0[125]}), .c ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, new_AGEMA_signal_1345, sbox_inst_31_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U1 ( .a ({input0_s3[122], input0_s2[122], input0_s1[122], input0_s0[122]}), .b ({input0_s3[121], input0_s2[121], input0_s1[121], input0_s0[121]}), .c ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, sbox_inst_30_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U1 ( .a ({input0_s3[118], input0_s2[118], input0_s1[118], input0_s0[118]}), .b ({input0_s3[117], input0_s2[117], input0_s1[117], input0_s0[117]}), .c ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, new_AGEMA_signal_1405, sbox_inst_29_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U1 ( .a ({input0_s3[114], input0_s2[114], input0_s1[114], input0_s0[114]}), .b ({input0_s3[113], input0_s2[113], input0_s1[113], input0_s0[113]}), .c ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, new_AGEMA_signal_1435, sbox_inst_28_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U1 ( .a ({input0_s3[110], input0_s2[110], input0_s1[110], input0_s0[110]}), .b ({input0_s3[109], input0_s2[109], input0_s1[109], input0_s0[109]}), .c ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, new_AGEMA_signal_1465, sbox_inst_27_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U1 ( .a ({input0_s3[106], input0_s2[106], input0_s1[106], input0_s0[106]}), .b ({input0_s3[105], input0_s2[105], input0_s1[105], input0_s0[105]}), .c ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, new_AGEMA_signal_1495, sbox_inst_26_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U1 ( .a ({input0_s3[102], input0_s2[102], input0_s1[102], input0_s0[102]}), .b ({input0_s3[101], input0_s2[101], input0_s1[101], input0_s0[101]}), .c ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, sbox_inst_25_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U1 ( .a ({input0_s3[98], input0_s2[98], input0_s1[98], input0_s0[98]}), .b ({input0_s3[97], input0_s2[97], input0_s1[97], input0_s0[97]}), .c ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, new_AGEMA_signal_1555, sbox_inst_24_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U1 ( .a ({input0_s3[94], input0_s2[94], input0_s1[94], input0_s0[94]}), .b ({input0_s3[93], input0_s2[93], input0_s1[93], input0_s0[93]}), .c ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, new_AGEMA_signal_1585, sbox_inst_23_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U1 ( .a ({input0_s3[90], input0_s2[90], input0_s1[90], input0_s0[90]}), .b ({input0_s3[89], input0_s2[89], input0_s1[89], input0_s0[89]}), .c ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, sbox_inst_22_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U1 ( .a ({input0_s3[86], input0_s2[86], input0_s1[86], input0_s0[86]}), .b ({input0_s3[85], input0_s2[85], input0_s1[85], input0_s0[85]}), .c ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, new_AGEMA_signal_1645, sbox_inst_21_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U1 ( .a ({input0_s3[82], input0_s2[82], input0_s1[82], input0_s0[82]}), .b ({input0_s3[81], input0_s2[81], input0_s1[81], input0_s0[81]}), .c ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, new_AGEMA_signal_1675, sbox_inst_20_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U1 ( .a ({input0_s3[78], input0_s2[78], input0_s1[78], input0_s0[78]}), .b ({input0_s3[77], input0_s2[77], input0_s1[77], input0_s0[77]}), .c ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, new_AGEMA_signal_1705, sbox_inst_19_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U1 ( .a ({input0_s3[74], input0_s2[74], input0_s1[74], input0_s0[74]}), .b ({input0_s3[73], input0_s2[73], input0_s1[73], input0_s0[73]}), .c ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, new_AGEMA_signal_1735, sbox_inst_18_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U1 ( .a ({input0_s3[70], input0_s2[70], input0_s1[70], input0_s0[70]}), .b ({input0_s3[69], input0_s2[69], input0_s1[69], input0_s0[69]}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, new_AGEMA_signal_1765, sbox_inst_17_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U1 ( .a ({input0_s3[66], input0_s2[66], input0_s1[66], input0_s0[66]}), .b ({input0_s3[65], input0_s2[65], input0_s1[65], input0_s0[65]}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, sbox_inst_16_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U1 ( .a ({input0_s3[62], input0_s2[62], input0_s1[62], input0_s0[62]}), .b ({input0_s3[61], input0_s2[61], input0_s1[61], input0_s0[61]}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, new_AGEMA_signal_1825, sbox_inst_15_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U1 ( .a ({input0_s3[58], input0_s2[58], input0_s1[58], input0_s0[58]}), .b ({input0_s3[57], input0_s2[57], input0_s1[57], input0_s0[57]}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, new_AGEMA_signal_1855, sbox_inst_14_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U1 ( .a ({input0_s3[54], input0_s2[54], input0_s1[54], input0_s0[54]}), .b ({input0_s3[53], input0_s2[53], input0_s1[53], input0_s0[53]}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, new_AGEMA_signal_1885, sbox_inst_13_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U1 ( .a ({input0_s3[50], input0_s2[50], input0_s1[50], input0_s0[50]}), .b ({input0_s3[49], input0_s2[49], input0_s1[49], input0_s0[49]}), .c ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, new_AGEMA_signal_1915, sbox_inst_12_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U1 ( .a ({input0_s3[46], input0_s2[46], input0_s1[46], input0_s0[46]}), .b ({input0_s3[45], input0_s2[45], input0_s1[45], input0_s0[45]}), .c ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, new_AGEMA_signal_1945, sbox_inst_11_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U1 ( .a ({input0_s3[42], input0_s2[42], input0_s1[42], input0_s0[42]}), .b ({input0_s3[41], input0_s2[41], input0_s1[41], input0_s0[41]}), .c ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, sbox_inst_10_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U1 ( .a ({input0_s3[38], input0_s2[38], input0_s1[38], input0_s0[38]}), .b ({input0_s3[37], input0_s2[37], input0_s1[37], input0_s0[37]}), .c ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, new_AGEMA_signal_2005, sbox_inst_9_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U1 ( .a ({input0_s3[34], input0_s2[34], input0_s1[34], input0_s0[34]}), .b ({input0_s3[33], input0_s2[33], input0_s1[33], input0_s0[33]}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, new_AGEMA_signal_2035, sbox_inst_8_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U1 ( .a ({input0_s3[30], input0_s2[30], input0_s1[30], input0_s0[30]}), .b ({input0_s3[29], input0_s2[29], input0_s1[29], input0_s0[29]}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, new_AGEMA_signal_2065, sbox_inst_7_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U1 ( .a ({input0_s3[26], input0_s2[26], input0_s1[26], input0_s0[26]}), .b ({input0_s3[25], input0_s2[25], input0_s1[25], input0_s0[25]}), .c ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, sbox_inst_6_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U1 ( .a ({input0_s3[22], input0_s2[22], input0_s1[22], input0_s0[22]}), .b ({input0_s3[21], input0_s2[21], input0_s1[21], input0_s0[21]}), .c ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, new_AGEMA_signal_2125, sbox_inst_5_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U1 ( .a ({input0_s3[18], input0_s2[18], input0_s1[18], input0_s0[18]}), .b ({input0_s3[17], input0_s2[17], input0_s1[17], input0_s0[17]}), .c ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, new_AGEMA_signal_2155, sbox_inst_4_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U1 ( .a ({input0_s3[14], input0_s2[14], input0_s1[14], input0_s0[14]}), .b ({input0_s3[13], input0_s2[13], input0_s1[13], input0_s0[13]}), .c ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, new_AGEMA_signal_2185, sbox_inst_3_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U1 ( .a ({input0_s3[10], input0_s2[10], input0_s1[10], input0_s0[10]}), .b ({input0_s3[9], input0_s2[9], input0_s1[9], input0_s0[9]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, new_AGEMA_signal_2215, sbox_inst_2_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U1 ( .a ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, input_array_6}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, input_array_5}), .c ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, new_AGEMA_signal_2818, sbox_inst_1_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U1 ( .a ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, new_AGEMA_signal_1120, input_array_2}), .b ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, input_array_1}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, new_AGEMA_signal_2839, sbox_inst_0_L0}) ) ;
    //ClockGatingController #(4) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U12 ( .a ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, new_AGEMA_signal_2251, sbox_inst_39_T3}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, new_AGEMA_signal_2863, sbox_inst_39_n17}), .c ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, new_AGEMA_signal_3460, sbox_inst_39_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U6 ( .a ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, sbox_inst_39_T4}), .b ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, new_AGEMA_signal_2248, sbox_inst_39_T2}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, new_AGEMA_signal_2857, sbox_inst_39_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U5 ( .a ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, new_AGEMA_signal_2245, sbox_inst_39_T1}), .b ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, input_array[158]}), .c ({new_AGEMA_signal_2862, new_AGEMA_signal_2861, new_AGEMA_signal_2860, sbox_inst_39_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U4 ( .a ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, new_AGEMA_signal_3469, sbox_inst_39_n11}), .b ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, input_array[157]}), .c ({output0_s3[39], output0_s2[39], output0_s1[39], output0_s0[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U3 ( .a ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, new_AGEMA_signal_1132, input_array[159]}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, new_AGEMA_signal_2863, sbox_inst_39_n17}), .c ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, new_AGEMA_signal_3469, sbox_inst_39_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U2 ( .a ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, new_AGEMA_signal_1144, input_array[156]}), .b ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, sbox_inst_39_T0}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, new_AGEMA_signal_2863, sbox_inst_39_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_t0_AND_U1 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, input_array[157]}), .b ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, input_array[158]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, new_AGEMA_signal_2242, sbox_inst_39_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_t1_AND_U1 ( .a ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, new_AGEMA_signal_1144, input_array[156]}), .b ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, new_AGEMA_signal_1132, input_array[159]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, new_AGEMA_signal_2245, sbox_inst_39_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_t2_AND_U1 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, input_array[157]}), .b ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, new_AGEMA_signal_1132, input_array[159]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, new_AGEMA_signal_2248, sbox_inst_39_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_t3_AND_U1 ( .a ({new_AGEMA_signal_1140, new_AGEMA_signal_1139, new_AGEMA_signal_1138, input_array[158]}), .b ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, new_AGEMA_signal_1132, input_array[159]}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, new_AGEMA_signal_2251, sbox_inst_39_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_t4_AND_U1 ( .a ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, new_AGEMA_signal_1144, input_array[156]}), .b ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, input_array[157]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, new_AGEMA_signal_2254, sbox_inst_39_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U12 ( .a ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, new_AGEMA_signal_2272, sbox_inst_38_T3}), .b ({new_AGEMA_signal_2880, new_AGEMA_signal_2879, new_AGEMA_signal_2878, sbox_inst_38_n17}), .c ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, new_AGEMA_signal_3475, sbox_inst_38_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U6 ( .a ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, new_AGEMA_signal_2275, sbox_inst_38_T4}), .b ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, new_AGEMA_signal_2269, sbox_inst_38_T2}), .c ({new_AGEMA_signal_2874, new_AGEMA_signal_2873, new_AGEMA_signal_2872, sbox_inst_38_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U5 ( .a ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, sbox_inst_38_T1}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, input_array[154]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, new_AGEMA_signal_2875, sbox_inst_38_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U4 ( .a ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, new_AGEMA_signal_3484, sbox_inst_38_n11}), .b ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, input_array[153]}), .c ({output0_s3[38], output0_s2[38], output0_s1[38], output0_s0[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U3 ( .a ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, input_array[155]}), .b ({new_AGEMA_signal_2880, new_AGEMA_signal_2879, new_AGEMA_signal_2878, sbox_inst_38_n17}), .c ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, new_AGEMA_signal_3484, sbox_inst_38_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U2 ( .a ({input0_s3[152], input0_s2[152], input0_s1[152], input0_s0[152]}), .b ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, new_AGEMA_signal_2260, sbox_inst_38_T0}), .c ({new_AGEMA_signal_2880, new_AGEMA_signal_2879, new_AGEMA_signal_2878, sbox_inst_38_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_t0_AND_U1 ( .a ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, input_array[153]}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, input_array[154]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, new_AGEMA_signal_2260, sbox_inst_38_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_t1_AND_U1 ( .a ({input0_s3[152], input0_s2[152], input0_s1[152], input0_s0[152]}), .b ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, input_array[155]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, sbox_inst_38_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_t2_AND_U1 ( .a ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, input_array[153]}), .b ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, input_array[155]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, new_AGEMA_signal_2269, sbox_inst_38_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_t3_AND_U1 ( .a ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, new_AGEMA_signal_1156, input_array[154]}), .b ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, input_array[155]}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, new_AGEMA_signal_2272, sbox_inst_38_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_t4_AND_U1 ( .a ({input0_s3[152], input0_s2[152], input0_s1[152], input0_s0[152]}), .b ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, input_array[153]}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, new_AGEMA_signal_2275, sbox_inst_38_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U12 ( .a ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, sbox_inst_37_T3}), .b ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, new_AGEMA_signal_2284, sbox_inst_37_n17}), .c ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, new_AGEMA_signal_2890, sbox_inst_37_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U6 ( .a ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, new_AGEMA_signal_1186, sbox_inst_37_T4}), .b ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, new_AGEMA_signal_1180, sbox_inst_37_T2}), .c ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, new_AGEMA_signal_2278, sbox_inst_37_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U5 ( .a ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, new_AGEMA_signal_1177, sbox_inst_37_T1}), .b ({input0_s3[150], input0_s2[150], input0_s1[150], input0_s0[150]}), .c ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, sbox_inst_37_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U4 ( .a ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, new_AGEMA_signal_2899, sbox_inst_37_n11}), .b ({input0_s3[149], input0_s2[149], input0_s1[149], input0_s0[149]}), .c ({output0_s3[37], output0_s2[37], output0_s1[37], output0_s0[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U3 ( .a ({input0_s3[151], input0_s2[151], input0_s1[151], input0_s0[151]}), .b ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, new_AGEMA_signal_2284, sbox_inst_37_n17}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, new_AGEMA_signal_2899, sbox_inst_37_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U2 ( .a ({input0_s3[148], input0_s2[148], input0_s1[148], input0_s0[148]}), .b ({new_AGEMA_signal_1170, new_AGEMA_signal_1169, new_AGEMA_signal_1168, sbox_inst_37_T0}), .c ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, new_AGEMA_signal_2284, sbox_inst_37_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_t0_AND_U1 ( .a ({input0_s3[149], input0_s2[149], input0_s1[149], input0_s0[149]}), .b ({input0_s3[150], input0_s2[150], input0_s1[150], input0_s0[150]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1170, new_AGEMA_signal_1169, new_AGEMA_signal_1168, sbox_inst_37_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_t1_AND_U1 ( .a ({input0_s3[148], input0_s2[148], input0_s1[148], input0_s0[148]}), .b ({input0_s3[151], input0_s2[151], input0_s1[151], input0_s0[151]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, new_AGEMA_signal_1177, sbox_inst_37_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_t2_AND_U1 ( .a ({input0_s3[149], input0_s2[149], input0_s1[149], input0_s0[149]}), .b ({input0_s3[151], input0_s2[151], input0_s1[151], input0_s0[151]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, new_AGEMA_signal_1180, sbox_inst_37_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_t3_AND_U1 ( .a ({input0_s3[150], input0_s2[150], input0_s1[150], input0_s0[150]}), .b ({input0_s3[151], input0_s2[151], input0_s1[151], input0_s0[151]}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, sbox_inst_37_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_t4_AND_U1 ( .a ({input0_s3[148], input0_s2[148], input0_s1[148], input0_s0[148]}), .b ({input0_s3[149], input0_s2[149], input0_s1[149], input0_s0[149]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, new_AGEMA_signal_1186, sbox_inst_37_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U12 ( .a ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, new_AGEMA_signal_1213, sbox_inst_36_T3}), .b ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, new_AGEMA_signal_2299, sbox_inst_36_n17}), .c ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, new_AGEMA_signal_2905, sbox_inst_36_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U6 ( .a ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, new_AGEMA_signal_1216, sbox_inst_36_T4}), .b ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, new_AGEMA_signal_1210, sbox_inst_36_T2}), .c ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, new_AGEMA_signal_2293, sbox_inst_36_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U5 ( .a ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, sbox_inst_36_T1}), .b ({input0_s3[146], input0_s2[146], input0_s1[146], input0_s0[146]}), .c ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, new_AGEMA_signal_2296, sbox_inst_36_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U4 ( .a ({new_AGEMA_signal_2916, new_AGEMA_signal_2915, new_AGEMA_signal_2914, sbox_inst_36_n11}), .b ({input0_s3[145], input0_s2[145], input0_s1[145], input0_s0[145]}), .c ({output0_s3[36], output0_s2[36], output0_s1[36], output0_s0[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U3 ( .a ({input0_s3[147], input0_s2[147], input0_s1[147], input0_s0[147]}), .b ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, new_AGEMA_signal_2299, sbox_inst_36_n17}), .c ({new_AGEMA_signal_2916, new_AGEMA_signal_2915, new_AGEMA_signal_2914, sbox_inst_36_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U2 ( .a ({input0_s3[144], input0_s2[144], input0_s1[144], input0_s0[144]}), .b ({new_AGEMA_signal_1200, new_AGEMA_signal_1199, new_AGEMA_signal_1198, sbox_inst_36_T0}), .c ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, new_AGEMA_signal_2299, sbox_inst_36_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_t0_AND_U1 ( .a ({input0_s3[145], input0_s2[145], input0_s1[145], input0_s0[145]}), .b ({input0_s3[146], input0_s2[146], input0_s1[146], input0_s0[146]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1200, new_AGEMA_signal_1199, new_AGEMA_signal_1198, sbox_inst_36_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_t1_AND_U1 ( .a ({input0_s3[144], input0_s2[144], input0_s1[144], input0_s0[144]}), .b ({input0_s3[147], input0_s2[147], input0_s1[147], input0_s0[147]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, sbox_inst_36_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_t2_AND_U1 ( .a ({input0_s3[145], input0_s2[145], input0_s1[145], input0_s0[145]}), .b ({input0_s3[147], input0_s2[147], input0_s1[147], input0_s0[147]}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, new_AGEMA_signal_1210, sbox_inst_36_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_t3_AND_U1 ( .a ({input0_s3[146], input0_s2[146], input0_s1[146], input0_s0[146]}), .b ({input0_s3[147], input0_s2[147], input0_s1[147], input0_s0[147]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, new_AGEMA_signal_1213, sbox_inst_36_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_t4_AND_U1 ( .a ({input0_s3[144], input0_s2[144], input0_s1[144], input0_s0[144]}), .b ({input0_s3[145], input0_s2[145], input0_s1[145], input0_s0[145]}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, new_AGEMA_signal_1216, sbox_inst_36_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U12 ( .a ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, sbox_inst_35_T3}), .b ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, sbox_inst_35_n17}), .c ({new_AGEMA_signal_2922, new_AGEMA_signal_2921, new_AGEMA_signal_2920, sbox_inst_35_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U6 ( .a ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, new_AGEMA_signal_1246, sbox_inst_35_T4}), .b ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, new_AGEMA_signal_1240, sbox_inst_35_T2}), .c ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, new_AGEMA_signal_2308, sbox_inst_35_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U5 ( .a ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, new_AGEMA_signal_1237, sbox_inst_35_T1}), .b ({input0_s3[142], input0_s2[142], input0_s1[142], input0_s0[142]}), .c ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, sbox_inst_35_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U4 ( .a ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, new_AGEMA_signal_2929, sbox_inst_35_n11}), .b ({input0_s3[141], input0_s2[141], input0_s1[141], input0_s0[141]}), .c ({output0_s3[35], output0_s2[35], output0_s1[35], output0_s0[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U3 ( .a ({input0_s3[143], input0_s2[143], input0_s1[143], input0_s0[143]}), .b ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, sbox_inst_35_n17}), .c ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, new_AGEMA_signal_2929, sbox_inst_35_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U2 ( .a ({input0_s3[140], input0_s2[140], input0_s1[140], input0_s0[140]}), .b ({new_AGEMA_signal_1230, new_AGEMA_signal_1229, new_AGEMA_signal_1228, sbox_inst_35_T0}), .c ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, new_AGEMA_signal_2314, sbox_inst_35_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_t0_AND_U1 ( .a ({input0_s3[141], input0_s2[141], input0_s1[141], input0_s0[141]}), .b ({input0_s3[142], input0_s2[142], input0_s1[142], input0_s0[142]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1230, new_AGEMA_signal_1229, new_AGEMA_signal_1228, sbox_inst_35_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_t1_AND_U1 ( .a ({input0_s3[140], input0_s2[140], input0_s1[140], input0_s0[140]}), .b ({input0_s3[143], input0_s2[143], input0_s1[143], input0_s0[143]}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, new_AGEMA_signal_1237, sbox_inst_35_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_t2_AND_U1 ( .a ({input0_s3[141], input0_s2[141], input0_s1[141], input0_s0[141]}), .b ({input0_s3[143], input0_s2[143], input0_s1[143], input0_s0[143]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, new_AGEMA_signal_1240, sbox_inst_35_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_t3_AND_U1 ( .a ({input0_s3[142], input0_s2[142], input0_s1[142], input0_s0[142]}), .b ({input0_s3[143], input0_s2[143], input0_s1[143], input0_s0[143]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, sbox_inst_35_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_t4_AND_U1 ( .a ({input0_s3[140], input0_s2[140], input0_s1[140], input0_s0[140]}), .b ({input0_s3[141], input0_s2[141], input0_s1[141], input0_s0[141]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, new_AGEMA_signal_1246, sbox_inst_35_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U12 ( .a ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, new_AGEMA_signal_1273, sbox_inst_34_T3}), .b ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, sbox_inst_34_n17}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, new_AGEMA_signal_2935, sbox_inst_34_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U6 ( .a ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, new_AGEMA_signal_1276, sbox_inst_34_T4}), .b ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, sbox_inst_34_T2}), .c ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, new_AGEMA_signal_2323, sbox_inst_34_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U5 ( .a ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, sbox_inst_34_T1}), .b ({input0_s3[138], input0_s2[138], input0_s1[138], input0_s0[138]}), .c ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, sbox_inst_34_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U4 ( .a ({new_AGEMA_signal_2946, new_AGEMA_signal_2945, new_AGEMA_signal_2944, sbox_inst_34_n11}), .b ({input0_s3[137], input0_s2[137], input0_s1[137], input0_s0[137]}), .c ({output0_s3[34], output0_s2[34], output0_s1[34], output0_s0[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U3 ( .a ({input0_s3[139], input0_s2[139], input0_s1[139], input0_s0[139]}), .b ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, sbox_inst_34_n17}), .c ({new_AGEMA_signal_2946, new_AGEMA_signal_2945, new_AGEMA_signal_2944, sbox_inst_34_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U2 ( .a ({input0_s3[136], input0_s2[136], input0_s1[136], input0_s0[136]}), .b ({new_AGEMA_signal_1260, new_AGEMA_signal_1259, new_AGEMA_signal_1258, sbox_inst_34_T0}), .c ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, new_AGEMA_signal_2329, sbox_inst_34_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_t0_AND_U1 ( .a ({input0_s3[137], input0_s2[137], input0_s1[137], input0_s0[137]}), .b ({input0_s3[138], input0_s2[138], input0_s1[138], input0_s0[138]}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1260, new_AGEMA_signal_1259, new_AGEMA_signal_1258, sbox_inst_34_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_t1_AND_U1 ( .a ({input0_s3[136], input0_s2[136], input0_s1[136], input0_s0[136]}), .b ({input0_s3[139], input0_s2[139], input0_s1[139], input0_s0[139]}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, sbox_inst_34_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_t2_AND_U1 ( .a ({input0_s3[137], input0_s2[137], input0_s1[137], input0_s0[137]}), .b ({input0_s3[139], input0_s2[139], input0_s1[139], input0_s0[139]}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, sbox_inst_34_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_t3_AND_U1 ( .a ({input0_s3[138], input0_s2[138], input0_s1[138], input0_s0[138]}), .b ({input0_s3[139], input0_s2[139], input0_s1[139], input0_s0[139]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, new_AGEMA_signal_1273, sbox_inst_34_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_t4_AND_U1 ( .a ({input0_s3[136], input0_s2[136], input0_s1[136], input0_s0[136]}), .b ({input0_s3[137], input0_s2[137], input0_s1[137], input0_s0[137]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, new_AGEMA_signal_1276, sbox_inst_34_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U12 ( .a ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, new_AGEMA_signal_1303, sbox_inst_33_T3}), .b ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, sbox_inst_33_n17}), .c ({new_AGEMA_signal_2952, new_AGEMA_signal_2951, new_AGEMA_signal_2950, sbox_inst_33_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U6 ( .a ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, sbox_inst_33_T4}), .b ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, new_AGEMA_signal_1300, sbox_inst_33_T2}), .c ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, sbox_inst_33_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U5 ( .a ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, new_AGEMA_signal_1297, sbox_inst_33_T1}), .b ({input0_s3[134], input0_s2[134], input0_s1[134], input0_s0[134]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, sbox_inst_33_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U4 ( .a ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, new_AGEMA_signal_2959, sbox_inst_33_n11}), .b ({input0_s3[133], input0_s2[133], input0_s1[133], input0_s0[133]}), .c ({output0_s3[33], output0_s2[33], output0_s1[33], output0_s0[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U3 ( .a ({input0_s3[135], input0_s2[135], input0_s1[135], input0_s0[135]}), .b ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, sbox_inst_33_n17}), .c ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, new_AGEMA_signal_2959, sbox_inst_33_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U2 ( .a ({input0_s3[132], input0_s2[132], input0_s1[132], input0_s0[132]}), .b ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, new_AGEMA_signal_1288, sbox_inst_33_T0}), .c ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, sbox_inst_33_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_t0_AND_U1 ( .a ({input0_s3[133], input0_s2[133], input0_s1[133], input0_s0[133]}), .b ({input0_s3[134], input0_s2[134], input0_s1[134], input0_s0[134]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, new_AGEMA_signal_1288, sbox_inst_33_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_t1_AND_U1 ( .a ({input0_s3[132], input0_s2[132], input0_s1[132], input0_s0[132]}), .b ({input0_s3[135], input0_s2[135], input0_s1[135], input0_s0[135]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, new_AGEMA_signal_1297, sbox_inst_33_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_t2_AND_U1 ( .a ({input0_s3[133], input0_s2[133], input0_s1[133], input0_s0[133]}), .b ({input0_s3[135], input0_s2[135], input0_s1[135], input0_s0[135]}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, new_AGEMA_signal_1300, sbox_inst_33_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_t3_AND_U1 ( .a ({input0_s3[134], input0_s2[134], input0_s1[134], input0_s0[134]}), .b ({input0_s3[135], input0_s2[135], input0_s1[135], input0_s0[135]}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, new_AGEMA_signal_1303, sbox_inst_33_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_t4_AND_U1 ( .a ({input0_s3[132], input0_s2[132], input0_s1[132], input0_s0[132]}), .b ({input0_s3[133], input0_s2[133], input0_s1[133], input0_s0[133]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, new_AGEMA_signal_1306, sbox_inst_33_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U12 ( .a ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, new_AGEMA_signal_1333, sbox_inst_32_T3}), .b ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, sbox_inst_32_n17}), .c ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, new_AGEMA_signal_2965, sbox_inst_32_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U6 ( .a ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, new_AGEMA_signal_1336, sbox_inst_32_T4}), .b ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, sbox_inst_32_T2}), .c ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, sbox_inst_32_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U5 ( .a ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, sbox_inst_32_T1}), .b ({input0_s3[130], input0_s2[130], input0_s1[130], input0_s0[130]}), .c ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, new_AGEMA_signal_2356, sbox_inst_32_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U4 ( .a ({new_AGEMA_signal_2976, new_AGEMA_signal_2975, new_AGEMA_signal_2974, sbox_inst_32_n11}), .b ({input0_s3[129], input0_s2[129], input0_s1[129], input0_s0[129]}), .c ({output0_s3[32], output0_s2[32], output0_s1[32], output0_s0[32]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U3 ( .a ({input0_s3[131], input0_s2[131], input0_s1[131], input0_s0[131]}), .b ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, sbox_inst_32_n17}), .c ({new_AGEMA_signal_2976, new_AGEMA_signal_2975, new_AGEMA_signal_2974, sbox_inst_32_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U2 ( .a ({input0_s3[128], input0_s2[128], input0_s1[128], input0_s0[128]}), .b ({new_AGEMA_signal_1320, new_AGEMA_signal_1319, new_AGEMA_signal_1318, sbox_inst_32_T0}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, sbox_inst_32_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_t0_AND_U1 ( .a ({input0_s3[129], input0_s2[129], input0_s1[129], input0_s0[129]}), .b ({input0_s3[130], input0_s2[130], input0_s1[130], input0_s0[130]}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1320, new_AGEMA_signal_1319, new_AGEMA_signal_1318, sbox_inst_32_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_t1_AND_U1 ( .a ({input0_s3[128], input0_s2[128], input0_s1[128], input0_s0[128]}), .b ({input0_s3[131], input0_s2[131], input0_s1[131], input0_s0[131]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, sbox_inst_32_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_t2_AND_U1 ( .a ({input0_s3[129], input0_s2[129], input0_s1[129], input0_s0[129]}), .b ({input0_s3[131], input0_s2[131], input0_s1[131], input0_s0[131]}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, sbox_inst_32_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_t3_AND_U1 ( .a ({input0_s3[130], input0_s2[130], input0_s1[130], input0_s0[130]}), .b ({input0_s3[131], input0_s2[131], input0_s1[131], input0_s0[131]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, new_AGEMA_signal_1333, sbox_inst_32_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_t4_AND_U1 ( .a ({input0_s3[128], input0_s2[128], input0_s1[128], input0_s0[128]}), .b ({input0_s3[129], input0_s2[129], input0_s1[129], input0_s0[129]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, new_AGEMA_signal_1336, sbox_inst_32_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U12 ( .a ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, new_AGEMA_signal_1363, sbox_inst_31_T3}), .b ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, sbox_inst_31_n17}), .c ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, new_AGEMA_signal_2980, sbox_inst_31_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U6 ( .a ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, sbox_inst_31_T4}), .b ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, new_AGEMA_signal_1360, sbox_inst_31_T2}), .c ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, new_AGEMA_signal_2368, sbox_inst_31_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U5 ( .a ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, new_AGEMA_signal_1357, sbox_inst_31_T1}), .b ({input0_s3[126], input0_s2[126], input0_s1[126], input0_s0[126]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, sbox_inst_31_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U4 ( .a ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, new_AGEMA_signal_2989, sbox_inst_31_n11}), .b ({input0_s3[125], input0_s2[125], input0_s1[125], input0_s0[125]}), .c ({output0_s3[31], output0_s2[31], output0_s1[31], output0_s0[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U3 ( .a ({input0_s3[127], input0_s2[127], input0_s1[127], input0_s0[127]}), .b ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, sbox_inst_31_n17}), .c ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, new_AGEMA_signal_2989, sbox_inst_31_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U2 ( .a ({input0_s3[124], input0_s2[124], input0_s1[124], input0_s0[124]}), .b ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, new_AGEMA_signal_1348, sbox_inst_31_T0}), .c ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, new_AGEMA_signal_2374, sbox_inst_31_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_t0_AND_U1 ( .a ({input0_s3[125], input0_s2[125], input0_s1[125], input0_s0[125]}), .b ({input0_s3[126], input0_s2[126], input0_s1[126], input0_s0[126]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, new_AGEMA_signal_1348, sbox_inst_31_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_t1_AND_U1 ( .a ({input0_s3[124], input0_s2[124], input0_s1[124], input0_s0[124]}), .b ({input0_s3[127], input0_s2[127], input0_s1[127], input0_s0[127]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, new_AGEMA_signal_1357, sbox_inst_31_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_t2_AND_U1 ( .a ({input0_s3[125], input0_s2[125], input0_s1[125], input0_s0[125]}), .b ({input0_s3[127], input0_s2[127], input0_s1[127], input0_s0[127]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, new_AGEMA_signal_1360, sbox_inst_31_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_t3_AND_U1 ( .a ({input0_s3[126], input0_s2[126], input0_s1[126], input0_s0[126]}), .b ({input0_s3[127], input0_s2[127], input0_s1[127], input0_s0[127]}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, new_AGEMA_signal_1363, sbox_inst_31_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_t4_AND_U1 ( .a ({input0_s3[124], input0_s2[124], input0_s1[124], input0_s0[124]}), .b ({input0_s3[125], input0_s2[125], input0_s1[125], input0_s0[125]}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, new_AGEMA_signal_1366, sbox_inst_31_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U12 ( .a ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, new_AGEMA_signal_1393, sbox_inst_30_T3}), .b ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, sbox_inst_30_n17}), .c ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, new_AGEMA_signal_2995, sbox_inst_30_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U6 ( .a ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, new_AGEMA_signal_1396, sbox_inst_30_T4}), .b ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, new_AGEMA_signal_1390, sbox_inst_30_T2}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, new_AGEMA_signal_2383, sbox_inst_30_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U5 ( .a ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, sbox_inst_30_T1}), .b ({input0_s3[122], input0_s2[122], input0_s1[122], input0_s0[122]}), .c ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, sbox_inst_30_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U4 ( .a ({new_AGEMA_signal_3006, new_AGEMA_signal_3005, new_AGEMA_signal_3004, sbox_inst_30_n11}), .b ({input0_s3[121], input0_s2[121], input0_s1[121], input0_s0[121]}), .c ({output0_s3[30], output0_s2[30], output0_s1[30], output0_s0[30]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U3 ( .a ({input0_s3[123], input0_s2[123], input0_s1[123], input0_s0[123]}), .b ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, sbox_inst_30_n17}), .c ({new_AGEMA_signal_3006, new_AGEMA_signal_3005, new_AGEMA_signal_3004, sbox_inst_30_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U2 ( .a ({input0_s3[120], input0_s2[120], input0_s1[120], input0_s0[120]}), .b ({new_AGEMA_signal_1380, new_AGEMA_signal_1379, new_AGEMA_signal_1378, sbox_inst_30_T0}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, sbox_inst_30_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_t0_AND_U1 ( .a ({input0_s3[121], input0_s2[121], input0_s1[121], input0_s0[121]}), .b ({input0_s3[122], input0_s2[122], input0_s1[122], input0_s0[122]}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1380, new_AGEMA_signal_1379, new_AGEMA_signal_1378, sbox_inst_30_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_t1_AND_U1 ( .a ({input0_s3[120], input0_s2[120], input0_s1[120], input0_s0[120]}), .b ({input0_s3[123], input0_s2[123], input0_s1[123], input0_s0[123]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, sbox_inst_30_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_t2_AND_U1 ( .a ({input0_s3[121], input0_s2[121], input0_s1[121], input0_s0[121]}), .b ({input0_s3[123], input0_s2[123], input0_s1[123], input0_s0[123]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, new_AGEMA_signal_1390, sbox_inst_30_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_t3_AND_U1 ( .a ({input0_s3[122], input0_s2[122], input0_s1[122], input0_s0[122]}), .b ({input0_s3[123], input0_s2[123], input0_s1[123], input0_s0[123]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, new_AGEMA_signal_1393, sbox_inst_30_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_t4_AND_U1 ( .a ({input0_s3[120], input0_s2[120], input0_s1[120], input0_s0[120]}), .b ({input0_s3[121], input0_s2[121], input0_s1[121], input0_s0[121]}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, new_AGEMA_signal_1396, sbox_inst_30_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U12 ( .a ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, sbox_inst_29_T3}), .b ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, sbox_inst_29_n17}), .c ({new_AGEMA_signal_3012, new_AGEMA_signal_3011, new_AGEMA_signal_3010, sbox_inst_29_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U6 ( .a ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, sbox_inst_29_T4}), .b ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, new_AGEMA_signal_1420, sbox_inst_29_T2}), .c ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, sbox_inst_29_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U5 ( .a ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, new_AGEMA_signal_1417, sbox_inst_29_T1}), .b ({input0_s3[118], input0_s2[118], input0_s1[118], input0_s0[118]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, sbox_inst_29_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U4 ( .a ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, new_AGEMA_signal_3019, sbox_inst_29_n11}), .b ({input0_s3[117], input0_s2[117], input0_s1[117], input0_s0[117]}), .c ({output0_s3[29], output0_s2[29], output0_s1[29], output0_s0[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U3 ( .a ({input0_s3[119], input0_s2[119], input0_s1[119], input0_s0[119]}), .b ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, sbox_inst_29_n17}), .c ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, new_AGEMA_signal_3019, sbox_inst_29_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U2 ( .a ({input0_s3[116], input0_s2[116], input0_s1[116], input0_s0[116]}), .b ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, new_AGEMA_signal_1408, sbox_inst_29_T0}), .c ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, sbox_inst_29_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_t0_AND_U1 ( .a ({input0_s3[117], input0_s2[117], input0_s1[117], input0_s0[117]}), .b ({input0_s3[118], input0_s2[118], input0_s1[118], input0_s0[118]}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, new_AGEMA_signal_1408, sbox_inst_29_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_t1_AND_U1 ( .a ({input0_s3[116], input0_s2[116], input0_s1[116], input0_s0[116]}), .b ({input0_s3[119], input0_s2[119], input0_s1[119], input0_s0[119]}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, new_AGEMA_signal_1417, sbox_inst_29_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_t2_AND_U1 ( .a ({input0_s3[117], input0_s2[117], input0_s1[117], input0_s0[117]}), .b ({input0_s3[119], input0_s2[119], input0_s1[119], input0_s0[119]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, new_AGEMA_signal_1420, sbox_inst_29_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_t3_AND_U1 ( .a ({input0_s3[118], input0_s2[118], input0_s1[118], input0_s0[118]}), .b ({input0_s3[119], input0_s2[119], input0_s1[119], input0_s0[119]}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, sbox_inst_29_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_t4_AND_U1 ( .a ({input0_s3[116], input0_s2[116], input0_s1[116], input0_s0[116]}), .b ({input0_s3[117], input0_s2[117], input0_s1[117], input0_s0[117]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, new_AGEMA_signal_1426, sbox_inst_29_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U12 ( .a ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, new_AGEMA_signal_1453, sbox_inst_28_T3}), .b ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, new_AGEMA_signal_2419, sbox_inst_28_n17}), .c ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, new_AGEMA_signal_3025, sbox_inst_28_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U6 ( .a ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, new_AGEMA_signal_1456, sbox_inst_28_T4}), .b ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, new_AGEMA_signal_1450, sbox_inst_28_T2}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2413, sbox_inst_28_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U5 ( .a ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, sbox_inst_28_T1}), .b ({input0_s3[114], input0_s2[114], input0_s1[114], input0_s0[114]}), .c ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, sbox_inst_28_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U4 ( .a ({new_AGEMA_signal_3036, new_AGEMA_signal_3035, new_AGEMA_signal_3034, sbox_inst_28_n11}), .b ({input0_s3[113], input0_s2[113], input0_s1[113], input0_s0[113]}), .c ({output0_s3[28], output0_s2[28], output0_s1[28], output0_s0[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U3 ( .a ({input0_s3[115], input0_s2[115], input0_s1[115], input0_s0[115]}), .b ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, new_AGEMA_signal_2419, sbox_inst_28_n17}), .c ({new_AGEMA_signal_3036, new_AGEMA_signal_3035, new_AGEMA_signal_3034, sbox_inst_28_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U2 ( .a ({input0_s3[112], input0_s2[112], input0_s1[112], input0_s0[112]}), .b ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, new_AGEMA_signal_1438, sbox_inst_28_T0}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, new_AGEMA_signal_2419, sbox_inst_28_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_t0_AND_U1 ( .a ({input0_s3[113], input0_s2[113], input0_s1[113], input0_s0[113]}), .b ({input0_s3[114], input0_s2[114], input0_s1[114], input0_s0[114]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1440, new_AGEMA_signal_1439, new_AGEMA_signal_1438, sbox_inst_28_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_t1_AND_U1 ( .a ({input0_s3[112], input0_s2[112], input0_s1[112], input0_s0[112]}), .b ({input0_s3[115], input0_s2[115], input0_s1[115], input0_s0[115]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, sbox_inst_28_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_t2_AND_U1 ( .a ({input0_s3[113], input0_s2[113], input0_s1[113], input0_s0[113]}), .b ({input0_s3[115], input0_s2[115], input0_s1[115], input0_s0[115]}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, new_AGEMA_signal_1450, sbox_inst_28_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_t3_AND_U1 ( .a ({input0_s3[114], input0_s2[114], input0_s1[114], input0_s0[114]}), .b ({input0_s3[115], input0_s2[115], input0_s1[115], input0_s0[115]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, new_AGEMA_signal_1453, sbox_inst_28_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_t4_AND_U1 ( .a ({input0_s3[112], input0_s2[112], input0_s1[112], input0_s0[112]}), .b ({input0_s3[113], input0_s2[113], input0_s1[113], input0_s0[113]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, new_AGEMA_signal_1456, sbox_inst_28_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U12 ( .a ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, sbox_inst_27_T3}), .b ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, sbox_inst_27_n17}), .c ({new_AGEMA_signal_3042, new_AGEMA_signal_3041, new_AGEMA_signal_3040, sbox_inst_27_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U6 ( .a ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, new_AGEMA_signal_1486, sbox_inst_27_T4}), .b ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, sbox_inst_27_T2}), .c ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, new_AGEMA_signal_2428, sbox_inst_27_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U5 ( .a ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, new_AGEMA_signal_1477, sbox_inst_27_T1}), .b ({input0_s3[110], input0_s2[110], input0_s1[110], input0_s0[110]}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, sbox_inst_27_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U4 ( .a ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, new_AGEMA_signal_3049, sbox_inst_27_n11}), .b ({input0_s3[109], input0_s2[109], input0_s1[109], input0_s0[109]}), .c ({output0_s3[27], output0_s2[27], output0_s1[27], output0_s0[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U3 ( .a ({input0_s3[111], input0_s2[111], input0_s1[111], input0_s0[111]}), .b ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, sbox_inst_27_n17}), .c ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, new_AGEMA_signal_3049, sbox_inst_27_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U2 ( .a ({input0_s3[108], input0_s2[108], input0_s1[108], input0_s0[108]}), .b ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, new_AGEMA_signal_1468, sbox_inst_27_T0}), .c ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, sbox_inst_27_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_t0_AND_U1 ( .a ({input0_s3[109], input0_s2[109], input0_s1[109], input0_s0[109]}), .b ({input0_s3[110], input0_s2[110], input0_s1[110], input0_s0[110]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, new_AGEMA_signal_1468, sbox_inst_27_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_t1_AND_U1 ( .a ({input0_s3[108], input0_s2[108], input0_s1[108], input0_s0[108]}), .b ({input0_s3[111], input0_s2[111], input0_s1[111], input0_s0[111]}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, new_AGEMA_signal_1477, sbox_inst_27_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_t2_AND_U1 ( .a ({input0_s3[109], input0_s2[109], input0_s1[109], input0_s0[109]}), .b ({input0_s3[111], input0_s2[111], input0_s1[111], input0_s0[111]}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, sbox_inst_27_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_t3_AND_U1 ( .a ({input0_s3[110], input0_s2[110], input0_s1[110], input0_s0[110]}), .b ({input0_s3[111], input0_s2[111], input0_s1[111], input0_s0[111]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, sbox_inst_27_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_t4_AND_U1 ( .a ({input0_s3[108], input0_s2[108], input0_s1[108], input0_s0[108]}), .b ({input0_s3[109], input0_s2[109], input0_s1[109], input0_s0[109]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, new_AGEMA_signal_1486, sbox_inst_27_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U12 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, new_AGEMA_signal_1513, sbox_inst_26_T3}), .b ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, sbox_inst_26_n17}), .c ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, new_AGEMA_signal_3055, sbox_inst_26_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U6 ( .a ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, sbox_inst_26_T4}), .b ({new_AGEMA_signal_1512, new_AGEMA_signal_1511, new_AGEMA_signal_1510, sbox_inst_26_T2}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, new_AGEMA_signal_2443, sbox_inst_26_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U5 ( .a ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, sbox_inst_26_T1}), .b ({input0_s3[106], input0_s2[106], input0_s1[106], input0_s0[106]}), .c ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, sbox_inst_26_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U4 ( .a ({new_AGEMA_signal_3066, new_AGEMA_signal_3065, new_AGEMA_signal_3064, sbox_inst_26_n11}), .b ({input0_s3[105], input0_s2[105], input0_s1[105], input0_s0[105]}), .c ({output0_s3[26], output0_s2[26], output0_s1[26], output0_s0[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U3 ( .a ({input0_s3[107], input0_s2[107], input0_s1[107], input0_s0[107]}), .b ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, sbox_inst_26_n17}), .c ({new_AGEMA_signal_3066, new_AGEMA_signal_3065, new_AGEMA_signal_3064, sbox_inst_26_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U2 ( .a ({input0_s3[104], input0_s2[104], input0_s1[104], input0_s0[104]}), .b ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, sbox_inst_26_T0}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, sbox_inst_26_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_t0_AND_U1 ( .a ({input0_s3[105], input0_s2[105], input0_s1[105], input0_s0[105]}), .b ({input0_s3[106], input0_s2[106], input0_s1[106], input0_s0[106]}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1500, new_AGEMA_signal_1499, new_AGEMA_signal_1498, sbox_inst_26_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_t1_AND_U1 ( .a ({input0_s3[104], input0_s2[104], input0_s1[104], input0_s0[104]}), .b ({input0_s3[107], input0_s2[107], input0_s1[107], input0_s0[107]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, sbox_inst_26_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_t2_AND_U1 ( .a ({input0_s3[105], input0_s2[105], input0_s1[105], input0_s0[105]}), .b ({input0_s3[107], input0_s2[107], input0_s1[107], input0_s0[107]}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1512, new_AGEMA_signal_1511, new_AGEMA_signal_1510, sbox_inst_26_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_t3_AND_U1 ( .a ({input0_s3[106], input0_s2[106], input0_s1[106], input0_s0[106]}), .b ({input0_s3[107], input0_s2[107], input0_s1[107], input0_s0[107]}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, new_AGEMA_signal_1513, sbox_inst_26_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_t4_AND_U1 ( .a ({input0_s3[104], input0_s2[104], input0_s1[104], input0_s0[104]}), .b ({input0_s3[105], input0_s2[105], input0_s1[105], input0_s0[105]}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, new_AGEMA_signal_1516, sbox_inst_26_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U12 ( .a ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, sbox_inst_25_T3}), .b ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, new_AGEMA_signal_2464, sbox_inst_25_n17}), .c ({new_AGEMA_signal_3072, new_AGEMA_signal_3071, new_AGEMA_signal_3070, sbox_inst_25_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U6 ( .a ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, new_AGEMA_signal_1546, sbox_inst_25_T4}), .b ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, new_AGEMA_signal_1540, sbox_inst_25_T2}), .c ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, sbox_inst_25_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U5 ( .a ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, new_AGEMA_signal_1537, sbox_inst_25_T1}), .b ({input0_s3[102], input0_s2[102], input0_s1[102], input0_s0[102]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, new_AGEMA_signal_2461, sbox_inst_25_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U4 ( .a ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, new_AGEMA_signal_3079, sbox_inst_25_n11}), .b ({input0_s3[101], input0_s2[101], input0_s1[101], input0_s0[101]}), .c ({output0_s3[25], output0_s2[25], output0_s1[25], output0_s0[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U3 ( .a ({input0_s3[103], input0_s2[103], input0_s1[103], input0_s0[103]}), .b ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, new_AGEMA_signal_2464, sbox_inst_25_n17}), .c ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, new_AGEMA_signal_3079, sbox_inst_25_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U2 ( .a ({input0_s3[100], input0_s2[100], input0_s1[100], input0_s0[100]}), .b ({new_AGEMA_signal_1530, new_AGEMA_signal_1529, new_AGEMA_signal_1528, sbox_inst_25_T0}), .c ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, new_AGEMA_signal_2464, sbox_inst_25_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_t0_AND_U1 ( .a ({input0_s3[101], input0_s2[101], input0_s1[101], input0_s0[101]}), .b ({input0_s3[102], input0_s2[102], input0_s1[102], input0_s0[102]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1530, new_AGEMA_signal_1529, new_AGEMA_signal_1528, sbox_inst_25_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_t1_AND_U1 ( .a ({input0_s3[100], input0_s2[100], input0_s1[100], input0_s0[100]}), .b ({input0_s3[103], input0_s2[103], input0_s1[103], input0_s0[103]}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, new_AGEMA_signal_1537, sbox_inst_25_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_t2_AND_U1 ( .a ({input0_s3[101], input0_s2[101], input0_s1[101], input0_s0[101]}), .b ({input0_s3[103], input0_s2[103], input0_s1[103], input0_s0[103]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, new_AGEMA_signal_1540, sbox_inst_25_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_t3_AND_U1 ( .a ({input0_s3[102], input0_s2[102], input0_s1[102], input0_s0[102]}), .b ({input0_s3[103], input0_s2[103], input0_s1[103], input0_s0[103]}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, sbox_inst_25_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_t4_AND_U1 ( .a ({input0_s3[100], input0_s2[100], input0_s1[100], input0_s0[100]}), .b ({input0_s3[101], input0_s2[101], input0_s1[101], input0_s0[101]}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, new_AGEMA_signal_1546, sbox_inst_25_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U12 ( .a ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, new_AGEMA_signal_1573, sbox_inst_24_T3}), .b ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, new_AGEMA_signal_2479, sbox_inst_24_n17}), .c ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, new_AGEMA_signal_3085, sbox_inst_24_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U6 ( .a ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, new_AGEMA_signal_1576, sbox_inst_24_T4}), .b ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, sbox_inst_24_T2}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, new_AGEMA_signal_2473, sbox_inst_24_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U5 ( .a ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, new_AGEMA_signal_1567, sbox_inst_24_T1}), .b ({input0_s3[98], input0_s2[98], input0_s1[98], input0_s0[98]}), .c ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, new_AGEMA_signal_2476, sbox_inst_24_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U4 ( .a ({new_AGEMA_signal_3096, new_AGEMA_signal_3095, new_AGEMA_signal_3094, sbox_inst_24_n11}), .b ({input0_s3[97], input0_s2[97], input0_s1[97], input0_s0[97]}), .c ({output0_s3[24], output0_s2[24], output0_s1[24], output0_s0[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U3 ( .a ({input0_s3[99], input0_s2[99], input0_s1[99], input0_s0[99]}), .b ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, new_AGEMA_signal_2479, sbox_inst_24_n17}), .c ({new_AGEMA_signal_3096, new_AGEMA_signal_3095, new_AGEMA_signal_3094, sbox_inst_24_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U2 ( .a ({input0_s3[96], input0_s2[96], input0_s1[96], input0_s0[96]}), .b ({new_AGEMA_signal_1560, new_AGEMA_signal_1559, new_AGEMA_signal_1558, sbox_inst_24_T0}), .c ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, new_AGEMA_signal_2479, sbox_inst_24_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_t0_AND_U1 ( .a ({input0_s3[97], input0_s2[97], input0_s1[97], input0_s0[97]}), .b ({input0_s3[98], input0_s2[98], input0_s1[98], input0_s0[98]}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1560, new_AGEMA_signal_1559, new_AGEMA_signal_1558, sbox_inst_24_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_t1_AND_U1 ( .a ({input0_s3[96], input0_s2[96], input0_s1[96], input0_s0[96]}), .b ({input0_s3[99], input0_s2[99], input0_s1[99], input0_s0[99]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, new_AGEMA_signal_1567, sbox_inst_24_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_t2_AND_U1 ( .a ({input0_s3[97], input0_s2[97], input0_s1[97], input0_s0[97]}), .b ({input0_s3[99], input0_s2[99], input0_s1[99], input0_s0[99]}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, sbox_inst_24_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_t3_AND_U1 ( .a ({input0_s3[98], input0_s2[98], input0_s1[98], input0_s0[98]}), .b ({input0_s3[99], input0_s2[99], input0_s1[99], input0_s0[99]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, new_AGEMA_signal_1573, sbox_inst_24_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_t4_AND_U1 ( .a ({input0_s3[96], input0_s2[96], input0_s1[96], input0_s0[96]}), .b ({input0_s3[97], input0_s2[97], input0_s1[97], input0_s0[97]}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, new_AGEMA_signal_1576, sbox_inst_24_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U12 ( .a ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, new_AGEMA_signal_1603, sbox_inst_23_T3}), .b ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, sbox_inst_23_n17}), .c ({new_AGEMA_signal_3102, new_AGEMA_signal_3101, new_AGEMA_signal_3100, sbox_inst_23_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U6 ( .a ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, sbox_inst_23_T4}), .b ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, new_AGEMA_signal_1600, sbox_inst_23_T2}), .c ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, new_AGEMA_signal_2488, sbox_inst_23_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U5 ( .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, sbox_inst_23_T1}), .b ({input0_s3[94], input0_s2[94], input0_s1[94], input0_s0[94]}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, new_AGEMA_signal_2491, sbox_inst_23_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U4 ( .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, new_AGEMA_signal_3109, sbox_inst_23_n11}), .b ({input0_s3[93], input0_s2[93], input0_s1[93], input0_s0[93]}), .c ({output0_s3[23], output0_s2[23], output0_s1[23], output0_s0[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U3 ( .a ({input0_s3[95], input0_s2[95], input0_s1[95], input0_s0[95]}), .b ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, sbox_inst_23_n17}), .c ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, new_AGEMA_signal_3109, sbox_inst_23_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U2 ( .a ({input0_s3[92], input0_s2[92], input0_s1[92], input0_s0[92]}), .b ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, new_AGEMA_signal_1588, sbox_inst_23_T0}), .c ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, sbox_inst_23_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_t0_AND_U1 ( .a ({input0_s3[93], input0_s2[93], input0_s1[93], input0_s0[93]}), .b ({input0_s3[94], input0_s2[94], input0_s1[94], input0_s0[94]}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, new_AGEMA_signal_1588, sbox_inst_23_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_t1_AND_U1 ( .a ({input0_s3[92], input0_s2[92], input0_s1[92], input0_s0[92]}), .b ({input0_s3[95], input0_s2[95], input0_s1[95], input0_s0[95]}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, sbox_inst_23_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_t2_AND_U1 ( .a ({input0_s3[93], input0_s2[93], input0_s1[93], input0_s0[93]}), .b ({input0_s3[95], input0_s2[95], input0_s1[95], input0_s0[95]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, new_AGEMA_signal_1600, sbox_inst_23_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_t3_AND_U1 ( .a ({input0_s3[94], input0_s2[94], input0_s1[94], input0_s0[94]}), .b ({input0_s3[95], input0_s2[95], input0_s1[95], input0_s0[95]}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, new_AGEMA_signal_1603, sbox_inst_23_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_t4_AND_U1 ( .a ({input0_s3[92], input0_s2[92], input0_s1[92], input0_s0[92]}), .b ({input0_s3[93], input0_s2[93], input0_s1[93], input0_s0[93]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, new_AGEMA_signal_1606, sbox_inst_23_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U12 ( .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, sbox_inst_22_T3}), .b ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, new_AGEMA_signal_2509, sbox_inst_22_n17}), .c ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, new_AGEMA_signal_3115, sbox_inst_22_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U6 ( .a ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, new_AGEMA_signal_1636, sbox_inst_22_T4}), .b ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, new_AGEMA_signal_1630, sbox_inst_22_T2}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, new_AGEMA_signal_2503, sbox_inst_22_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U5 ( .a ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, new_AGEMA_signal_1627, sbox_inst_22_T1}), .b ({input0_s3[90], input0_s2[90], input0_s1[90], input0_s0[90]}), .c ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, new_AGEMA_signal_2506, sbox_inst_22_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U4 ( .a ({new_AGEMA_signal_3126, new_AGEMA_signal_3125, new_AGEMA_signal_3124, sbox_inst_22_n11}), .b ({input0_s3[89], input0_s2[89], input0_s1[89], input0_s0[89]}), .c ({output0_s3[22], output0_s2[22], output0_s1[22], output0_s0[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U3 ( .a ({input0_s3[91], input0_s2[91], input0_s1[91], input0_s0[91]}), .b ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, new_AGEMA_signal_2509, sbox_inst_22_n17}), .c ({new_AGEMA_signal_3126, new_AGEMA_signal_3125, new_AGEMA_signal_3124, sbox_inst_22_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U2 ( .a ({input0_s3[88], input0_s2[88], input0_s1[88], input0_s0[88]}), .b ({new_AGEMA_signal_1620, new_AGEMA_signal_1619, new_AGEMA_signal_1618, sbox_inst_22_T0}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, new_AGEMA_signal_2509, sbox_inst_22_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_t0_AND_U1 ( .a ({input0_s3[89], input0_s2[89], input0_s1[89], input0_s0[89]}), .b ({input0_s3[90], input0_s2[90], input0_s1[90], input0_s0[90]}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1620, new_AGEMA_signal_1619, new_AGEMA_signal_1618, sbox_inst_22_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_t1_AND_U1 ( .a ({input0_s3[88], input0_s2[88], input0_s1[88], input0_s0[88]}), .b ({input0_s3[91], input0_s2[91], input0_s1[91], input0_s0[91]}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, new_AGEMA_signal_1627, sbox_inst_22_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_t2_AND_U1 ( .a ({input0_s3[89], input0_s2[89], input0_s1[89], input0_s0[89]}), .b ({input0_s3[91], input0_s2[91], input0_s1[91], input0_s0[91]}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, new_AGEMA_signal_1630, sbox_inst_22_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_t3_AND_U1 ( .a ({input0_s3[90], input0_s2[90], input0_s1[90], input0_s0[90]}), .b ({input0_s3[91], input0_s2[91], input0_s1[91], input0_s0[91]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, sbox_inst_22_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_t4_AND_U1 ( .a ({input0_s3[88], input0_s2[88], input0_s1[88], input0_s0[88]}), .b ({input0_s3[89], input0_s2[89], input0_s1[89], input0_s0[89]}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, new_AGEMA_signal_1636, sbox_inst_22_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U12 ( .a ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, new_AGEMA_signal_1663, sbox_inst_21_T3}), .b ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, new_AGEMA_signal_2524, sbox_inst_21_n17}), .c ({new_AGEMA_signal_3132, new_AGEMA_signal_3131, new_AGEMA_signal_3130, sbox_inst_21_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U6 ( .a ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, new_AGEMA_signal_1666, sbox_inst_21_T4}), .b ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, sbox_inst_21_T2}), .c ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, new_AGEMA_signal_2518, sbox_inst_21_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U5 ( .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, new_AGEMA_signal_1657, sbox_inst_21_T1}), .b ({input0_s3[86], input0_s2[86], input0_s1[86], input0_s0[86]}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, new_AGEMA_signal_2521, sbox_inst_21_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U4 ( .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, new_AGEMA_signal_3139, sbox_inst_21_n11}), .b ({input0_s3[85], input0_s2[85], input0_s1[85], input0_s0[85]}), .c ({output0_s3[21], output0_s2[21], output0_s1[21], output0_s0[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U3 ( .a ({input0_s3[87], input0_s2[87], input0_s1[87], input0_s0[87]}), .b ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, new_AGEMA_signal_2524, sbox_inst_21_n17}), .c ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, new_AGEMA_signal_3139, sbox_inst_21_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U2 ( .a ({input0_s3[84], input0_s2[84], input0_s1[84], input0_s0[84]}), .b ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, new_AGEMA_signal_1648, sbox_inst_21_T0}), .c ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, new_AGEMA_signal_2524, sbox_inst_21_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_t0_AND_U1 ( .a ({input0_s3[85], input0_s2[85], input0_s1[85], input0_s0[85]}), .b ({input0_s3[86], input0_s2[86], input0_s1[86], input0_s0[86]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, new_AGEMA_signal_1648, sbox_inst_21_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_t1_AND_U1 ( .a ({input0_s3[84], input0_s2[84], input0_s1[84], input0_s0[84]}), .b ({input0_s3[87], input0_s2[87], input0_s1[87], input0_s0[87]}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, new_AGEMA_signal_1657, sbox_inst_21_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_t2_AND_U1 ( .a ({input0_s3[85], input0_s2[85], input0_s1[85], input0_s0[85]}), .b ({input0_s3[87], input0_s2[87], input0_s1[87], input0_s0[87]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, sbox_inst_21_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_t3_AND_U1 ( .a ({input0_s3[86], input0_s2[86], input0_s1[86], input0_s0[86]}), .b ({input0_s3[87], input0_s2[87], input0_s1[87], input0_s0[87]}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, new_AGEMA_signal_1663, sbox_inst_21_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_t4_AND_U1 ( .a ({input0_s3[84], input0_s2[84], input0_s1[84], input0_s0[84]}), .b ({input0_s3[85], input0_s2[85], input0_s1[85], input0_s0[85]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, new_AGEMA_signal_1666, sbox_inst_21_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U12 ( .a ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, new_AGEMA_signal_1693, sbox_inst_20_T3}), .b ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, new_AGEMA_signal_2539, sbox_inst_20_n17}), .c ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, new_AGEMA_signal_3145, sbox_inst_20_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U6 ( .a ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, new_AGEMA_signal_1696, sbox_inst_20_T4}), .b ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, new_AGEMA_signal_1690, sbox_inst_20_T2}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, new_AGEMA_signal_2533, sbox_inst_20_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U5 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, sbox_inst_20_T1}), .b ({input0_s3[82], input0_s2[82], input0_s1[82], input0_s0[82]}), .c ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, new_AGEMA_signal_2536, sbox_inst_20_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U4 ( .a ({new_AGEMA_signal_3156, new_AGEMA_signal_3155, new_AGEMA_signal_3154, sbox_inst_20_n11}), .b ({input0_s3[81], input0_s2[81], input0_s1[81], input0_s0[81]}), .c ({output0_s3[20], output0_s2[20], output0_s1[20], output0_s0[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U3 ( .a ({input0_s3[83], input0_s2[83], input0_s1[83], input0_s0[83]}), .b ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, new_AGEMA_signal_2539, sbox_inst_20_n17}), .c ({new_AGEMA_signal_3156, new_AGEMA_signal_3155, new_AGEMA_signal_3154, sbox_inst_20_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U2 ( .a ({input0_s3[80], input0_s2[80], input0_s1[80], input0_s0[80]}), .b ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, sbox_inst_20_T0}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, new_AGEMA_signal_2539, sbox_inst_20_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_t0_AND_U1 ( .a ({input0_s3[81], input0_s2[81], input0_s1[81], input0_s0[81]}), .b ({input0_s3[82], input0_s2[82], input0_s1[82], input0_s0[82]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_1680, new_AGEMA_signal_1679, new_AGEMA_signal_1678, sbox_inst_20_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_t1_AND_U1 ( .a ({input0_s3[80], input0_s2[80], input0_s1[80], input0_s0[80]}), .b ({input0_s3[83], input0_s2[83], input0_s1[83], input0_s0[83]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, sbox_inst_20_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_t2_AND_U1 ( .a ({input0_s3[81], input0_s2[81], input0_s1[81], input0_s0[81]}), .b ({input0_s3[83], input0_s2[83], input0_s1[83], input0_s0[83]}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, new_AGEMA_signal_1690, sbox_inst_20_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_t3_AND_U1 ( .a ({input0_s3[82], input0_s2[82], input0_s1[82], input0_s0[82]}), .b ({input0_s3[83], input0_s2[83], input0_s1[83], input0_s0[83]}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, new_AGEMA_signal_1693, sbox_inst_20_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_t4_AND_U1 ( .a ({input0_s3[80], input0_s2[80], input0_s1[80], input0_s0[80]}), .b ({input0_s3[81], input0_s2[81], input0_s1[81], input0_s0[81]}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, new_AGEMA_signal_1696, sbox_inst_20_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U12 ( .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, sbox_inst_19_T3}), .b ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, new_AGEMA_signal_2554, sbox_inst_19_n17}), .c ({new_AGEMA_signal_3162, new_AGEMA_signal_3161, new_AGEMA_signal_3160, sbox_inst_19_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U6 ( .a ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, new_AGEMA_signal_1726, sbox_inst_19_T4}), .b ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, new_AGEMA_signal_1720, sbox_inst_19_T2}), .c ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, new_AGEMA_signal_2548, sbox_inst_19_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U5 ( .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, new_AGEMA_signal_1717, sbox_inst_19_T1}), .b ({input0_s3[78], input0_s2[78], input0_s1[78], input0_s0[78]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, new_AGEMA_signal_2551, sbox_inst_19_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U4 ( .a ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, new_AGEMA_signal_3169, sbox_inst_19_n11}), .b ({input0_s3[77], input0_s2[77], input0_s1[77], input0_s0[77]}), .c ({output0_s3[19], output0_s2[19], output0_s1[19], output0_s0[19]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U3 ( .a ({input0_s3[79], input0_s2[79], input0_s1[79], input0_s0[79]}), .b ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, new_AGEMA_signal_2554, sbox_inst_19_n17}), .c ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, new_AGEMA_signal_3169, sbox_inst_19_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U2 ( .a ({input0_s3[76], input0_s2[76], input0_s1[76], input0_s0[76]}), .b ({new_AGEMA_signal_1710, new_AGEMA_signal_1709, new_AGEMA_signal_1708, sbox_inst_19_T0}), .c ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, new_AGEMA_signal_2554, sbox_inst_19_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_t0_AND_U1 ( .a ({input0_s3[77], input0_s2[77], input0_s1[77], input0_s0[77]}), .b ({input0_s3[78], input0_s2[78], input0_s1[78], input0_s0[78]}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_1710, new_AGEMA_signal_1709, new_AGEMA_signal_1708, sbox_inst_19_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_t1_AND_U1 ( .a ({input0_s3[76], input0_s2[76], input0_s1[76], input0_s0[76]}), .b ({input0_s3[79], input0_s2[79], input0_s1[79], input0_s0[79]}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, new_AGEMA_signal_1717, sbox_inst_19_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_t2_AND_U1 ( .a ({input0_s3[77], input0_s2[77], input0_s1[77], input0_s0[77]}), .b ({input0_s3[79], input0_s2[79], input0_s1[79], input0_s0[79]}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, new_AGEMA_signal_1720, sbox_inst_19_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_t3_AND_U1 ( .a ({input0_s3[78], input0_s2[78], input0_s1[78], input0_s0[78]}), .b ({input0_s3[79], input0_s2[79], input0_s1[79], input0_s0[79]}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, sbox_inst_19_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_t4_AND_U1 ( .a ({input0_s3[76], input0_s2[76], input0_s1[76], input0_s0[76]}), .b ({input0_s3[77], input0_s2[77], input0_s1[77], input0_s0[77]}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, new_AGEMA_signal_1726, sbox_inst_19_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U12 ( .a ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, new_AGEMA_signal_1753, sbox_inst_18_T3}), .b ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, new_AGEMA_signal_2569, sbox_inst_18_n17}), .c ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, new_AGEMA_signal_3175, sbox_inst_18_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U6 ( .a ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, new_AGEMA_signal_1756, sbox_inst_18_T4}), .b ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, sbox_inst_18_T2}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, new_AGEMA_signal_2563, sbox_inst_18_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U5 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, sbox_inst_18_T1}), .b ({input0_s3[74], input0_s2[74], input0_s1[74], input0_s0[74]}), .c ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, sbox_inst_18_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U4 ( .a ({new_AGEMA_signal_3186, new_AGEMA_signal_3185, new_AGEMA_signal_3184, sbox_inst_18_n11}), .b ({input0_s3[73], input0_s2[73], input0_s1[73], input0_s0[73]}), .c ({output0_s3[18], output0_s2[18], output0_s1[18], output0_s0[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U3 ( .a ({input0_s3[75], input0_s2[75], input0_s1[75], input0_s0[75]}), .b ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, new_AGEMA_signal_2569, sbox_inst_18_n17}), .c ({new_AGEMA_signal_3186, new_AGEMA_signal_3185, new_AGEMA_signal_3184, sbox_inst_18_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U2 ( .a ({input0_s3[72], input0_s2[72], input0_s1[72], input0_s0[72]}), .b ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, new_AGEMA_signal_1738, sbox_inst_18_T0}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, new_AGEMA_signal_2569, sbox_inst_18_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_t0_AND_U1 ( .a ({input0_s3[73], input0_s2[73], input0_s1[73], input0_s0[73]}), .b ({input0_s3[74], input0_s2[74], input0_s1[74], input0_s0[74]}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_1740, new_AGEMA_signal_1739, new_AGEMA_signal_1738, sbox_inst_18_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_t1_AND_U1 ( .a ({input0_s3[72], input0_s2[72], input0_s1[72], input0_s0[72]}), .b ({input0_s3[75], input0_s2[75], input0_s1[75], input0_s0[75]}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, sbox_inst_18_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_t2_AND_U1 ( .a ({input0_s3[73], input0_s2[73], input0_s1[73], input0_s0[73]}), .b ({input0_s3[75], input0_s2[75], input0_s1[75], input0_s0[75]}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, sbox_inst_18_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_t3_AND_U1 ( .a ({input0_s3[74], input0_s2[74], input0_s1[74], input0_s0[74]}), .b ({input0_s3[75], input0_s2[75], input0_s1[75], input0_s0[75]}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, new_AGEMA_signal_1753, sbox_inst_18_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_t4_AND_U1 ( .a ({input0_s3[72], input0_s2[72], input0_s1[72], input0_s0[72]}), .b ({input0_s3[73], input0_s2[73], input0_s1[73], input0_s0[73]}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, new_AGEMA_signal_1756, sbox_inst_18_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U12 ( .a ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, new_AGEMA_signal_1783, sbox_inst_17_T3}), .b ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, new_AGEMA_signal_2584, sbox_inst_17_n17}), .c ({new_AGEMA_signal_3192, new_AGEMA_signal_3191, new_AGEMA_signal_3190, sbox_inst_17_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U6 ( .a ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, sbox_inst_17_T4}), .b ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, new_AGEMA_signal_1780, sbox_inst_17_T2}), .c ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, sbox_inst_17_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U5 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, sbox_inst_17_T1}), .b ({input0_s3[70], input0_s2[70], input0_s1[70], input0_s0[70]}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, new_AGEMA_signal_2581, sbox_inst_17_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U4 ( .a ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, new_AGEMA_signal_3199, sbox_inst_17_n11}), .b ({input0_s3[69], input0_s2[69], input0_s1[69], input0_s0[69]}), .c ({output0_s3[17], output0_s2[17], output0_s1[17], output0_s0[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U3 ( .a ({input0_s3[71], input0_s2[71], input0_s1[71], input0_s0[71]}), .b ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, new_AGEMA_signal_2584, sbox_inst_17_n17}), .c ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, new_AGEMA_signal_3199, sbox_inst_17_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U2 ( .a ({input0_s3[68], input0_s2[68], input0_s1[68], input0_s0[68]}), .b ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, new_AGEMA_signal_1768, sbox_inst_17_T0}), .c ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, new_AGEMA_signal_2584, sbox_inst_17_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_t0_AND_U1 ( .a ({input0_s3[69], input0_s2[69], input0_s1[69], input0_s0[69]}), .b ({input0_s3[70], input0_s2[70], input0_s1[70], input0_s0[70]}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, new_AGEMA_signal_1768, sbox_inst_17_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_t1_AND_U1 ( .a ({input0_s3[68], input0_s2[68], input0_s1[68], input0_s0[68]}), .b ({input0_s3[71], input0_s2[71], input0_s1[71], input0_s0[71]}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, sbox_inst_17_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_t2_AND_U1 ( .a ({input0_s3[69], input0_s2[69], input0_s1[69], input0_s0[69]}), .b ({input0_s3[71], input0_s2[71], input0_s1[71], input0_s0[71]}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, new_AGEMA_signal_1780, sbox_inst_17_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_t3_AND_U1 ( .a ({input0_s3[70], input0_s2[70], input0_s1[70], input0_s0[70]}), .b ({input0_s3[71], input0_s2[71], input0_s1[71], input0_s0[71]}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, new_AGEMA_signal_1783, sbox_inst_17_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_t4_AND_U1 ( .a ({input0_s3[68], input0_s2[68], input0_s1[68], input0_s0[68]}), .b ({input0_s3[69], input0_s2[69], input0_s1[69], input0_s0[69]}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, new_AGEMA_signal_1786, sbox_inst_17_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U12 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, sbox_inst_16_T3}), .b ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, new_AGEMA_signal_2599, sbox_inst_16_n17}), .c ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, new_AGEMA_signal_3205, sbox_inst_16_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U6 ( .a ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, new_AGEMA_signal_1816, sbox_inst_16_T4}), .b ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, new_AGEMA_signal_1810, sbox_inst_16_T2}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, new_AGEMA_signal_2593, sbox_inst_16_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U5 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, new_AGEMA_signal_1807, sbox_inst_16_T1}), .b ({input0_s3[66], input0_s2[66], input0_s1[66], input0_s0[66]}), .c ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, new_AGEMA_signal_2596, sbox_inst_16_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U4 ( .a ({new_AGEMA_signal_3216, new_AGEMA_signal_3215, new_AGEMA_signal_3214, sbox_inst_16_n11}), .b ({input0_s3[65], input0_s2[65], input0_s1[65], input0_s0[65]}), .c ({output0_s3[16], output0_s2[16], output0_s1[16], output0_s0[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U3 ( .a ({input0_s3[67], input0_s2[67], input0_s1[67], input0_s0[67]}), .b ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, new_AGEMA_signal_2599, sbox_inst_16_n17}), .c ({new_AGEMA_signal_3216, new_AGEMA_signal_3215, new_AGEMA_signal_3214, sbox_inst_16_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U2 ( .a ({input0_s3[64], input0_s2[64], input0_s1[64], input0_s0[64]}), .b ({new_AGEMA_signal_1800, new_AGEMA_signal_1799, new_AGEMA_signal_1798, sbox_inst_16_T0}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, new_AGEMA_signal_2599, sbox_inst_16_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_t0_AND_U1 ( .a ({input0_s3[65], input0_s2[65], input0_s1[65], input0_s0[65]}), .b ({input0_s3[66], input0_s2[66], input0_s1[66], input0_s0[66]}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_1800, new_AGEMA_signal_1799, new_AGEMA_signal_1798, sbox_inst_16_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_t1_AND_U1 ( .a ({input0_s3[64], input0_s2[64], input0_s1[64], input0_s0[64]}), .b ({input0_s3[67], input0_s2[67], input0_s1[67], input0_s0[67]}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, new_AGEMA_signal_1807, sbox_inst_16_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_t2_AND_U1 ( .a ({input0_s3[65], input0_s2[65], input0_s1[65], input0_s0[65]}), .b ({input0_s3[67], input0_s2[67], input0_s1[67], input0_s0[67]}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, new_AGEMA_signal_1810, sbox_inst_16_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_t3_AND_U1 ( .a ({input0_s3[66], input0_s2[66], input0_s1[66], input0_s0[66]}), .b ({input0_s3[67], input0_s2[67], input0_s1[67], input0_s0[67]}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, sbox_inst_16_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_t4_AND_U1 ( .a ({input0_s3[64], input0_s2[64], input0_s1[64], input0_s0[64]}), .b ({input0_s3[65], input0_s2[65], input0_s1[65], input0_s0[65]}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, new_AGEMA_signal_1816, sbox_inst_16_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U12 ( .a ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, new_AGEMA_signal_1843, sbox_inst_15_T3}), .b ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, new_AGEMA_signal_2614, sbox_inst_15_n17}), .c ({new_AGEMA_signal_3222, new_AGEMA_signal_3221, new_AGEMA_signal_3220, sbox_inst_15_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U6 ( .a ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, new_AGEMA_signal_1846, sbox_inst_15_T4}), .b ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, sbox_inst_15_T2}), .c ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, new_AGEMA_signal_2608, sbox_inst_15_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U5 ( .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, new_AGEMA_signal_1837, sbox_inst_15_T1}), .b ({input0_s3[62], input0_s2[62], input0_s1[62], input0_s0[62]}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, new_AGEMA_signal_2611, sbox_inst_15_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U4 ( .a ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, new_AGEMA_signal_3229, sbox_inst_15_n11}), .b ({input0_s3[61], input0_s2[61], input0_s1[61], input0_s0[61]}), .c ({output0_s3[15], output0_s2[15], output0_s1[15], output0_s0[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U3 ( .a ({input0_s3[63], input0_s2[63], input0_s1[63], input0_s0[63]}), .b ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, new_AGEMA_signal_2614, sbox_inst_15_n17}), .c ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, new_AGEMA_signal_3229, sbox_inst_15_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U2 ( .a ({input0_s3[60], input0_s2[60], input0_s1[60], input0_s0[60]}), .b ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, new_AGEMA_signal_1828, sbox_inst_15_T0}), .c ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, new_AGEMA_signal_2614, sbox_inst_15_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_t0_AND_U1 ( .a ({input0_s3[61], input0_s2[61], input0_s1[61], input0_s0[61]}), .b ({input0_s3[62], input0_s2[62], input0_s1[62], input0_s0[62]}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, new_AGEMA_signal_1828, sbox_inst_15_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_t1_AND_U1 ( .a ({input0_s3[60], input0_s2[60], input0_s1[60], input0_s0[60]}), .b ({input0_s3[63], input0_s2[63], input0_s1[63], input0_s0[63]}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, new_AGEMA_signal_1837, sbox_inst_15_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_t2_AND_U1 ( .a ({input0_s3[61], input0_s2[61], input0_s1[61], input0_s0[61]}), .b ({input0_s3[63], input0_s2[63], input0_s1[63], input0_s0[63]}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, sbox_inst_15_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_t3_AND_U1 ( .a ({input0_s3[62], input0_s2[62], input0_s1[62], input0_s0[62]}), .b ({input0_s3[63], input0_s2[63], input0_s1[63], input0_s0[63]}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, new_AGEMA_signal_1843, sbox_inst_15_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_t4_AND_U1 ( .a ({input0_s3[60], input0_s2[60], input0_s1[60], input0_s0[60]}), .b ({input0_s3[61], input0_s2[61], input0_s1[61], input0_s0[61]}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, new_AGEMA_signal_1846, sbox_inst_15_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U12 ( .a ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, new_AGEMA_signal_1873, sbox_inst_14_T3}), .b ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, new_AGEMA_signal_2629, sbox_inst_14_n17}), .c ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, new_AGEMA_signal_3235, sbox_inst_14_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U6 ( .a ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, new_AGEMA_signal_1876, sbox_inst_14_T4}), .b ({new_AGEMA_signal_1872, new_AGEMA_signal_1871, new_AGEMA_signal_1870, sbox_inst_14_T2}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, new_AGEMA_signal_2623, sbox_inst_14_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U5 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, sbox_inst_14_T1}), .b ({input0_s3[58], input0_s2[58], input0_s1[58], input0_s0[58]}), .c ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, new_AGEMA_signal_2626, sbox_inst_14_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U4 ( .a ({new_AGEMA_signal_3246, new_AGEMA_signal_3245, new_AGEMA_signal_3244, sbox_inst_14_n11}), .b ({input0_s3[57], input0_s2[57], input0_s1[57], input0_s0[57]}), .c ({output0_s3[14], output0_s2[14], output0_s1[14], output0_s0[14]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U3 ( .a ({input0_s3[59], input0_s2[59], input0_s1[59], input0_s0[59]}), .b ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, new_AGEMA_signal_2629, sbox_inst_14_n17}), .c ({new_AGEMA_signal_3246, new_AGEMA_signal_3245, new_AGEMA_signal_3244, sbox_inst_14_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U2 ( .a ({input0_s3[56], input0_s2[56], input0_s1[56], input0_s0[56]}), .b ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, sbox_inst_14_T0}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, new_AGEMA_signal_2629, sbox_inst_14_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_t0_AND_U1 ( .a ({input0_s3[57], input0_s2[57], input0_s1[57], input0_s0[57]}), .b ({input0_s3[58], input0_s2[58], input0_s1[58], input0_s0[58]}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, new_AGEMA_signal_1858, sbox_inst_14_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_t1_AND_U1 ( .a ({input0_s3[56], input0_s2[56], input0_s1[56], input0_s0[56]}), .b ({input0_s3[59], input0_s2[59], input0_s1[59], input0_s0[59]}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, sbox_inst_14_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_t2_AND_U1 ( .a ({input0_s3[57], input0_s2[57], input0_s1[57], input0_s0[57]}), .b ({input0_s3[59], input0_s2[59], input0_s1[59], input0_s0[59]}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_1872, new_AGEMA_signal_1871, new_AGEMA_signal_1870, sbox_inst_14_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_t3_AND_U1 ( .a ({input0_s3[58], input0_s2[58], input0_s1[58], input0_s0[58]}), .b ({input0_s3[59], input0_s2[59], input0_s1[59], input0_s0[59]}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, new_AGEMA_signal_1873, sbox_inst_14_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_t4_AND_U1 ( .a ({input0_s3[56], input0_s2[56], input0_s1[56], input0_s0[56]}), .b ({input0_s3[57], input0_s2[57], input0_s1[57], input0_s0[57]}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, new_AGEMA_signal_1876, sbox_inst_14_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U12 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, sbox_inst_13_T3}), .b ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, new_AGEMA_signal_2644, sbox_inst_13_n17}), .c ({new_AGEMA_signal_3252, new_AGEMA_signal_3251, new_AGEMA_signal_3250, sbox_inst_13_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U6 ( .a ({new_AGEMA_signal_1908, new_AGEMA_signal_1907, new_AGEMA_signal_1906, sbox_inst_13_T4}), .b ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, new_AGEMA_signal_1900, sbox_inst_13_T2}), .c ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, sbox_inst_13_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U5 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, new_AGEMA_signal_1897, sbox_inst_13_T1}), .b ({input0_s3[54], input0_s2[54], input0_s1[54], input0_s0[54]}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, new_AGEMA_signal_2641, sbox_inst_13_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U4 ( .a ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, new_AGEMA_signal_3259, sbox_inst_13_n11}), .b ({input0_s3[53], input0_s2[53], input0_s1[53], input0_s0[53]}), .c ({output0_s3[13], output0_s2[13], output0_s1[13], output0_s0[13]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U3 ( .a ({input0_s3[55], input0_s2[55], input0_s1[55], input0_s0[55]}), .b ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, new_AGEMA_signal_2644, sbox_inst_13_n17}), .c ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, new_AGEMA_signal_3259, sbox_inst_13_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U2 ( .a ({input0_s3[52], input0_s2[52], input0_s1[52], input0_s0[52]}), .b ({new_AGEMA_signal_1890, new_AGEMA_signal_1889, new_AGEMA_signal_1888, sbox_inst_13_T0}), .c ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, new_AGEMA_signal_2644, sbox_inst_13_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_t0_AND_U1 ( .a ({input0_s3[53], input0_s2[53], input0_s1[53], input0_s0[53]}), .b ({input0_s3[54], input0_s2[54], input0_s1[54], input0_s0[54]}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_1890, new_AGEMA_signal_1889, new_AGEMA_signal_1888, sbox_inst_13_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_t1_AND_U1 ( .a ({input0_s3[52], input0_s2[52], input0_s1[52], input0_s0[52]}), .b ({input0_s3[55], input0_s2[55], input0_s1[55], input0_s0[55]}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, new_AGEMA_signal_1897, sbox_inst_13_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_t2_AND_U1 ( .a ({input0_s3[53], input0_s2[53], input0_s1[53], input0_s0[53]}), .b ({input0_s3[55], input0_s2[55], input0_s1[55], input0_s0[55]}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, new_AGEMA_signal_1900, sbox_inst_13_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_t3_AND_U1 ( .a ({input0_s3[54], input0_s2[54], input0_s1[54], input0_s0[54]}), .b ({input0_s3[55], input0_s2[55], input0_s1[55], input0_s0[55]}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, sbox_inst_13_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_t4_AND_U1 ( .a ({input0_s3[52], input0_s2[52], input0_s1[52], input0_s0[52]}), .b ({input0_s3[53], input0_s2[53], input0_s1[53], input0_s0[53]}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_1908, new_AGEMA_signal_1907, new_AGEMA_signal_1906, sbox_inst_13_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U12 ( .a ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, new_AGEMA_signal_1933, sbox_inst_12_T3}), .b ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, new_AGEMA_signal_2659, sbox_inst_12_n17}), .c ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, new_AGEMA_signal_3265, sbox_inst_12_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U6 ( .a ({new_AGEMA_signal_1938, new_AGEMA_signal_1937, new_AGEMA_signal_1936, sbox_inst_12_T4}), .b ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, sbox_inst_12_T2}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, new_AGEMA_signal_2653, sbox_inst_12_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U5 ( .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, sbox_inst_12_T1}), .b ({input0_s3[50], input0_s2[50], input0_s1[50], input0_s0[50]}), .c ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, new_AGEMA_signal_2656, sbox_inst_12_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U4 ( .a ({new_AGEMA_signal_3276, new_AGEMA_signal_3275, new_AGEMA_signal_3274, sbox_inst_12_n11}), .b ({input0_s3[49], input0_s2[49], input0_s1[49], input0_s0[49]}), .c ({output0_s3[12], output0_s2[12], output0_s1[12], output0_s0[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U3 ( .a ({input0_s3[51], input0_s2[51], input0_s1[51], input0_s0[51]}), .b ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, new_AGEMA_signal_2659, sbox_inst_12_n17}), .c ({new_AGEMA_signal_3276, new_AGEMA_signal_3275, new_AGEMA_signal_3274, sbox_inst_12_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U2 ( .a ({input0_s3[48], input0_s2[48], input0_s1[48], input0_s0[48]}), .b ({new_AGEMA_signal_1920, new_AGEMA_signal_1919, new_AGEMA_signal_1918, sbox_inst_12_T0}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, new_AGEMA_signal_2659, sbox_inst_12_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_t0_AND_U1 ( .a ({input0_s3[49], input0_s2[49], input0_s1[49], input0_s0[49]}), .b ({input0_s3[50], input0_s2[50], input0_s1[50], input0_s0[50]}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_1920, new_AGEMA_signal_1919, new_AGEMA_signal_1918, sbox_inst_12_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_t1_AND_U1 ( .a ({input0_s3[48], input0_s2[48], input0_s1[48], input0_s0[48]}), .b ({input0_s3[51], input0_s2[51], input0_s1[51], input0_s0[51]}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, sbox_inst_12_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_t2_AND_U1 ( .a ({input0_s3[49], input0_s2[49], input0_s1[49], input0_s0[49]}), .b ({input0_s3[51], input0_s2[51], input0_s1[51], input0_s0[51]}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, sbox_inst_12_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_t3_AND_U1 ( .a ({input0_s3[50], input0_s2[50], input0_s1[50], input0_s0[50]}), .b ({input0_s3[51], input0_s2[51], input0_s1[51], input0_s0[51]}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, new_AGEMA_signal_1933, sbox_inst_12_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_t4_AND_U1 ( .a ({input0_s3[48], input0_s2[48], input0_s1[48], input0_s0[48]}), .b ({input0_s3[49], input0_s2[49], input0_s1[49], input0_s0[49]}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_1938, new_AGEMA_signal_1937, new_AGEMA_signal_1936, sbox_inst_12_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U12 ( .a ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, new_AGEMA_signal_1963, sbox_inst_11_T3}), .b ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, sbox_inst_11_n17}), .c ({new_AGEMA_signal_3282, new_AGEMA_signal_3281, new_AGEMA_signal_3280, sbox_inst_11_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U6 ( .a ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, sbox_inst_11_T4}), .b ({new_AGEMA_signal_1962, new_AGEMA_signal_1961, new_AGEMA_signal_1960, sbox_inst_11_T2}), .c ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, new_AGEMA_signal_2668, sbox_inst_11_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U5 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, sbox_inst_11_T1}), .b ({input0_s3[46], input0_s2[46], input0_s1[46], input0_s0[46]}), .c ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, new_AGEMA_signal_2671, sbox_inst_11_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U4 ( .a ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, new_AGEMA_signal_3289, sbox_inst_11_n11}), .b ({input0_s3[45], input0_s2[45], input0_s1[45], input0_s0[45]}), .c ({output0_s3[11], output0_s2[11], output0_s1[11], output0_s0[11]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U3 ( .a ({input0_s3[47], input0_s2[47], input0_s1[47], input0_s0[47]}), .b ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, sbox_inst_11_n17}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, new_AGEMA_signal_3289, sbox_inst_11_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U2 ( .a ({input0_s3[44], input0_s2[44], input0_s1[44], input0_s0[44]}), .b ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, new_AGEMA_signal_1948, sbox_inst_11_T0}), .c ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, sbox_inst_11_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_t0_AND_U1 ( .a ({input0_s3[45], input0_s2[45], input0_s1[45], input0_s0[45]}), .b ({input0_s3[46], input0_s2[46], input0_s1[46], input0_s0[46]}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, new_AGEMA_signal_1948, sbox_inst_11_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_t1_AND_U1 ( .a ({input0_s3[44], input0_s2[44], input0_s1[44], input0_s0[44]}), .b ({input0_s3[47], input0_s2[47], input0_s1[47], input0_s0[47]}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, sbox_inst_11_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_t2_AND_U1 ( .a ({input0_s3[45], input0_s2[45], input0_s1[45], input0_s0[45]}), .b ({input0_s3[47], input0_s2[47], input0_s1[47], input0_s0[47]}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_1962, new_AGEMA_signal_1961, new_AGEMA_signal_1960, sbox_inst_11_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_t3_AND_U1 ( .a ({input0_s3[46], input0_s2[46], input0_s1[46], input0_s0[46]}), .b ({input0_s3[47], input0_s2[47], input0_s1[47], input0_s0[47]}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, new_AGEMA_signal_1963, sbox_inst_11_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_t4_AND_U1 ( .a ({input0_s3[44], input0_s2[44], input0_s1[44], input0_s0[44]}), .b ({input0_s3[45], input0_s2[45], input0_s1[45], input0_s0[45]}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, new_AGEMA_signal_1966, sbox_inst_11_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U12 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, sbox_inst_10_T3}), .b ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, new_AGEMA_signal_2689, sbox_inst_10_n17}), .c ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, new_AGEMA_signal_3295, sbox_inst_10_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U6 ( .a ({new_AGEMA_signal_1998, new_AGEMA_signal_1997, new_AGEMA_signal_1996, sbox_inst_10_T4}), .b ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, new_AGEMA_signal_1990, sbox_inst_10_T2}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, new_AGEMA_signal_2683, sbox_inst_10_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U5 ( .a ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, new_AGEMA_signal_1987, sbox_inst_10_T1}), .b ({input0_s3[42], input0_s2[42], input0_s1[42], input0_s0[42]}), .c ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, sbox_inst_10_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U4 ( .a ({new_AGEMA_signal_3306, new_AGEMA_signal_3305, new_AGEMA_signal_3304, sbox_inst_10_n11}), .b ({input0_s3[41], input0_s2[41], input0_s1[41], input0_s0[41]}), .c ({output0_s3[10], output0_s2[10], output0_s1[10], output0_s0[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U3 ( .a ({input0_s3[43], input0_s2[43], input0_s1[43], input0_s0[43]}), .b ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, new_AGEMA_signal_2689, sbox_inst_10_n17}), .c ({new_AGEMA_signal_3306, new_AGEMA_signal_3305, new_AGEMA_signal_3304, sbox_inst_10_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U2 ( .a ({input0_s3[40], input0_s2[40], input0_s1[40], input0_s0[40]}), .b ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, new_AGEMA_signal_1978, sbox_inst_10_T0}), .c ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, new_AGEMA_signal_2689, sbox_inst_10_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_t0_AND_U1 ( .a ({input0_s3[41], input0_s2[41], input0_s1[41], input0_s0[41]}), .b ({input0_s3[42], input0_s2[42], input0_s1[42], input0_s0[42]}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, new_AGEMA_signal_1978, sbox_inst_10_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_t1_AND_U1 ( .a ({input0_s3[40], input0_s2[40], input0_s1[40], input0_s0[40]}), .b ({input0_s3[43], input0_s2[43], input0_s1[43], input0_s0[43]}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, new_AGEMA_signal_1987, sbox_inst_10_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_t2_AND_U1 ( .a ({input0_s3[41], input0_s2[41], input0_s1[41], input0_s0[41]}), .b ({input0_s3[43], input0_s2[43], input0_s1[43], input0_s0[43]}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, new_AGEMA_signal_1990, sbox_inst_10_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_t3_AND_U1 ( .a ({input0_s3[42], input0_s2[42], input0_s1[42], input0_s0[42]}), .b ({input0_s3[43], input0_s2[43], input0_s1[43], input0_s0[43]}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, sbox_inst_10_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_t4_AND_U1 ( .a ({input0_s3[40], input0_s2[40], input0_s1[40], input0_s0[40]}), .b ({input0_s3[41], input0_s2[41], input0_s1[41], input0_s0[41]}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_1998, new_AGEMA_signal_1997, new_AGEMA_signal_1996, sbox_inst_10_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U12 ( .a ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, new_AGEMA_signal_2023, sbox_inst_9_T3}), .b ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, new_AGEMA_signal_2704, sbox_inst_9_n17}), .c ({new_AGEMA_signal_3312, new_AGEMA_signal_3311, new_AGEMA_signal_3310, sbox_inst_9_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U6 ( .a ({new_AGEMA_signal_2028, new_AGEMA_signal_2027, new_AGEMA_signal_2026, sbox_inst_9_T4}), .b ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, sbox_inst_9_T2}), .c ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, new_AGEMA_signal_2698, sbox_inst_9_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U5 ( .a ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, new_AGEMA_signal_2017, sbox_inst_9_T1}), .b ({input0_s3[38], input0_s2[38], input0_s1[38], input0_s0[38]}), .c ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, new_AGEMA_signal_2701, sbox_inst_9_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U4 ( .a ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, new_AGEMA_signal_3319, sbox_inst_9_n11}), .b ({input0_s3[37], input0_s2[37], input0_s1[37], input0_s0[37]}), .c ({output0_s3[9], output0_s2[9], output0_s1[9], output0_s0[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U3 ( .a ({input0_s3[39], input0_s2[39], input0_s1[39], input0_s0[39]}), .b ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, new_AGEMA_signal_2704, sbox_inst_9_n17}), .c ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, new_AGEMA_signal_3319, sbox_inst_9_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U2 ( .a ({input0_s3[36], input0_s2[36], input0_s1[36], input0_s0[36]}), .b ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, new_AGEMA_signal_2008, sbox_inst_9_T0}), .c ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, new_AGEMA_signal_2704, sbox_inst_9_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_t0_AND_U1 ( .a ({input0_s3[37], input0_s2[37], input0_s1[37], input0_s0[37]}), .b ({input0_s3[38], input0_s2[38], input0_s1[38], input0_s0[38]}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, new_AGEMA_signal_2008, sbox_inst_9_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_t1_AND_U1 ( .a ({input0_s3[36], input0_s2[36], input0_s1[36], input0_s0[36]}), .b ({input0_s3[39], input0_s2[39], input0_s1[39], input0_s0[39]}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, new_AGEMA_signal_2017, sbox_inst_9_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_t2_AND_U1 ( .a ({input0_s3[37], input0_s2[37], input0_s1[37], input0_s0[37]}), .b ({input0_s3[39], input0_s2[39], input0_s1[39], input0_s0[39]}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, sbox_inst_9_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_t3_AND_U1 ( .a ({input0_s3[38], input0_s2[38], input0_s1[38], input0_s0[38]}), .b ({input0_s3[39], input0_s2[39], input0_s1[39], input0_s0[39]}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, new_AGEMA_signal_2023, sbox_inst_9_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_t4_AND_U1 ( .a ({input0_s3[36], input0_s2[36], input0_s1[36], input0_s0[36]}), .b ({input0_s3[37], input0_s2[37], input0_s1[37], input0_s0[37]}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_2028, new_AGEMA_signal_2027, new_AGEMA_signal_2026, sbox_inst_9_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U12 ( .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, new_AGEMA_signal_2053, sbox_inst_8_T3}), .b ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, new_AGEMA_signal_2719, sbox_inst_8_n17}), .c ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, new_AGEMA_signal_3325, sbox_inst_8_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U6 ( .a ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, new_AGEMA_signal_2056, sbox_inst_8_T4}), .b ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, new_AGEMA_signal_2050, sbox_inst_8_T2}), .c ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, new_AGEMA_signal_2713, sbox_inst_8_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U5 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, sbox_inst_8_T1}), .b ({input0_s3[34], input0_s2[34], input0_s1[34], input0_s0[34]}), .c ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, new_AGEMA_signal_2716, sbox_inst_8_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U4 ( .a ({new_AGEMA_signal_3336, new_AGEMA_signal_3335, new_AGEMA_signal_3334, sbox_inst_8_n11}), .b ({input0_s3[33], input0_s2[33], input0_s1[33], input0_s0[33]}), .c ({output0_s3[8], output0_s2[8], output0_s1[8], output0_s0[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U3 ( .a ({input0_s3[35], input0_s2[35], input0_s1[35], input0_s0[35]}), .b ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, new_AGEMA_signal_2719, sbox_inst_8_n17}), .c ({new_AGEMA_signal_3336, new_AGEMA_signal_3335, new_AGEMA_signal_3334, sbox_inst_8_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U2 ( .a ({input0_s3[32], input0_s2[32], input0_s1[32], input0_s0[32]}), .b ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, sbox_inst_8_T0}), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, new_AGEMA_signal_2719, sbox_inst_8_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_t0_AND_U1 ( .a ({input0_s3[33], input0_s2[33], input0_s1[33], input0_s0[33]}), .b ({input0_s3[34], input0_s2[34], input0_s1[34], input0_s0[34]}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, new_AGEMA_signal_2038, sbox_inst_8_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_t1_AND_U1 ( .a ({input0_s3[32], input0_s2[32], input0_s1[32], input0_s0[32]}), .b ({input0_s3[35], input0_s2[35], input0_s1[35], input0_s0[35]}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, sbox_inst_8_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_t2_AND_U1 ( .a ({input0_s3[33], input0_s2[33], input0_s1[33], input0_s0[33]}), .b ({input0_s3[35], input0_s2[35], input0_s1[35], input0_s0[35]}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, new_AGEMA_signal_2050, sbox_inst_8_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_t3_AND_U1 ( .a ({input0_s3[34], input0_s2[34], input0_s1[34], input0_s0[34]}), .b ({input0_s3[35], input0_s2[35], input0_s1[35], input0_s0[35]}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, new_AGEMA_signal_2053, sbox_inst_8_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_t4_AND_U1 ( .a ({input0_s3[32], input0_s2[32], input0_s1[32], input0_s0[32]}), .b ({input0_s3[33], input0_s2[33], input0_s1[33], input0_s0[33]}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, new_AGEMA_signal_2056, sbox_inst_8_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U12 ( .a ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, sbox_inst_7_T3}), .b ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, new_AGEMA_signal_2734, sbox_inst_7_n17}), .c ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, new_AGEMA_signal_3340, sbox_inst_7_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U6 ( .a ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, sbox_inst_7_T4}), .b ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, sbox_inst_7_T2}), .c ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, new_AGEMA_signal_2728, sbox_inst_7_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U5 ( .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, new_AGEMA_signal_2077, sbox_inst_7_T1}), .b ({input0_s3[30], input0_s2[30], input0_s1[30], input0_s0[30]}), .c ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, new_AGEMA_signal_2731, sbox_inst_7_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U4 ( .a ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, new_AGEMA_signal_3349, sbox_inst_7_n11}), .b ({input0_s3[29], input0_s2[29], input0_s1[29], input0_s0[29]}), .c ({output0_s3[7], output0_s2[7], output0_s1[7], output0_s0[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U3 ( .a ({input0_s3[31], input0_s2[31], input0_s1[31], input0_s0[31]}), .b ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, new_AGEMA_signal_2734, sbox_inst_7_n17}), .c ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, new_AGEMA_signal_3349, sbox_inst_7_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U2 ( .a ({input0_s3[28], input0_s2[28], input0_s1[28], input0_s0[28]}), .b ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, new_AGEMA_signal_2068, sbox_inst_7_T0}), .c ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, new_AGEMA_signal_2734, sbox_inst_7_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_t0_AND_U1 ( .a ({input0_s3[29], input0_s2[29], input0_s1[29], input0_s0[29]}), .b ({input0_s3[30], input0_s2[30], input0_s1[30], input0_s0[30]}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, new_AGEMA_signal_2068, sbox_inst_7_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_t1_AND_U1 ( .a ({input0_s3[28], input0_s2[28], input0_s1[28], input0_s0[28]}), .b ({input0_s3[31], input0_s2[31], input0_s1[31], input0_s0[31]}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, new_AGEMA_signal_2077, sbox_inst_7_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_t2_AND_U1 ( .a ({input0_s3[29], input0_s2[29], input0_s1[29], input0_s0[29]}), .b ({input0_s3[31], input0_s2[31], input0_s1[31], input0_s0[31]}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, sbox_inst_7_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_t3_AND_U1 ( .a ({input0_s3[30], input0_s2[30], input0_s1[30], input0_s0[30]}), .b ({input0_s3[31], input0_s2[31], input0_s1[31], input0_s0[31]}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, sbox_inst_7_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_t4_AND_U1 ( .a ({input0_s3[28], input0_s2[28], input0_s1[28], input0_s0[28]}), .b ({input0_s3[29], input0_s2[29], input0_s1[29], input0_s0[29]}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, new_AGEMA_signal_2086, sbox_inst_7_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U12 ( .a ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, sbox_inst_6_T3}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, new_AGEMA_signal_2749, sbox_inst_6_n17}), .c ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, new_AGEMA_signal_3355, sbox_inst_6_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U6 ( .a ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, new_AGEMA_signal_2116, sbox_inst_6_T4}), .b ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, sbox_inst_6_T2}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, new_AGEMA_signal_2743, sbox_inst_6_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U5 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, sbox_inst_6_T1}), .b ({input0_s3[26], input0_s2[26], input0_s1[26], input0_s0[26]}), .c ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, new_AGEMA_signal_2746, sbox_inst_6_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U4 ( .a ({new_AGEMA_signal_3366, new_AGEMA_signal_3365, new_AGEMA_signal_3364, sbox_inst_6_n11}), .b ({input0_s3[25], input0_s2[25], input0_s1[25], input0_s0[25]}), .c ({output0_s3[6], output0_s2[6], output0_s1[6], output0_s0[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U3 ( .a ({input0_s3[27], input0_s2[27], input0_s1[27], input0_s0[27]}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, new_AGEMA_signal_2749, sbox_inst_6_n17}), .c ({new_AGEMA_signal_3366, new_AGEMA_signal_3365, new_AGEMA_signal_3364, sbox_inst_6_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U2 ( .a ({input0_s3[24], input0_s2[24], input0_s1[24], input0_s0[24]}), .b ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, sbox_inst_6_T0}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, new_AGEMA_signal_2749, sbox_inst_6_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_t0_AND_U1 ( .a ({input0_s3[25], input0_s2[25], input0_s1[25], input0_s0[25]}), .b ({input0_s3[26], input0_s2[26], input0_s1[26], input0_s0[26]}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, new_AGEMA_signal_2098, sbox_inst_6_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_t1_AND_U1 ( .a ({input0_s3[24], input0_s2[24], input0_s1[24], input0_s0[24]}), .b ({input0_s3[27], input0_s2[27], input0_s1[27], input0_s0[27]}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, sbox_inst_6_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_t2_AND_U1 ( .a ({input0_s3[25], input0_s2[25], input0_s1[25], input0_s0[25]}), .b ({input0_s3[27], input0_s2[27], input0_s1[27], input0_s0[27]}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, sbox_inst_6_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_t3_AND_U1 ( .a ({input0_s3[26], input0_s2[26], input0_s1[26], input0_s0[26]}), .b ({input0_s3[27], input0_s2[27], input0_s1[27], input0_s0[27]}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, sbox_inst_6_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_t4_AND_U1 ( .a ({input0_s3[24], input0_s2[24], input0_s1[24], input0_s0[24]}), .b ({input0_s3[25], input0_s2[25], input0_s1[25], input0_s0[25]}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, new_AGEMA_signal_2116, sbox_inst_6_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U12 ( .a ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, sbox_inst_5_T3}), .b ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, new_AGEMA_signal_2764, sbox_inst_5_n17}), .c ({new_AGEMA_signal_3372, new_AGEMA_signal_3371, new_AGEMA_signal_3370, sbox_inst_5_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U6 ( .a ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, sbox_inst_5_T4}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, new_AGEMA_signal_2140, sbox_inst_5_T2}), .c ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, new_AGEMA_signal_2758, sbox_inst_5_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U5 ( .a ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, sbox_inst_5_T1}), .b ({input0_s3[22], input0_s2[22], input0_s1[22], input0_s0[22]}), .c ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, new_AGEMA_signal_2761, sbox_inst_5_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U4 ( .a ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, new_AGEMA_signal_3379, sbox_inst_5_n11}), .b ({input0_s3[21], input0_s2[21], input0_s1[21], input0_s0[21]}), .c ({output0_s3[5], output0_s2[5], output0_s1[5], output0_s0[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U3 ( .a ({input0_s3[23], input0_s2[23], input0_s1[23], input0_s0[23]}), .b ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, new_AGEMA_signal_2764, sbox_inst_5_n17}), .c ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, new_AGEMA_signal_3379, sbox_inst_5_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U2 ( .a ({input0_s3[20], input0_s2[20], input0_s1[20], input0_s0[20]}), .b ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, new_AGEMA_signal_2128, sbox_inst_5_T0}), .c ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, new_AGEMA_signal_2764, sbox_inst_5_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_t0_AND_U1 ( .a ({input0_s3[21], input0_s2[21], input0_s1[21], input0_s0[21]}), .b ({input0_s3[22], input0_s2[22], input0_s1[22], input0_s0[22]}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, new_AGEMA_signal_2128, sbox_inst_5_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_t1_AND_U1 ( .a ({input0_s3[20], input0_s2[20], input0_s1[20], input0_s0[20]}), .b ({input0_s3[23], input0_s2[23], input0_s1[23], input0_s0[23]}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, sbox_inst_5_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_t2_AND_U1 ( .a ({input0_s3[21], input0_s2[21], input0_s1[21], input0_s0[21]}), .b ({input0_s3[23], input0_s2[23], input0_s1[23], input0_s0[23]}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, new_AGEMA_signal_2140, sbox_inst_5_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_t3_AND_U1 ( .a ({input0_s3[22], input0_s2[22], input0_s1[22], input0_s0[22]}), .b ({input0_s3[23], input0_s2[23], input0_s1[23], input0_s0[23]}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, sbox_inst_5_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_t4_AND_U1 ( .a ({input0_s3[20], input0_s2[20], input0_s1[20], input0_s0[20]}), .b ({input0_s3[21], input0_s2[21], input0_s1[21], input0_s0[21]}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, new_AGEMA_signal_2146, sbox_inst_5_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U12 ( .a ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, new_AGEMA_signal_2173, sbox_inst_4_T3}), .b ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, new_AGEMA_signal_2779, sbox_inst_4_n17}), .c ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, new_AGEMA_signal_3385, sbox_inst_4_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U6 ( .a ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, new_AGEMA_signal_2176, sbox_inst_4_T4}), .b ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, sbox_inst_4_T2}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, new_AGEMA_signal_2773, sbox_inst_4_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U5 ( .a ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, sbox_inst_4_T1}), .b ({input0_s3[18], input0_s2[18], input0_s1[18], input0_s0[18]}), .c ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, new_AGEMA_signal_2776, sbox_inst_4_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U4 ( .a ({new_AGEMA_signal_3396, new_AGEMA_signal_3395, new_AGEMA_signal_3394, sbox_inst_4_n11}), .b ({input0_s3[17], input0_s2[17], input0_s1[17], input0_s0[17]}), .c ({output0_s3[4], output0_s2[4], output0_s1[4], output0_s0[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U3 ( .a ({input0_s3[19], input0_s2[19], input0_s1[19], input0_s0[19]}), .b ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, new_AGEMA_signal_2779, sbox_inst_4_n17}), .c ({new_AGEMA_signal_3396, new_AGEMA_signal_3395, new_AGEMA_signal_3394, sbox_inst_4_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U2 ( .a ({input0_s3[16], input0_s2[16], input0_s1[16], input0_s0[16]}), .b ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, sbox_inst_4_T0}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, new_AGEMA_signal_2779, sbox_inst_4_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_t0_AND_U1 ( .a ({input0_s3[17], input0_s2[17], input0_s1[17], input0_s0[17]}), .b ({input0_s3[18], input0_s2[18], input0_s1[18], input0_s0[18]}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, new_AGEMA_signal_2158, sbox_inst_4_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_t1_AND_U1 ( .a ({input0_s3[16], input0_s2[16], input0_s1[16], input0_s0[16]}), .b ({input0_s3[19], input0_s2[19], input0_s1[19], input0_s0[19]}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, sbox_inst_4_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_t2_AND_U1 ( .a ({input0_s3[17], input0_s2[17], input0_s1[17], input0_s0[17]}), .b ({input0_s3[19], input0_s2[19], input0_s1[19], input0_s0[19]}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, sbox_inst_4_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_t3_AND_U1 ( .a ({input0_s3[18], input0_s2[18], input0_s1[18], input0_s0[18]}), .b ({input0_s3[19], input0_s2[19], input0_s1[19], input0_s0[19]}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, new_AGEMA_signal_2173, sbox_inst_4_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_t4_AND_U1 ( .a ({input0_s3[16], input0_s2[16], input0_s1[16], input0_s0[16]}), .b ({input0_s3[17], input0_s2[17], input0_s1[17], input0_s0[17]}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, new_AGEMA_signal_2176, sbox_inst_4_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U12 ( .a ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, new_AGEMA_signal_2203, sbox_inst_3_T3}), .b ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, new_AGEMA_signal_2794, sbox_inst_3_n17}), .c ({new_AGEMA_signal_3402, new_AGEMA_signal_3401, new_AGEMA_signal_3400, sbox_inst_3_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U6 ( .a ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, sbox_inst_3_T4}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, new_AGEMA_signal_2200, sbox_inst_3_T2}), .c ({new_AGEMA_signal_2790, new_AGEMA_signal_2789, new_AGEMA_signal_2788, sbox_inst_3_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U5 ( .a ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, new_AGEMA_signal_2197, sbox_inst_3_T1}), .b ({input0_s3[14], input0_s2[14], input0_s1[14], input0_s0[14]}), .c ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, new_AGEMA_signal_2791, sbox_inst_3_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U4 ( .a ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, new_AGEMA_signal_3409, sbox_inst_3_n11}), .b ({input0_s3[13], input0_s2[13], input0_s1[13], input0_s0[13]}), .c ({output0_s3[3], output0_s2[3], output0_s1[3], output0_s0[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U3 ( .a ({input0_s3[15], input0_s2[15], input0_s1[15], input0_s0[15]}), .b ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, new_AGEMA_signal_2794, sbox_inst_3_n17}), .c ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, new_AGEMA_signal_3409, sbox_inst_3_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U2 ( .a ({input0_s3[12], input0_s2[12], input0_s1[12], input0_s0[12]}), .b ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, new_AGEMA_signal_2188, sbox_inst_3_T0}), .c ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, new_AGEMA_signal_2794, sbox_inst_3_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_t0_AND_U1 ( .a ({input0_s3[13], input0_s2[13], input0_s1[13], input0_s0[13]}), .b ({input0_s3[14], input0_s2[14], input0_s1[14], input0_s0[14]}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, new_AGEMA_signal_2188, sbox_inst_3_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_t1_AND_U1 ( .a ({input0_s3[12], input0_s2[12], input0_s1[12], input0_s0[12]}), .b ({input0_s3[15], input0_s2[15], input0_s1[15], input0_s0[15]}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, new_AGEMA_signal_2197, sbox_inst_3_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_t2_AND_U1 ( .a ({input0_s3[13], input0_s2[13], input0_s1[13], input0_s0[13]}), .b ({input0_s3[15], input0_s2[15], input0_s1[15], input0_s0[15]}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, new_AGEMA_signal_2200, sbox_inst_3_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_t3_AND_U1 ( .a ({input0_s3[14], input0_s2[14], input0_s1[14], input0_s0[14]}), .b ({input0_s3[15], input0_s2[15], input0_s1[15], input0_s0[15]}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, new_AGEMA_signal_2203, sbox_inst_3_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_t4_AND_U1 ( .a ({input0_s3[12], input0_s2[12], input0_s1[12], input0_s0[12]}), .b ({input0_s3[13], input0_s2[13], input0_s1[13], input0_s0[13]}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, new_AGEMA_signal_2206, sbox_inst_3_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U12 ( .a ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, sbox_inst_2_T3}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, new_AGEMA_signal_2809, sbox_inst_2_n17}), .c ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, new_AGEMA_signal_3415, sbox_inst_2_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U6 ( .a ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, new_AGEMA_signal_2236, sbox_inst_2_T4}), .b ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, sbox_inst_2_T2}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, new_AGEMA_signal_2803, sbox_inst_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U5 ( .a ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, new_AGEMA_signal_2227, sbox_inst_2_T1}), .b ({input0_s3[10], input0_s2[10], input0_s1[10], input0_s0[10]}), .c ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, new_AGEMA_signal_2806, sbox_inst_2_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U4 ( .a ({new_AGEMA_signal_3426, new_AGEMA_signal_3425, new_AGEMA_signal_3424, sbox_inst_2_n11}), .b ({input0_s3[9], input0_s2[9], input0_s1[9], input0_s0[9]}), .c ({output0_s3[2], output0_s2[2], output0_s1[2], output0_s0[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U3 ( .a ({input0_s3[11], input0_s2[11], input0_s1[11], input0_s0[11]}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, new_AGEMA_signal_2809, sbox_inst_2_n17}), .c ({new_AGEMA_signal_3426, new_AGEMA_signal_3425, new_AGEMA_signal_3424, sbox_inst_2_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U2 ( .a ({input0_s3[8], input0_s2[8], input0_s1[8], input0_s0[8]}), .b ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, sbox_inst_2_T0}), .c ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, new_AGEMA_signal_2809, sbox_inst_2_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_t0_AND_U1 ( .a ({input0_s3[9], input0_s2[9], input0_s1[9], input0_s0[9]}), .b ({input0_s3[10], input0_s2[10], input0_s1[10], input0_s0[10]}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, new_AGEMA_signal_2218, sbox_inst_2_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_t1_AND_U1 ( .a ({input0_s3[8], input0_s2[8], input0_s1[8], input0_s0[8]}), .b ({input0_s3[11], input0_s2[11], input0_s1[11], input0_s0[11]}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, new_AGEMA_signal_2227, sbox_inst_2_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_t2_AND_U1 ( .a ({input0_s3[9], input0_s2[9], input0_s1[9], input0_s0[9]}), .b ({input0_s3[11], input0_s2[11], input0_s1[11], input0_s0[11]}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, sbox_inst_2_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_t3_AND_U1 ( .a ({input0_s3[10], input0_s2[10], input0_s1[10], input0_s0[10]}), .b ({input0_s3[11], input0_s2[11], input0_s1[11], input0_s0[11]}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, sbox_inst_2_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_t4_AND_U1 ( .a ({input0_s3[8], input0_s2[8], input0_s1[8], input0_s0[8]}), .b ({input0_s3[9], input0_s2[9], input0_s1[9], input0_s0[9]}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, new_AGEMA_signal_2236, sbox_inst_2_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U12 ( .a ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, new_AGEMA_signal_2833, sbox_inst_1_T3}), .b ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, new_AGEMA_signal_3433, sbox_inst_1_n17}), .c ({new_AGEMA_signal_3924, new_AGEMA_signal_3923, new_AGEMA_signal_3922, sbox_inst_1_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U6 ( .a ({new_AGEMA_signal_2838, new_AGEMA_signal_2837, new_AGEMA_signal_2836, sbox_inst_1_T4}), .b ({new_AGEMA_signal_2832, new_AGEMA_signal_2831, new_AGEMA_signal_2830, sbox_inst_1_T2}), .c ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, new_AGEMA_signal_3427, sbox_inst_1_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U5 ( .a ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, new_AGEMA_signal_2827, sbox_inst_1_T1}), .b ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, input_array_6}), .c ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, new_AGEMA_signal_3430, sbox_inst_1_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U4 ( .a ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, new_AGEMA_signal_3931, sbox_inst_1_n11}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, input_array_5}), .c ({output0_s3[1], output0_s2[1], output0_s1[1], output0_s0[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U3 ( .a ({input0_s3[7], input0_s2[7], input0_s1[7], input0_s0[7]}), .b ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, new_AGEMA_signal_3433, sbox_inst_1_n17}), .c ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, new_AGEMA_signal_3931, sbox_inst_1_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U2 ( .a ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, new_AGEMA_signal_1108, input_array_4}), .b ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, new_AGEMA_signal_2821, sbox_inst_1_T0}), .c ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, new_AGEMA_signal_3433, sbox_inst_1_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_t0_AND_U1 ( .a ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, input_array_5}), .b ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, input_array_6}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, new_AGEMA_signal_2821, sbox_inst_1_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_t1_AND_U1 ( .a ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, new_AGEMA_signal_1108, input_array_4}), .b ({input0_s3[7], input0_s2[7], input0_s1[7], input0_s0[7]}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, new_AGEMA_signal_2827, sbox_inst_1_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_t2_AND_U1 ( .a ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, input_array_5}), .b ({input0_s3[7], input0_s2[7], input0_s1[7], input0_s0[7]}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_2832, new_AGEMA_signal_2831, new_AGEMA_signal_2830, sbox_inst_1_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_t3_AND_U1 ( .a ({new_AGEMA_signal_1104, new_AGEMA_signal_1103, new_AGEMA_signal_1102, input_array_6}), .b ({input0_s3[7], input0_s2[7], input0_s1[7], input0_s0[7]}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, new_AGEMA_signal_2833, sbox_inst_1_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_t4_AND_U1 ( .a ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, new_AGEMA_signal_1108, input_array_4}), .b ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, input_array_5}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_2838, new_AGEMA_signal_2837, new_AGEMA_signal_2836, sbox_inst_1_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U12 ( .a ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, new_AGEMA_signal_2851, sbox_inst_0_T3}), .b ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, new_AGEMA_signal_3448, sbox_inst_0_n17}), .c ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, new_AGEMA_signal_3937, sbox_inst_0_n19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U6 ( .a ({new_AGEMA_signal_2856, new_AGEMA_signal_2855, new_AGEMA_signal_2854, sbox_inst_0_T4}), .b ({new_AGEMA_signal_2850, new_AGEMA_signal_2849, new_AGEMA_signal_2848, sbox_inst_0_T2}), .c ({new_AGEMA_signal_3444, new_AGEMA_signal_3443, new_AGEMA_signal_3442, sbox_inst_0_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U5 ( .a ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, new_AGEMA_signal_2845, sbox_inst_0_T1}), .b ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, new_AGEMA_signal_1120, input_array_2}), .c ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, new_AGEMA_signal_3445, sbox_inst_0_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U4 ( .a ({new_AGEMA_signal_3948, new_AGEMA_signal_3947, new_AGEMA_signal_3946, sbox_inst_0_n11}), .b ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, input_array_1}), .c ({output0_s3[0], output0_s2[0], output0_s1[0], output0_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U3 ( .a ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, new_AGEMA_signal_1114, input_array_3}), .b ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, new_AGEMA_signal_3448, sbox_inst_0_n17}), .c ({new_AGEMA_signal_3948, new_AGEMA_signal_3947, new_AGEMA_signal_3946, sbox_inst_0_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U2 ( .a ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, input_array_0}), .b ({new_AGEMA_signal_2844, new_AGEMA_signal_2843, new_AGEMA_signal_2842, sbox_inst_0_T0}), .c ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, new_AGEMA_signal_3448, sbox_inst_0_n17}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_t0_AND_U1 ( .a ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, input_array_1}), .b ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, new_AGEMA_signal_1120, input_array_2}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_2844, new_AGEMA_signal_2843, new_AGEMA_signal_2842, sbox_inst_0_T0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_t1_AND_U1 ( .a ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, input_array_0}), .b ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, new_AGEMA_signal_1114, input_array_3}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, new_AGEMA_signal_2845, sbox_inst_0_T1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_t2_AND_U1 ( .a ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, input_array_1}), .b ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, new_AGEMA_signal_1114, input_array_3}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_2850, new_AGEMA_signal_2849, new_AGEMA_signal_2848, sbox_inst_0_T2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_t3_AND_U1 ( .a ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, new_AGEMA_signal_1120, input_array_2}), .b ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, new_AGEMA_signal_1114, input_array_3}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, new_AGEMA_signal_2851, sbox_inst_0_T3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_t4_AND_U1 ( .a ({new_AGEMA_signal_1128, new_AGEMA_signal_1127, new_AGEMA_signal_1126, input_array_0}), .b ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, input_array_1}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_2856, new_AGEMA_signal_2855, new_AGEMA_signal_2854, sbox_inst_0_T4}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U15 ( .a ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, new_AGEMA_signal_2248, sbox_inst_39_T2}), .b ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, new_AGEMA_signal_3949, sbox_inst_39_n20}), .c ({output0_s3[79], output0_s2[79], output0_s1[79], output0_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U14 ( .a ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, new_AGEMA_signal_3460, sbox_inst_39_n19}), .b ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, new_AGEMA_signal_3457, sbox_inst_39_n18}), .c ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, new_AGEMA_signal_3949, sbox_inst_39_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U13 ( .a ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, new_AGEMA_signal_2245, sbox_inst_39_T1}), .b ({new_AGEMA_signal_2868, new_AGEMA_signal_2867, new_AGEMA_signal_2866, sbox_inst_39_T5}), .c ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, new_AGEMA_signal_3457, sbox_inst_39_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U11 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, input_array[157]}), .b ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, new_AGEMA_signal_3463, sbox_inst_39_n16}), .c ({output0_s3[119], output0_s2[119], output0_s1[119], output0_s0[119]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U10 ( .a ({new_AGEMA_signal_2862, new_AGEMA_signal_2861, new_AGEMA_signal_2860, sbox_inst_39_n15}), .b ({new_AGEMA_signal_2868, new_AGEMA_signal_2867, new_AGEMA_signal_2866, sbox_inst_39_T5}), .c ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, new_AGEMA_signal_3463, sbox_inst_39_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U9 ( .a ({new_AGEMA_signal_2862, new_AGEMA_signal_2861, new_AGEMA_signal_2860, sbox_inst_39_n15}), .b ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, new_AGEMA_signal_3955, sbox_inst_39_n14}), .c ({output0_s3[159], output0_s2[159], output0_s1[159], output0_s0[159]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U8 ( .a ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, new_AGEMA_signal_2857, sbox_inst_39_n13}), .b ({new_AGEMA_signal_3468, new_AGEMA_signal_3467, new_AGEMA_signal_3466, sbox_inst_39_n12}), .c ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, new_AGEMA_signal_3955, sbox_inst_39_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_U7 ( .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, new_AGEMA_signal_2869, sbox_inst_39_T6}), .b ({new_AGEMA_signal_1134, new_AGEMA_signal_1133, new_AGEMA_signal_1132, input_array[159]}), .c ({new_AGEMA_signal_3468, new_AGEMA_signal_3467, new_AGEMA_signal_3466, sbox_inst_39_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_t5_AND_U1 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, new_AGEMA_signal_1084, input_array[157]}), .b ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, new_AGEMA_signal_2251, sbox_inst_39_T3}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_2868, new_AGEMA_signal_2867, new_AGEMA_signal_2866, sbox_inst_39_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_39_t6_AND_U1 ( .a ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, new_AGEMA_signal_2239, sbox_inst_39_L0}), .b ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, new_AGEMA_signal_2245, sbox_inst_39_T1}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, new_AGEMA_signal_2869, sbox_inst_39_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U15 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, new_AGEMA_signal_2269, sbox_inst_38_T2}), .b ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, new_AGEMA_signal_3961, sbox_inst_38_n20}), .c ({output0_s3[78], output0_s2[78], output0_s1[78], output0_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U14 ( .a ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, new_AGEMA_signal_3475, sbox_inst_38_n19}), .b ({new_AGEMA_signal_3474, new_AGEMA_signal_3473, new_AGEMA_signal_3472, sbox_inst_38_n18}), .c ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, new_AGEMA_signal_3961, sbox_inst_38_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U13 ( .a ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, sbox_inst_38_T1}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, new_AGEMA_signal_2881, sbox_inst_38_T5}), .c ({new_AGEMA_signal_3474, new_AGEMA_signal_3473, new_AGEMA_signal_3472, sbox_inst_38_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U11 ( .a ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, input_array[153]}), .b ({new_AGEMA_signal_3480, new_AGEMA_signal_3479, new_AGEMA_signal_3478, sbox_inst_38_n16}), .c ({output0_s3[118], output0_s2[118], output0_s1[118], output0_s0[118]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U10 ( .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, new_AGEMA_signal_2875, sbox_inst_38_n15}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, new_AGEMA_signal_2881, sbox_inst_38_T5}), .c ({new_AGEMA_signal_3480, new_AGEMA_signal_3479, new_AGEMA_signal_3478, sbox_inst_38_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U9 ( .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, new_AGEMA_signal_2875, sbox_inst_38_n15}), .b ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, new_AGEMA_signal_3967, sbox_inst_38_n14}), .c ({output0_s3[158], output0_s2[158], output0_s1[158], output0_s0[158]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U8 ( .a ({new_AGEMA_signal_2874, new_AGEMA_signal_2873, new_AGEMA_signal_2872, sbox_inst_38_n13}), .b ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, new_AGEMA_signal_3481, sbox_inst_38_n12}), .c ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, new_AGEMA_signal_3967, sbox_inst_38_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_U7 ( .a ({new_AGEMA_signal_2886, new_AGEMA_signal_2885, new_AGEMA_signal_2884, sbox_inst_38_T6}), .b ({new_AGEMA_signal_1152, new_AGEMA_signal_1151, new_AGEMA_signal_1150, input_array[155]}), .c ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, new_AGEMA_signal_3481, sbox_inst_38_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_t5_AND_U1 ( .a ({new_AGEMA_signal_1092, new_AGEMA_signal_1091, new_AGEMA_signal_1090, input_array[153]}), .b ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, new_AGEMA_signal_2272, sbox_inst_38_T3}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, new_AGEMA_signal_2881, sbox_inst_38_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_38_t6_AND_U1 ( .a ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, new_AGEMA_signal_2257, sbox_inst_38_L0}), .b ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, new_AGEMA_signal_2266, sbox_inst_38_T1}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_2886, new_AGEMA_signal_2885, new_AGEMA_signal_2884, sbox_inst_38_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U15 ( .a ({new_AGEMA_signal_1182, new_AGEMA_signal_1181, new_AGEMA_signal_1180, sbox_inst_37_T2}), .b ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, new_AGEMA_signal_3487, sbox_inst_37_n20}), .c ({output0_s3[77], output0_s2[77], output0_s1[77], output0_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U14 ( .a ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, new_AGEMA_signal_2890, sbox_inst_37_n19}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, new_AGEMA_signal_2887, sbox_inst_37_n18}), .c ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, new_AGEMA_signal_3487, sbox_inst_37_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U13 ( .a ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, new_AGEMA_signal_1177, sbox_inst_37_T1}), .b ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, sbox_inst_37_T5}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, new_AGEMA_signal_2887, sbox_inst_37_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U11 ( .a ({input0_s3[149], input0_s2[149], input0_s1[149], input0_s0[149]}), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, new_AGEMA_signal_2893, sbox_inst_37_n16}), .c ({output0_s3[117], output0_s2[117], output0_s1[117], output0_s0[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U10 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, sbox_inst_37_n15}), .b ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, sbox_inst_37_T5}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, new_AGEMA_signal_2893, sbox_inst_37_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U9 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, new_AGEMA_signal_2281, sbox_inst_37_n15}), .b ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, new_AGEMA_signal_3493, sbox_inst_37_n14}), .c ({output0_s3[157], output0_s2[157], output0_s1[157], output0_s0[157]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U8 ( .a ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, new_AGEMA_signal_2278, sbox_inst_37_n13}), .b ({new_AGEMA_signal_2898, new_AGEMA_signal_2897, new_AGEMA_signal_2896, sbox_inst_37_n12}), .c ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, new_AGEMA_signal_3493, sbox_inst_37_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_U7 ( .a ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, sbox_inst_37_T6}), .b ({input0_s3[151], input0_s2[151], input0_s1[151], input0_s0[151]}), .c ({new_AGEMA_signal_2898, new_AGEMA_signal_2897, new_AGEMA_signal_2896, sbox_inst_37_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_t5_AND_U1 ( .a ({input0_s3[149], input0_s2[149], input0_s1[149], input0_s0[149]}), .b ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, new_AGEMA_signal_1183, sbox_inst_37_T3}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, new_AGEMA_signal_2287, sbox_inst_37_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_37_t6_AND_U1 ( .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, new_AGEMA_signal_1165, sbox_inst_37_L0}), .b ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, new_AGEMA_signal_1177, sbox_inst_37_T1}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, new_AGEMA_signal_2290, sbox_inst_37_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U15 ( .a ({new_AGEMA_signal_1212, new_AGEMA_signal_1211, new_AGEMA_signal_1210, sbox_inst_36_T2}), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, new_AGEMA_signal_3499, sbox_inst_36_n20}), .c ({output0_s3[76], output0_s2[76], output0_s1[76], output0_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U14 ( .a ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, new_AGEMA_signal_2905, sbox_inst_36_n19}), .b ({new_AGEMA_signal_2904, new_AGEMA_signal_2903, new_AGEMA_signal_2902, sbox_inst_36_n18}), .c ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, new_AGEMA_signal_3499, sbox_inst_36_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U13 ( .a ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, sbox_inst_36_T1}), .b ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, sbox_inst_36_T5}), .c ({new_AGEMA_signal_2904, new_AGEMA_signal_2903, new_AGEMA_signal_2902, sbox_inst_36_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U11 ( .a ({input0_s3[145], input0_s2[145], input0_s1[145], input0_s0[145]}), .b ({new_AGEMA_signal_2910, new_AGEMA_signal_2909, new_AGEMA_signal_2908, sbox_inst_36_n16}), .c ({output0_s3[116], output0_s2[116], output0_s1[116], output0_s0[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U10 ( .a ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, new_AGEMA_signal_2296, sbox_inst_36_n15}), .b ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, sbox_inst_36_T5}), .c ({new_AGEMA_signal_2910, new_AGEMA_signal_2909, new_AGEMA_signal_2908, sbox_inst_36_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U9 ( .a ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, new_AGEMA_signal_2296, sbox_inst_36_n15}), .b ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, new_AGEMA_signal_3505, sbox_inst_36_n14}), .c ({output0_s3[156], output0_s2[156], output0_s1[156], output0_s0[156]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U8 ( .a ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, new_AGEMA_signal_2293, sbox_inst_36_n13}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, new_AGEMA_signal_2911, sbox_inst_36_n12}), .c ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, new_AGEMA_signal_3505, sbox_inst_36_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_U7 ( .a ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, new_AGEMA_signal_2305, sbox_inst_36_T6}), .b ({input0_s3[147], input0_s2[147], input0_s1[147], input0_s0[147]}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, new_AGEMA_signal_2911, sbox_inst_36_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_t5_AND_U1 ( .a ({input0_s3[145], input0_s2[145], input0_s1[145], input0_s0[145]}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, new_AGEMA_signal_1213, sbox_inst_36_T3}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, new_AGEMA_signal_2302, sbox_inst_36_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_36_t6_AND_U1 ( .a ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, new_AGEMA_signal_1195, sbox_inst_36_L0}), .b ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, new_AGEMA_signal_1207, sbox_inst_36_T1}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, new_AGEMA_signal_2305, sbox_inst_36_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U15 ( .a ({new_AGEMA_signal_1242, new_AGEMA_signal_1241, new_AGEMA_signal_1240, sbox_inst_35_T2}), .b ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, new_AGEMA_signal_3511, sbox_inst_35_n20}), .c ({output0_s3[75], output0_s2[75], output0_s1[75], output0_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U14 ( .a ({new_AGEMA_signal_2922, new_AGEMA_signal_2921, new_AGEMA_signal_2920, sbox_inst_35_n19}), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, new_AGEMA_signal_2917, sbox_inst_35_n18}), .c ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, new_AGEMA_signal_3511, sbox_inst_35_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U13 ( .a ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, new_AGEMA_signal_1237, sbox_inst_35_T1}), .b ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, new_AGEMA_signal_2317, sbox_inst_35_T5}), .c ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, new_AGEMA_signal_2917, sbox_inst_35_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U11 ( .a ({input0_s3[141], input0_s2[141], input0_s1[141], input0_s0[141]}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, new_AGEMA_signal_2923, sbox_inst_35_n16}), .c ({output0_s3[115], output0_s2[115], output0_s1[115], output0_s0[115]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U10 ( .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, sbox_inst_35_n15}), .b ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, new_AGEMA_signal_2317, sbox_inst_35_T5}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, new_AGEMA_signal_2923, sbox_inst_35_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U9 ( .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, new_AGEMA_signal_2311, sbox_inst_35_n15}), .b ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, new_AGEMA_signal_3517, sbox_inst_35_n14}), .c ({output0_s3[155], output0_s2[155], output0_s1[155], output0_s0[155]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U8 ( .a ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, new_AGEMA_signal_2308, sbox_inst_35_n13}), .b ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, new_AGEMA_signal_2926, sbox_inst_35_n12}), .c ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, new_AGEMA_signal_3517, sbox_inst_35_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_U7 ( .a ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, new_AGEMA_signal_2320, sbox_inst_35_T6}), .b ({input0_s3[143], input0_s2[143], input0_s1[143], input0_s0[143]}), .c ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, new_AGEMA_signal_2926, sbox_inst_35_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_t5_AND_U1 ( .a ({input0_s3[141], input0_s2[141], input0_s1[141], input0_s0[141]}), .b ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, new_AGEMA_signal_1243, sbox_inst_35_T3}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, new_AGEMA_signal_2317, sbox_inst_35_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_35_t6_AND_U1 ( .a ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, new_AGEMA_signal_1225, sbox_inst_35_L0}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, new_AGEMA_signal_1237, sbox_inst_35_T1}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, new_AGEMA_signal_2320, sbox_inst_35_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U15 ( .a ({new_AGEMA_signal_1272, new_AGEMA_signal_1271, new_AGEMA_signal_1270, sbox_inst_34_T2}), .b ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, new_AGEMA_signal_3523, sbox_inst_34_n20}), .c ({output0_s3[74], output0_s2[74], output0_s1[74], output0_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U14 ( .a ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, new_AGEMA_signal_2935, sbox_inst_34_n19}), .b ({new_AGEMA_signal_2934, new_AGEMA_signal_2933, new_AGEMA_signal_2932, sbox_inst_34_n18}), .c ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, new_AGEMA_signal_3523, sbox_inst_34_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U13 ( .a ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, sbox_inst_34_T1}), .b ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, new_AGEMA_signal_2332, sbox_inst_34_T5}), .c ({new_AGEMA_signal_2934, new_AGEMA_signal_2933, new_AGEMA_signal_2932, sbox_inst_34_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U11 ( .a ({input0_s3[137], input0_s2[137], input0_s1[137], input0_s0[137]}), .b ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, new_AGEMA_signal_2938, sbox_inst_34_n16}), .c ({output0_s3[114], output0_s2[114], output0_s1[114], output0_s0[114]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U10 ( .a ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, sbox_inst_34_n15}), .b ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, new_AGEMA_signal_2332, sbox_inst_34_T5}), .c ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, new_AGEMA_signal_2938, sbox_inst_34_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U9 ( .a ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, new_AGEMA_signal_2326, sbox_inst_34_n15}), .b ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, new_AGEMA_signal_3529, sbox_inst_34_n14}), .c ({output0_s3[154], output0_s2[154], output0_s1[154], output0_s0[154]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U8 ( .a ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, new_AGEMA_signal_2323, sbox_inst_34_n13}), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, new_AGEMA_signal_2941, sbox_inst_34_n12}), .c ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, new_AGEMA_signal_3529, sbox_inst_34_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_U7 ( .a ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, new_AGEMA_signal_2335, sbox_inst_34_T6}), .b ({input0_s3[139], input0_s2[139], input0_s1[139], input0_s0[139]}), .c ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, new_AGEMA_signal_2941, sbox_inst_34_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_t5_AND_U1 ( .a ({input0_s3[137], input0_s2[137], input0_s1[137], input0_s0[137]}), .b ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, new_AGEMA_signal_1273, sbox_inst_34_T3}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, new_AGEMA_signal_2332, sbox_inst_34_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_34_t6_AND_U1 ( .a ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, new_AGEMA_signal_1255, sbox_inst_34_L0}), .b ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, new_AGEMA_signal_1267, sbox_inst_34_T1}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, new_AGEMA_signal_2335, sbox_inst_34_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U15 ( .a ({new_AGEMA_signal_1302, new_AGEMA_signal_1301, new_AGEMA_signal_1300, sbox_inst_33_T2}), .b ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, sbox_inst_33_n20}), .c ({output0_s3[73], output0_s2[73], output0_s1[73], output0_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U14 ( .a ({new_AGEMA_signal_2952, new_AGEMA_signal_2951, new_AGEMA_signal_2950, sbox_inst_33_n19}), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, new_AGEMA_signal_2947, sbox_inst_33_n18}), .c ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, sbox_inst_33_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U13 ( .a ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, new_AGEMA_signal_1297, sbox_inst_33_T1}), .b ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, new_AGEMA_signal_2347, sbox_inst_33_T5}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, new_AGEMA_signal_2947, sbox_inst_33_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U11 ( .a ({input0_s3[133], input0_s2[133], input0_s1[133], input0_s0[133]}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, new_AGEMA_signal_2953, sbox_inst_33_n16}), .c ({output0_s3[113], output0_s2[113], output0_s1[113], output0_s0[113]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U10 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, sbox_inst_33_n15}), .b ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, new_AGEMA_signal_2347, sbox_inst_33_T5}), .c ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, new_AGEMA_signal_2953, sbox_inst_33_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U9 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, sbox_inst_33_n15}), .b ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, new_AGEMA_signal_3541, sbox_inst_33_n14}), .c ({output0_s3[153], output0_s2[153], output0_s1[153], output0_s0[153]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U8 ( .a ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, new_AGEMA_signal_2338, sbox_inst_33_n13}), .b ({new_AGEMA_signal_2958, new_AGEMA_signal_2957, new_AGEMA_signal_2956, sbox_inst_33_n12}), .c ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, new_AGEMA_signal_3541, sbox_inst_33_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_U7 ( .a ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, sbox_inst_33_T6}), .b ({input0_s3[135], input0_s2[135], input0_s1[135], input0_s0[135]}), .c ({new_AGEMA_signal_2958, new_AGEMA_signal_2957, new_AGEMA_signal_2956, sbox_inst_33_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_t5_AND_U1 ( .a ({input0_s3[133], input0_s2[133], input0_s1[133], input0_s0[133]}), .b ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, new_AGEMA_signal_1303, sbox_inst_33_T3}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, new_AGEMA_signal_2347, sbox_inst_33_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_33_t6_AND_U1 ( .a ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, new_AGEMA_signal_1285, sbox_inst_33_L0}), .b ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, new_AGEMA_signal_1297, sbox_inst_33_T1}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, sbox_inst_33_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U15 ( .a ({new_AGEMA_signal_1332, new_AGEMA_signal_1331, new_AGEMA_signal_1330, sbox_inst_32_T2}), .b ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, new_AGEMA_signal_3547, sbox_inst_32_n20}), .c ({output0_s3[72], output0_s2[72], output0_s1[72], output0_s0[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U14 ( .a ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, new_AGEMA_signal_2965, sbox_inst_32_n19}), .b ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, new_AGEMA_signal_2962, sbox_inst_32_n18}), .c ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, new_AGEMA_signal_3547, sbox_inst_32_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U13 ( .a ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, sbox_inst_32_T1}), .b ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, sbox_inst_32_T5}), .c ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, new_AGEMA_signal_2962, sbox_inst_32_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U11 ( .a ({input0_s3[129], input0_s2[129], input0_s1[129], input0_s0[129]}), .b ({new_AGEMA_signal_2970, new_AGEMA_signal_2969, new_AGEMA_signal_2968, sbox_inst_32_n16}), .c ({output0_s3[112], output0_s2[112], output0_s1[112], output0_s0[112]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U10 ( .a ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, new_AGEMA_signal_2356, sbox_inst_32_n15}), .b ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, sbox_inst_32_T5}), .c ({new_AGEMA_signal_2970, new_AGEMA_signal_2969, new_AGEMA_signal_2968, sbox_inst_32_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U9 ( .a ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, new_AGEMA_signal_2356, sbox_inst_32_n15}), .b ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, new_AGEMA_signal_3553, sbox_inst_32_n14}), .c ({output0_s3[152], output0_s2[152], output0_s1[152], output0_s0[152]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U8 ( .a ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, sbox_inst_32_n13}), .b ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, new_AGEMA_signal_2971, sbox_inst_32_n12}), .c ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, new_AGEMA_signal_3553, sbox_inst_32_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_U7 ( .a ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, new_AGEMA_signal_2365, sbox_inst_32_T6}), .b ({input0_s3[131], input0_s2[131], input0_s1[131], input0_s0[131]}), .c ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, new_AGEMA_signal_2971, sbox_inst_32_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_t5_AND_U1 ( .a ({input0_s3[129], input0_s2[129], input0_s1[129], input0_s0[129]}), .b ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, new_AGEMA_signal_1333, sbox_inst_32_T3}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, sbox_inst_32_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_32_t6_AND_U1 ( .a ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, new_AGEMA_signal_1315, sbox_inst_32_L0}), .b ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, new_AGEMA_signal_1327, sbox_inst_32_T1}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, new_AGEMA_signal_2365, sbox_inst_32_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U15 ( .a ({new_AGEMA_signal_1362, new_AGEMA_signal_1361, new_AGEMA_signal_1360, sbox_inst_31_T2}), .b ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, sbox_inst_31_n20}), .c ({output0_s3[71], output0_s2[71], output0_s1[71], output0_s0[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U14 ( .a ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, new_AGEMA_signal_2980, sbox_inst_31_n19}), .b ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, new_AGEMA_signal_2977, sbox_inst_31_n18}), .c ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, sbox_inst_31_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U13 ( .a ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, new_AGEMA_signal_1357, sbox_inst_31_T1}), .b ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, sbox_inst_31_T5}), .c ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, new_AGEMA_signal_2977, sbox_inst_31_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U11 ( .a ({input0_s3[125], input0_s2[125], input0_s1[125], input0_s0[125]}), .b ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, new_AGEMA_signal_2983, sbox_inst_31_n16}), .c ({output0_s3[111], output0_s2[111], output0_s1[111], output0_s0[111]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U10 ( .a ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, sbox_inst_31_n15}), .b ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, sbox_inst_31_T5}), .c ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, new_AGEMA_signal_2983, sbox_inst_31_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U9 ( .a ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, sbox_inst_31_n15}), .b ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, new_AGEMA_signal_3565, sbox_inst_31_n14}), .c ({output0_s3[151], output0_s2[151], output0_s1[151], output0_s0[151]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U8 ( .a ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, new_AGEMA_signal_2368, sbox_inst_31_n13}), .b ({new_AGEMA_signal_2988, new_AGEMA_signal_2987, new_AGEMA_signal_2986, sbox_inst_31_n12}), .c ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, new_AGEMA_signal_3565, sbox_inst_31_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_U7 ( .a ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, new_AGEMA_signal_2380, sbox_inst_31_T6}), .b ({input0_s3[127], input0_s2[127], input0_s1[127], input0_s0[127]}), .c ({new_AGEMA_signal_2988, new_AGEMA_signal_2987, new_AGEMA_signal_2986, sbox_inst_31_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_t5_AND_U1 ( .a ({input0_s3[125], input0_s2[125], input0_s1[125], input0_s0[125]}), .b ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, new_AGEMA_signal_1363, sbox_inst_31_T3}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, sbox_inst_31_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_31_t6_AND_U1 ( .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, new_AGEMA_signal_1345, sbox_inst_31_L0}), .b ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, new_AGEMA_signal_1357, sbox_inst_31_T1}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, new_AGEMA_signal_2380, sbox_inst_31_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U15 ( .a ({new_AGEMA_signal_1392, new_AGEMA_signal_1391, new_AGEMA_signal_1390, sbox_inst_30_T2}), .b ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, new_AGEMA_signal_3571, sbox_inst_30_n20}), .c ({output0_s3[70], output0_s2[70], output0_s1[70], output0_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U14 ( .a ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, new_AGEMA_signal_2995, sbox_inst_30_n19}), .b ({new_AGEMA_signal_2994, new_AGEMA_signal_2993, new_AGEMA_signal_2992, sbox_inst_30_n18}), .c ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, new_AGEMA_signal_3571, sbox_inst_30_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U13 ( .a ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, sbox_inst_30_T1}), .b ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, new_AGEMA_signal_2392, sbox_inst_30_T5}), .c ({new_AGEMA_signal_2994, new_AGEMA_signal_2993, new_AGEMA_signal_2992, sbox_inst_30_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U11 ( .a ({input0_s3[121], input0_s2[121], input0_s1[121], input0_s0[121]}), .b ({new_AGEMA_signal_3000, new_AGEMA_signal_2999, new_AGEMA_signal_2998, sbox_inst_30_n16}), .c ({output0_s3[110], output0_s2[110], output0_s1[110], output0_s0[110]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U10 ( .a ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, sbox_inst_30_n15}), .b ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, new_AGEMA_signal_2392, sbox_inst_30_T5}), .c ({new_AGEMA_signal_3000, new_AGEMA_signal_2999, new_AGEMA_signal_2998, sbox_inst_30_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U9 ( .a ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, sbox_inst_30_n15}), .b ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, new_AGEMA_signal_3577, sbox_inst_30_n14}), .c ({output0_s3[150], output0_s2[150], output0_s1[150], output0_s0[150]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U8 ( .a ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, new_AGEMA_signal_2383, sbox_inst_30_n13}), .b ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, new_AGEMA_signal_3001, sbox_inst_30_n12}), .c ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, new_AGEMA_signal_3577, sbox_inst_30_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_U7 ( .a ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, new_AGEMA_signal_2395, sbox_inst_30_T6}), .b ({input0_s3[123], input0_s2[123], input0_s1[123], input0_s0[123]}), .c ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, new_AGEMA_signal_3001, sbox_inst_30_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_t5_AND_U1 ( .a ({input0_s3[121], input0_s2[121], input0_s1[121], input0_s0[121]}), .b ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, new_AGEMA_signal_1393, sbox_inst_30_T3}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, new_AGEMA_signal_2392, sbox_inst_30_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_30_t6_AND_U1 ( .a ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, new_AGEMA_signal_1375, sbox_inst_30_L0}), .b ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, new_AGEMA_signal_1387, sbox_inst_30_T1}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, new_AGEMA_signal_2395, sbox_inst_30_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U15 ( .a ({new_AGEMA_signal_1422, new_AGEMA_signal_1421, new_AGEMA_signal_1420, sbox_inst_29_T2}), .b ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, sbox_inst_29_n20}), .c ({output0_s3[69], output0_s2[69], output0_s1[69], output0_s0[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U14 ( .a ({new_AGEMA_signal_3012, new_AGEMA_signal_3011, new_AGEMA_signal_3010, sbox_inst_29_n19}), .b ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, new_AGEMA_signal_3007, sbox_inst_29_n18}), .c ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, sbox_inst_29_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U13 ( .a ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, new_AGEMA_signal_1417, sbox_inst_29_T1}), .b ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, sbox_inst_29_T5}), .c ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, new_AGEMA_signal_3007, sbox_inst_29_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U11 ( .a ({input0_s3[117], input0_s2[117], input0_s1[117], input0_s0[117]}), .b ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, new_AGEMA_signal_3013, sbox_inst_29_n16}), .c ({output0_s3[109], output0_s2[109], output0_s1[109], output0_s0[109]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U10 ( .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, sbox_inst_29_n15}), .b ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, sbox_inst_29_T5}), .c ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, new_AGEMA_signal_3013, sbox_inst_29_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U9 ( .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_2401, sbox_inst_29_n15}), .b ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, new_AGEMA_signal_3589, sbox_inst_29_n14}), .c ({output0_s3[149], output0_s2[149], output0_s1[149], output0_s0[149]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U8 ( .a ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, sbox_inst_29_n13}), .b ({new_AGEMA_signal_3018, new_AGEMA_signal_3017, new_AGEMA_signal_3016, sbox_inst_29_n12}), .c ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, new_AGEMA_signal_3589, sbox_inst_29_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_U7 ( .a ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, sbox_inst_29_T6}), .b ({input0_s3[119], input0_s2[119], input0_s1[119], input0_s0[119]}), .c ({new_AGEMA_signal_3018, new_AGEMA_signal_3017, new_AGEMA_signal_3016, sbox_inst_29_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_t5_AND_U1 ( .a ({input0_s3[117], input0_s2[117], input0_s1[117], input0_s0[117]}), .b ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, new_AGEMA_signal_1423, sbox_inst_29_T3}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, sbox_inst_29_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_29_t6_AND_U1 ( .a ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, new_AGEMA_signal_1405, sbox_inst_29_L0}), .b ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, new_AGEMA_signal_1417, sbox_inst_29_T1}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, new_AGEMA_signal_2410, sbox_inst_29_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U15 ( .a ({new_AGEMA_signal_1452, new_AGEMA_signal_1451, new_AGEMA_signal_1450, sbox_inst_28_T2}), .b ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, new_AGEMA_signal_3595, sbox_inst_28_n20}), .c ({output0_s3[68], output0_s2[68], output0_s1[68], output0_s0[68]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U14 ( .a ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, new_AGEMA_signal_3025, sbox_inst_28_n19}), .b ({new_AGEMA_signal_3024, new_AGEMA_signal_3023, new_AGEMA_signal_3022, sbox_inst_28_n18}), .c ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, new_AGEMA_signal_3595, sbox_inst_28_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U13 ( .a ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, sbox_inst_28_T1}), .b ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, sbox_inst_28_T5}), .c ({new_AGEMA_signal_3024, new_AGEMA_signal_3023, new_AGEMA_signal_3022, sbox_inst_28_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U11 ( .a ({input0_s3[113], input0_s2[113], input0_s1[113], input0_s0[113]}), .b ({new_AGEMA_signal_3030, new_AGEMA_signal_3029, new_AGEMA_signal_3028, sbox_inst_28_n16}), .c ({output0_s3[108], output0_s2[108], output0_s1[108], output0_s0[108]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U10 ( .a ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, sbox_inst_28_n15}), .b ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, sbox_inst_28_T5}), .c ({new_AGEMA_signal_3030, new_AGEMA_signal_3029, new_AGEMA_signal_3028, sbox_inst_28_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U9 ( .a ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, sbox_inst_28_n15}), .b ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, new_AGEMA_signal_3601, sbox_inst_28_n14}), .c ({output0_s3[148], output0_s2[148], output0_s1[148], output0_s0[148]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U8 ( .a ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2413, sbox_inst_28_n13}), .b ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, new_AGEMA_signal_3031, sbox_inst_28_n12}), .c ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, new_AGEMA_signal_3601, sbox_inst_28_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_U7 ( .a ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, sbox_inst_28_T6}), .b ({input0_s3[115], input0_s2[115], input0_s1[115], input0_s0[115]}), .c ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, new_AGEMA_signal_3031, sbox_inst_28_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_t5_AND_U1 ( .a ({input0_s3[113], input0_s2[113], input0_s1[113], input0_s0[113]}), .b ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, new_AGEMA_signal_1453, sbox_inst_28_T3}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, sbox_inst_28_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_28_t6_AND_U1 ( .a ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, new_AGEMA_signal_1435, sbox_inst_28_L0}), .b ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, new_AGEMA_signal_1447, sbox_inst_28_T1}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, sbox_inst_28_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U15 ( .a ({new_AGEMA_signal_1482, new_AGEMA_signal_1481, new_AGEMA_signal_1480, sbox_inst_27_T2}), .b ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, new_AGEMA_signal_3607, sbox_inst_27_n20}), .c ({output0_s3[67], output0_s2[67], output0_s1[67], output0_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U14 ( .a ({new_AGEMA_signal_3042, new_AGEMA_signal_3041, new_AGEMA_signal_3040, sbox_inst_27_n19}), .b ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, new_AGEMA_signal_3037, sbox_inst_27_n18}), .c ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, new_AGEMA_signal_3607, sbox_inst_27_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U13 ( .a ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, new_AGEMA_signal_1477, sbox_inst_27_T1}), .b ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, new_AGEMA_signal_2437, sbox_inst_27_T5}), .c ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, new_AGEMA_signal_3037, sbox_inst_27_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U11 ( .a ({input0_s3[109], input0_s2[109], input0_s1[109], input0_s0[109]}), .b ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, new_AGEMA_signal_3043, sbox_inst_27_n16}), .c ({output0_s3[107], output0_s2[107], output0_s1[107], output0_s0[107]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U10 ( .a ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, sbox_inst_27_n15}), .b ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, new_AGEMA_signal_2437, sbox_inst_27_T5}), .c ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, new_AGEMA_signal_3043, sbox_inst_27_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U9 ( .a ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, sbox_inst_27_n15}), .b ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, new_AGEMA_signal_3613, sbox_inst_27_n14}), .c ({output0_s3[147], output0_s2[147], output0_s1[147], output0_s0[147]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U8 ( .a ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, new_AGEMA_signal_2428, sbox_inst_27_n13}), .b ({new_AGEMA_signal_3048, new_AGEMA_signal_3047, new_AGEMA_signal_3046, sbox_inst_27_n12}), .c ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, new_AGEMA_signal_3613, sbox_inst_27_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_U7 ( .a ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, sbox_inst_27_T6}), .b ({input0_s3[111], input0_s2[111], input0_s1[111], input0_s0[111]}), .c ({new_AGEMA_signal_3048, new_AGEMA_signal_3047, new_AGEMA_signal_3046, sbox_inst_27_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_t5_AND_U1 ( .a ({input0_s3[109], input0_s2[109], input0_s1[109], input0_s0[109]}), .b ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, new_AGEMA_signal_1483, sbox_inst_27_T3}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, new_AGEMA_signal_2437, sbox_inst_27_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_27_t6_AND_U1 ( .a ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, new_AGEMA_signal_1465, sbox_inst_27_L0}), .b ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, new_AGEMA_signal_1477, sbox_inst_27_T1}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, sbox_inst_27_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U15 ( .a ({new_AGEMA_signal_1512, new_AGEMA_signal_1511, new_AGEMA_signal_1510, sbox_inst_26_T2}), .b ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, new_AGEMA_signal_3619, sbox_inst_26_n20}), .c ({output0_s3[66], output0_s2[66], output0_s1[66], output0_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U14 ( .a ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, new_AGEMA_signal_3055, sbox_inst_26_n19}), .b ({new_AGEMA_signal_3054, new_AGEMA_signal_3053, new_AGEMA_signal_3052, sbox_inst_26_n18}), .c ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, new_AGEMA_signal_3619, sbox_inst_26_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U13 ( .a ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, sbox_inst_26_T1}), .b ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, sbox_inst_26_T5}), .c ({new_AGEMA_signal_3054, new_AGEMA_signal_3053, new_AGEMA_signal_3052, sbox_inst_26_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U11 ( .a ({input0_s3[105], input0_s2[105], input0_s1[105], input0_s0[105]}), .b ({new_AGEMA_signal_3060, new_AGEMA_signal_3059, new_AGEMA_signal_3058, sbox_inst_26_n16}), .c ({output0_s3[106], output0_s2[106], output0_s1[106], output0_s0[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U10 ( .a ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, sbox_inst_26_n15}), .b ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, sbox_inst_26_T5}), .c ({new_AGEMA_signal_3060, new_AGEMA_signal_3059, new_AGEMA_signal_3058, sbox_inst_26_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U9 ( .a ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, new_AGEMA_signal_2446, sbox_inst_26_n15}), .b ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, new_AGEMA_signal_3625, sbox_inst_26_n14}), .c ({output0_s3[146], output0_s2[146], output0_s1[146], output0_s0[146]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U8 ( .a ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, new_AGEMA_signal_2443, sbox_inst_26_n13}), .b ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, new_AGEMA_signal_3061, sbox_inst_26_n12}), .c ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, new_AGEMA_signal_3625, sbox_inst_26_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_U7 ( .a ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, new_AGEMA_signal_2455, sbox_inst_26_T6}), .b ({input0_s3[107], input0_s2[107], input0_s1[107], input0_s0[107]}), .c ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, new_AGEMA_signal_3061, sbox_inst_26_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_t5_AND_U1 ( .a ({input0_s3[105], input0_s2[105], input0_s1[105], input0_s0[105]}), .b ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, new_AGEMA_signal_1513, sbox_inst_26_T3}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, sbox_inst_26_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_26_t6_AND_U1 ( .a ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, new_AGEMA_signal_1495, sbox_inst_26_L0}), .b ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, new_AGEMA_signal_1507, sbox_inst_26_T1}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, new_AGEMA_signal_2455, sbox_inst_26_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U15 ( .a ({new_AGEMA_signal_1542, new_AGEMA_signal_1541, new_AGEMA_signal_1540, sbox_inst_25_T2}), .b ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, new_AGEMA_signal_3631, sbox_inst_25_n20}), .c ({output0_s3[65], output0_s2[65], output0_s1[65], output0_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U14 ( .a ({new_AGEMA_signal_3072, new_AGEMA_signal_3071, new_AGEMA_signal_3070, sbox_inst_25_n19}), .b ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, new_AGEMA_signal_3067, sbox_inst_25_n18}), .c ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, new_AGEMA_signal_3631, sbox_inst_25_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U13 ( .a ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, new_AGEMA_signal_1537, sbox_inst_25_T1}), .b ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, sbox_inst_25_T5}), .c ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, new_AGEMA_signal_3067, sbox_inst_25_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U11 ( .a ({input0_s3[101], input0_s2[101], input0_s1[101], input0_s0[101]}), .b ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, new_AGEMA_signal_3073, sbox_inst_25_n16}), .c ({output0_s3[105], output0_s2[105], output0_s1[105], output0_s0[105]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U10 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, new_AGEMA_signal_2461, sbox_inst_25_n15}), .b ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, sbox_inst_25_T5}), .c ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, new_AGEMA_signal_3073, sbox_inst_25_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U9 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, new_AGEMA_signal_2461, sbox_inst_25_n15}), .b ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, new_AGEMA_signal_3637, sbox_inst_25_n14}), .c ({output0_s3[145], output0_s2[145], output0_s1[145], output0_s0[145]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U8 ( .a ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, sbox_inst_25_n13}), .b ({new_AGEMA_signal_3078, new_AGEMA_signal_3077, new_AGEMA_signal_3076, sbox_inst_25_n12}), .c ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, new_AGEMA_signal_3637, sbox_inst_25_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_U7 ( .a ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, sbox_inst_25_T6}), .b ({input0_s3[103], input0_s2[103], input0_s1[103], input0_s0[103]}), .c ({new_AGEMA_signal_3078, new_AGEMA_signal_3077, new_AGEMA_signal_3076, sbox_inst_25_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_t5_AND_U1 ( .a ({input0_s3[101], input0_s2[101], input0_s1[101], input0_s0[101]}), .b ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, new_AGEMA_signal_1543, sbox_inst_25_T3}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, sbox_inst_25_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_25_t6_AND_U1 ( .a ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, new_AGEMA_signal_1525, sbox_inst_25_L0}), .b ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, new_AGEMA_signal_1537, sbox_inst_25_T1}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, sbox_inst_25_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U15 ( .a ({new_AGEMA_signal_1572, new_AGEMA_signal_1571, new_AGEMA_signal_1570, sbox_inst_24_T2}), .b ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, new_AGEMA_signal_3643, sbox_inst_24_n20}), .c ({output0_s3[64], output0_s2[64], output0_s1[64], output0_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U14 ( .a ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, new_AGEMA_signal_3085, sbox_inst_24_n19}), .b ({new_AGEMA_signal_3084, new_AGEMA_signal_3083, new_AGEMA_signal_3082, sbox_inst_24_n18}), .c ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, new_AGEMA_signal_3643, sbox_inst_24_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U13 ( .a ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, new_AGEMA_signal_1567, sbox_inst_24_T1}), .b ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, sbox_inst_24_T5}), .c ({new_AGEMA_signal_3084, new_AGEMA_signal_3083, new_AGEMA_signal_3082, sbox_inst_24_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U11 ( .a ({input0_s3[97], input0_s2[97], input0_s1[97], input0_s0[97]}), .b ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, new_AGEMA_signal_3088, sbox_inst_24_n16}), .c ({output0_s3[104], output0_s2[104], output0_s1[104], output0_s0[104]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U10 ( .a ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, new_AGEMA_signal_2476, sbox_inst_24_n15}), .b ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, sbox_inst_24_T5}), .c ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, new_AGEMA_signal_3088, sbox_inst_24_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U9 ( .a ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, new_AGEMA_signal_2476, sbox_inst_24_n15}), .b ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, new_AGEMA_signal_3649, sbox_inst_24_n14}), .c ({output0_s3[144], output0_s2[144], output0_s1[144], output0_s0[144]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U8 ( .a ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, new_AGEMA_signal_2473, sbox_inst_24_n13}), .b ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, new_AGEMA_signal_3091, sbox_inst_24_n12}), .c ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, new_AGEMA_signal_3649, sbox_inst_24_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_U7 ( .a ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, new_AGEMA_signal_2485, sbox_inst_24_T6}), .b ({input0_s3[99], input0_s2[99], input0_s1[99], input0_s0[99]}), .c ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, new_AGEMA_signal_3091, sbox_inst_24_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_t5_AND_U1 ( .a ({input0_s3[97], input0_s2[97], input0_s1[97], input0_s0[97]}), .b ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, new_AGEMA_signal_1573, sbox_inst_24_T3}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, new_AGEMA_signal_2482, sbox_inst_24_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_24_t6_AND_U1 ( .a ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, new_AGEMA_signal_1555, sbox_inst_24_L0}), .b ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, new_AGEMA_signal_1567, sbox_inst_24_T1}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, new_AGEMA_signal_2485, sbox_inst_24_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U15 ( .a ({new_AGEMA_signal_1602, new_AGEMA_signal_1601, new_AGEMA_signal_1600, sbox_inst_23_T2}), .b ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, new_AGEMA_signal_3655, sbox_inst_23_n20}), .c ({output0_s3[63], output0_s2[63], output0_s1[63], output0_s0[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U14 ( .a ({new_AGEMA_signal_3102, new_AGEMA_signal_3101, new_AGEMA_signal_3100, sbox_inst_23_n19}), .b ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, new_AGEMA_signal_3097, sbox_inst_23_n18}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, new_AGEMA_signal_3655, sbox_inst_23_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U13 ( .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, sbox_inst_23_T1}), .b ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, new_AGEMA_signal_2497, sbox_inst_23_T5}), .c ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, new_AGEMA_signal_3097, sbox_inst_23_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U11 ( .a ({input0_s3[93], input0_s2[93], input0_s1[93], input0_s0[93]}), .b ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, new_AGEMA_signal_3103, sbox_inst_23_n16}), .c ({output0_s3[103], output0_s2[103], output0_s1[103], output0_s0[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U10 ( .a ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, new_AGEMA_signal_2491, sbox_inst_23_n15}), .b ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, new_AGEMA_signal_2497, sbox_inst_23_T5}), .c ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, new_AGEMA_signal_3103, sbox_inst_23_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U9 ( .a ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, new_AGEMA_signal_2491, sbox_inst_23_n15}), .b ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, new_AGEMA_signal_3661, sbox_inst_23_n14}), .c ({output0_s3[143], output0_s2[143], output0_s1[143], output0_s0[143]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U8 ( .a ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, new_AGEMA_signal_2488, sbox_inst_23_n13}), .b ({new_AGEMA_signal_3108, new_AGEMA_signal_3107, new_AGEMA_signal_3106, sbox_inst_23_n12}), .c ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, new_AGEMA_signal_3661, sbox_inst_23_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_U7 ( .a ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, new_AGEMA_signal_2500, sbox_inst_23_T6}), .b ({input0_s3[95], input0_s2[95], input0_s1[95], input0_s0[95]}), .c ({new_AGEMA_signal_3108, new_AGEMA_signal_3107, new_AGEMA_signal_3106, sbox_inst_23_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_t5_AND_U1 ( .a ({input0_s3[93], input0_s2[93], input0_s1[93], input0_s0[93]}), .b ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, new_AGEMA_signal_1603, sbox_inst_23_T3}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, new_AGEMA_signal_2497, sbox_inst_23_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_23_t6_AND_U1 ( .a ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, new_AGEMA_signal_1585, sbox_inst_23_L0}), .b ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, new_AGEMA_signal_1597, sbox_inst_23_T1}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, new_AGEMA_signal_2500, sbox_inst_23_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U15 ( .a ({new_AGEMA_signal_1632, new_AGEMA_signal_1631, new_AGEMA_signal_1630, sbox_inst_22_T2}), .b ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, new_AGEMA_signal_3667, sbox_inst_22_n20}), .c ({output0_s3[62], output0_s2[62], output0_s1[62], output0_s0[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U14 ( .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, new_AGEMA_signal_3115, sbox_inst_22_n19}), .b ({new_AGEMA_signal_3114, new_AGEMA_signal_3113, new_AGEMA_signal_3112, sbox_inst_22_n18}), .c ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, new_AGEMA_signal_3667, sbox_inst_22_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U13 ( .a ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, new_AGEMA_signal_1627, sbox_inst_22_T1}), .b ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, new_AGEMA_signal_2512, sbox_inst_22_T5}), .c ({new_AGEMA_signal_3114, new_AGEMA_signal_3113, new_AGEMA_signal_3112, sbox_inst_22_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U11 ( .a ({input0_s3[89], input0_s2[89], input0_s1[89], input0_s0[89]}), .b ({new_AGEMA_signal_3120, new_AGEMA_signal_3119, new_AGEMA_signal_3118, sbox_inst_22_n16}), .c ({output0_s3[102], output0_s2[102], output0_s1[102], output0_s0[102]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U10 ( .a ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, new_AGEMA_signal_2506, sbox_inst_22_n15}), .b ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, new_AGEMA_signal_2512, sbox_inst_22_T5}), .c ({new_AGEMA_signal_3120, new_AGEMA_signal_3119, new_AGEMA_signal_3118, sbox_inst_22_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U9 ( .a ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, new_AGEMA_signal_2506, sbox_inst_22_n15}), .b ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, new_AGEMA_signal_3673, sbox_inst_22_n14}), .c ({output0_s3[142], output0_s2[142], output0_s1[142], output0_s0[142]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U8 ( .a ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, new_AGEMA_signal_2503, sbox_inst_22_n13}), .b ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, new_AGEMA_signal_3121, sbox_inst_22_n12}), .c ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, new_AGEMA_signal_3673, sbox_inst_22_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_U7 ( .a ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, new_AGEMA_signal_2515, sbox_inst_22_T6}), .b ({input0_s3[91], input0_s2[91], input0_s1[91], input0_s0[91]}), .c ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, new_AGEMA_signal_3121, sbox_inst_22_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_t5_AND_U1 ( .a ({input0_s3[89], input0_s2[89], input0_s1[89], input0_s0[89]}), .b ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, new_AGEMA_signal_1633, sbox_inst_22_T3}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, new_AGEMA_signal_2512, sbox_inst_22_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_22_t6_AND_U1 ( .a ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, new_AGEMA_signal_1615, sbox_inst_22_L0}), .b ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, new_AGEMA_signal_1627, sbox_inst_22_T1}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, new_AGEMA_signal_2515, sbox_inst_22_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U15 ( .a ({new_AGEMA_signal_1662, new_AGEMA_signal_1661, new_AGEMA_signal_1660, sbox_inst_21_T2}), .b ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, new_AGEMA_signal_3679, sbox_inst_21_n20}), .c ({output0_s3[61], output0_s2[61], output0_s1[61], output0_s0[61]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U14 ( .a ({new_AGEMA_signal_3132, new_AGEMA_signal_3131, new_AGEMA_signal_3130, sbox_inst_21_n19}), .b ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, new_AGEMA_signal_3127, sbox_inst_21_n18}), .c ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, new_AGEMA_signal_3679, sbox_inst_21_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U13 ( .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, new_AGEMA_signal_1657, sbox_inst_21_T1}), .b ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, new_AGEMA_signal_2527, sbox_inst_21_T5}), .c ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, new_AGEMA_signal_3127, sbox_inst_21_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U11 ( .a ({input0_s3[85], input0_s2[85], input0_s1[85], input0_s0[85]}), .b ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, new_AGEMA_signal_3133, sbox_inst_21_n16}), .c ({output0_s3[101], output0_s2[101], output0_s1[101], output0_s0[101]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U10 ( .a ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, new_AGEMA_signal_2521, sbox_inst_21_n15}), .b ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, new_AGEMA_signal_2527, sbox_inst_21_T5}), .c ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, new_AGEMA_signal_3133, sbox_inst_21_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U9 ( .a ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, new_AGEMA_signal_2521, sbox_inst_21_n15}), .b ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, new_AGEMA_signal_3685, sbox_inst_21_n14}), .c ({output0_s3[141], output0_s2[141], output0_s1[141], output0_s0[141]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U8 ( .a ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, new_AGEMA_signal_2518, sbox_inst_21_n13}), .b ({new_AGEMA_signal_3138, new_AGEMA_signal_3137, new_AGEMA_signal_3136, sbox_inst_21_n12}), .c ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, new_AGEMA_signal_3685, sbox_inst_21_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_U7 ( .a ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, new_AGEMA_signal_2530, sbox_inst_21_T6}), .b ({input0_s3[87], input0_s2[87], input0_s1[87], input0_s0[87]}), .c ({new_AGEMA_signal_3138, new_AGEMA_signal_3137, new_AGEMA_signal_3136, sbox_inst_21_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_t5_AND_U1 ( .a ({input0_s3[85], input0_s2[85], input0_s1[85], input0_s0[85]}), .b ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, new_AGEMA_signal_1663, sbox_inst_21_T3}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, new_AGEMA_signal_2527, sbox_inst_21_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_21_t6_AND_U1 ( .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, new_AGEMA_signal_1645, sbox_inst_21_L0}), .b ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, new_AGEMA_signal_1657, sbox_inst_21_T1}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, new_AGEMA_signal_2530, sbox_inst_21_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U15 ( .a ({new_AGEMA_signal_1692, new_AGEMA_signal_1691, new_AGEMA_signal_1690, sbox_inst_20_T2}), .b ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, new_AGEMA_signal_3691, sbox_inst_20_n20}), .c ({output0_s3[60], output0_s2[60], output0_s1[60], output0_s0[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U14 ( .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, new_AGEMA_signal_3145, sbox_inst_20_n19}), .b ({new_AGEMA_signal_3144, new_AGEMA_signal_3143, new_AGEMA_signal_3142, sbox_inst_20_n18}), .c ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, new_AGEMA_signal_3691, sbox_inst_20_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U13 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, sbox_inst_20_T1}), .b ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, sbox_inst_20_T5}), .c ({new_AGEMA_signal_3144, new_AGEMA_signal_3143, new_AGEMA_signal_3142, sbox_inst_20_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U11 ( .a ({input0_s3[81], input0_s2[81], input0_s1[81], input0_s0[81]}), .b ({new_AGEMA_signal_3150, new_AGEMA_signal_3149, new_AGEMA_signal_3148, sbox_inst_20_n16}), .c ({output0_s3[100], output0_s2[100], output0_s1[100], output0_s0[100]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U10 ( .a ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, new_AGEMA_signal_2536, sbox_inst_20_n15}), .b ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, sbox_inst_20_T5}), .c ({new_AGEMA_signal_3150, new_AGEMA_signal_3149, new_AGEMA_signal_3148, sbox_inst_20_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U9 ( .a ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, new_AGEMA_signal_2536, sbox_inst_20_n15}), .b ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, new_AGEMA_signal_3697, sbox_inst_20_n14}), .c ({output0_s3[140], output0_s2[140], output0_s1[140], output0_s0[140]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U8 ( .a ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, new_AGEMA_signal_2533, sbox_inst_20_n13}), .b ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, new_AGEMA_signal_3151, sbox_inst_20_n12}), .c ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, new_AGEMA_signal_3697, sbox_inst_20_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_U7 ( .a ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, new_AGEMA_signal_2545, sbox_inst_20_T6}), .b ({input0_s3[83], input0_s2[83], input0_s1[83], input0_s0[83]}), .c ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, new_AGEMA_signal_3151, sbox_inst_20_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_t5_AND_U1 ( .a ({input0_s3[81], input0_s2[81], input0_s1[81], input0_s0[81]}), .b ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, new_AGEMA_signal_1693, sbox_inst_20_T3}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, sbox_inst_20_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_20_t6_AND_U1 ( .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, new_AGEMA_signal_1675, sbox_inst_20_L0}), .b ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, new_AGEMA_signal_1687, sbox_inst_20_T1}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, new_AGEMA_signal_2545, sbox_inst_20_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U15 ( .a ({new_AGEMA_signal_1722, new_AGEMA_signal_1721, new_AGEMA_signal_1720, sbox_inst_19_T2}), .b ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, new_AGEMA_signal_3703, sbox_inst_19_n20}), .c ({output0_s3[59], output0_s2[59], output0_s1[59], output0_s0[59]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U14 ( .a ({new_AGEMA_signal_3162, new_AGEMA_signal_3161, new_AGEMA_signal_3160, sbox_inst_19_n19}), .b ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, new_AGEMA_signal_3157, sbox_inst_19_n18}), .c ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, new_AGEMA_signal_3703, sbox_inst_19_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U13 ( .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, new_AGEMA_signal_1717, sbox_inst_19_T1}), .b ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, new_AGEMA_signal_2557, sbox_inst_19_T5}), .c ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, new_AGEMA_signal_3157, sbox_inst_19_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U11 ( .a ({input0_s3[77], input0_s2[77], input0_s1[77], input0_s0[77]}), .b ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, new_AGEMA_signal_3163, sbox_inst_19_n16}), .c ({output0_s3[99], output0_s2[99], output0_s1[99], output0_s0[99]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U10 ( .a ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, new_AGEMA_signal_2551, sbox_inst_19_n15}), .b ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, new_AGEMA_signal_2557, sbox_inst_19_T5}), .c ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, new_AGEMA_signal_3163, sbox_inst_19_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U9 ( .a ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, new_AGEMA_signal_2551, sbox_inst_19_n15}), .b ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, new_AGEMA_signal_3709, sbox_inst_19_n14}), .c ({output0_s3[139], output0_s2[139], output0_s1[139], output0_s0[139]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U8 ( .a ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, new_AGEMA_signal_2548, sbox_inst_19_n13}), .b ({new_AGEMA_signal_3168, new_AGEMA_signal_3167, new_AGEMA_signal_3166, sbox_inst_19_n12}), .c ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, new_AGEMA_signal_3709, sbox_inst_19_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_U7 ( .a ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, new_AGEMA_signal_2560, sbox_inst_19_T6}), .b ({input0_s3[79], input0_s2[79], input0_s1[79], input0_s0[79]}), .c ({new_AGEMA_signal_3168, new_AGEMA_signal_3167, new_AGEMA_signal_3166, sbox_inst_19_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_t5_AND_U1 ( .a ({input0_s3[77], input0_s2[77], input0_s1[77], input0_s0[77]}), .b ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, new_AGEMA_signal_1723, sbox_inst_19_T3}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, new_AGEMA_signal_2557, sbox_inst_19_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_19_t6_AND_U1 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, new_AGEMA_signal_1705, sbox_inst_19_L0}), .b ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, new_AGEMA_signal_1717, sbox_inst_19_T1}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, new_AGEMA_signal_2560, sbox_inst_19_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U15 ( .a ({new_AGEMA_signal_1752, new_AGEMA_signal_1751, new_AGEMA_signal_1750, sbox_inst_18_T2}), .b ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, new_AGEMA_signal_3715, sbox_inst_18_n20}), .c ({output0_s3[58], output0_s2[58], output0_s1[58], output0_s0[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U14 ( .a ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, new_AGEMA_signal_3175, sbox_inst_18_n19}), .b ({new_AGEMA_signal_3174, new_AGEMA_signal_3173, new_AGEMA_signal_3172, sbox_inst_18_n18}), .c ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, new_AGEMA_signal_3715, sbox_inst_18_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U13 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, sbox_inst_18_T1}), .b ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, new_AGEMA_signal_2572, sbox_inst_18_T5}), .c ({new_AGEMA_signal_3174, new_AGEMA_signal_3173, new_AGEMA_signal_3172, sbox_inst_18_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U11 ( .a ({input0_s3[73], input0_s2[73], input0_s1[73], input0_s0[73]}), .b ({new_AGEMA_signal_3180, new_AGEMA_signal_3179, new_AGEMA_signal_3178, sbox_inst_18_n16}), .c ({output0_s3[98], output0_s2[98], output0_s1[98], output0_s0[98]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U10 ( .a ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, sbox_inst_18_n15}), .b ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, new_AGEMA_signal_2572, sbox_inst_18_T5}), .c ({new_AGEMA_signal_3180, new_AGEMA_signal_3179, new_AGEMA_signal_3178, sbox_inst_18_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U9 ( .a ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, sbox_inst_18_n15}), .b ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, new_AGEMA_signal_3721, sbox_inst_18_n14}), .c ({output0_s3[138], output0_s2[138], output0_s1[138], output0_s0[138]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U8 ( .a ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, new_AGEMA_signal_2563, sbox_inst_18_n13}), .b ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, new_AGEMA_signal_3181, sbox_inst_18_n12}), .c ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, new_AGEMA_signal_3721, sbox_inst_18_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_U7 ( .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, new_AGEMA_signal_2575, sbox_inst_18_T6}), .b ({input0_s3[75], input0_s2[75], input0_s1[75], input0_s0[75]}), .c ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, new_AGEMA_signal_3181, sbox_inst_18_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_t5_AND_U1 ( .a ({input0_s3[73], input0_s2[73], input0_s1[73], input0_s0[73]}), .b ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, new_AGEMA_signal_1753, sbox_inst_18_T3}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, new_AGEMA_signal_2572, sbox_inst_18_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_18_t6_AND_U1 ( .a ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, new_AGEMA_signal_1735, sbox_inst_18_L0}), .b ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, new_AGEMA_signal_1747, sbox_inst_18_T1}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, new_AGEMA_signal_2575, sbox_inst_18_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U15 ( .a ({new_AGEMA_signal_1782, new_AGEMA_signal_1781, new_AGEMA_signal_1780, sbox_inst_17_T2}), .b ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, new_AGEMA_signal_3727, sbox_inst_17_n20}), .c ({output0_s3[57], output0_s2[57], output0_s1[57], output0_s0[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U14 ( .a ({new_AGEMA_signal_3192, new_AGEMA_signal_3191, new_AGEMA_signal_3190, sbox_inst_17_n19}), .b ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, new_AGEMA_signal_3187, sbox_inst_17_n18}), .c ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, new_AGEMA_signal_3727, sbox_inst_17_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U13 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, sbox_inst_17_T1}), .b ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2587, sbox_inst_17_T5}), .c ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, new_AGEMA_signal_3187, sbox_inst_17_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U11 ( .a ({input0_s3[69], input0_s2[69], input0_s1[69], input0_s0[69]}), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, new_AGEMA_signal_3193, sbox_inst_17_n16}), .c ({output0_s3[97], output0_s2[97], output0_s1[97], output0_s0[97]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U10 ( .a ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, new_AGEMA_signal_2581, sbox_inst_17_n15}), .b ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2587, sbox_inst_17_T5}), .c ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, new_AGEMA_signal_3193, sbox_inst_17_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U9 ( .a ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, new_AGEMA_signal_2581, sbox_inst_17_n15}), .b ({new_AGEMA_signal_3735, new_AGEMA_signal_3734, new_AGEMA_signal_3733, sbox_inst_17_n14}), .c ({output0_s3[137], output0_s2[137], output0_s1[137], output0_s0[137]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U8 ( .a ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, sbox_inst_17_n13}), .b ({new_AGEMA_signal_3198, new_AGEMA_signal_3197, new_AGEMA_signal_3196, sbox_inst_17_n12}), .c ({new_AGEMA_signal_3735, new_AGEMA_signal_3734, new_AGEMA_signal_3733, sbox_inst_17_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_U7 ( .a ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, new_AGEMA_signal_2590, sbox_inst_17_T6}), .b ({input0_s3[71], input0_s2[71], input0_s1[71], input0_s0[71]}), .c ({new_AGEMA_signal_3198, new_AGEMA_signal_3197, new_AGEMA_signal_3196, sbox_inst_17_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_t5_AND_U1 ( .a ({input0_s3[69], input0_s2[69], input0_s1[69], input0_s0[69]}), .b ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, new_AGEMA_signal_1783, sbox_inst_17_T3}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2587, sbox_inst_17_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_17_t6_AND_U1 ( .a ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, new_AGEMA_signal_1765, sbox_inst_17_L0}), .b ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, new_AGEMA_signal_1777, sbox_inst_17_T1}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, new_AGEMA_signal_2590, sbox_inst_17_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U15 ( .a ({new_AGEMA_signal_1812, new_AGEMA_signal_1811, new_AGEMA_signal_1810, sbox_inst_16_T2}), .b ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, new_AGEMA_signal_3739, sbox_inst_16_n20}), .c ({output0_s3[56], output0_s2[56], output0_s1[56], output0_s0[56]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U14 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, new_AGEMA_signal_3205, sbox_inst_16_n19}), .b ({new_AGEMA_signal_3204, new_AGEMA_signal_3203, new_AGEMA_signal_3202, sbox_inst_16_n18}), .c ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, new_AGEMA_signal_3739, sbox_inst_16_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U13 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, new_AGEMA_signal_1807, sbox_inst_16_T1}), .b ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, new_AGEMA_signal_2602, sbox_inst_16_T5}), .c ({new_AGEMA_signal_3204, new_AGEMA_signal_3203, new_AGEMA_signal_3202, sbox_inst_16_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U11 ( .a ({input0_s3[65], input0_s2[65], input0_s1[65], input0_s0[65]}), .b ({new_AGEMA_signal_3210, new_AGEMA_signal_3209, new_AGEMA_signal_3208, sbox_inst_16_n16}), .c ({output0_s3[96], output0_s2[96], output0_s1[96], output0_s0[96]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U10 ( .a ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, new_AGEMA_signal_2596, sbox_inst_16_n15}), .b ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, new_AGEMA_signal_2602, sbox_inst_16_T5}), .c ({new_AGEMA_signal_3210, new_AGEMA_signal_3209, new_AGEMA_signal_3208, sbox_inst_16_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U9 ( .a ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, new_AGEMA_signal_2596, sbox_inst_16_n15}), .b ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, new_AGEMA_signal_3745, sbox_inst_16_n14}), .c ({output0_s3[136], output0_s2[136], output0_s1[136], output0_s0[136]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U8 ( .a ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, new_AGEMA_signal_2593, sbox_inst_16_n13}), .b ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, new_AGEMA_signal_3211, sbox_inst_16_n12}), .c ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, new_AGEMA_signal_3745, sbox_inst_16_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_U7 ( .a ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, new_AGEMA_signal_2605, sbox_inst_16_T6}), .b ({input0_s3[67], input0_s2[67], input0_s1[67], input0_s0[67]}), .c ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, new_AGEMA_signal_3211, sbox_inst_16_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_t5_AND_U1 ( .a ({input0_s3[65], input0_s2[65], input0_s1[65], input0_s0[65]}), .b ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, new_AGEMA_signal_1813, sbox_inst_16_T3}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, new_AGEMA_signal_2602, sbox_inst_16_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_16_t6_AND_U1 ( .a ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, new_AGEMA_signal_1795, sbox_inst_16_L0}), .b ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, new_AGEMA_signal_1807, sbox_inst_16_T1}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, new_AGEMA_signal_2605, sbox_inst_16_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U15 ( .a ({new_AGEMA_signal_1842, new_AGEMA_signal_1841, new_AGEMA_signal_1840, sbox_inst_15_T2}), .b ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, new_AGEMA_signal_3751, sbox_inst_15_n20}), .c ({output0_s3[55], output0_s2[55], output0_s1[55], output0_s0[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U14 ( .a ({new_AGEMA_signal_3222, new_AGEMA_signal_3221, new_AGEMA_signal_3220, sbox_inst_15_n19}), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, new_AGEMA_signal_3217, sbox_inst_15_n18}), .c ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, new_AGEMA_signal_3751, sbox_inst_15_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U13 ( .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, new_AGEMA_signal_1837, sbox_inst_15_T1}), .b ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, new_AGEMA_signal_2617, sbox_inst_15_T5}), .c ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, new_AGEMA_signal_3217, sbox_inst_15_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U11 ( .a ({input0_s3[61], input0_s2[61], input0_s1[61], input0_s0[61]}), .b ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, new_AGEMA_signal_3223, sbox_inst_15_n16}), .c ({output0_s3[95], output0_s2[95], output0_s1[95], output0_s0[95]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U10 ( .a ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, new_AGEMA_signal_2611, sbox_inst_15_n15}), .b ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, new_AGEMA_signal_2617, sbox_inst_15_T5}), .c ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, new_AGEMA_signal_3223, sbox_inst_15_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U9 ( .a ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, new_AGEMA_signal_2611, sbox_inst_15_n15}), .b ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, new_AGEMA_signal_3757, sbox_inst_15_n14}), .c ({output0_s3[135], output0_s2[135], output0_s1[135], output0_s0[135]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U8 ( .a ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, new_AGEMA_signal_2608, sbox_inst_15_n13}), .b ({new_AGEMA_signal_3228, new_AGEMA_signal_3227, new_AGEMA_signal_3226, sbox_inst_15_n12}), .c ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, new_AGEMA_signal_3757, sbox_inst_15_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_U7 ( .a ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, new_AGEMA_signal_2620, sbox_inst_15_T6}), .b ({input0_s3[63], input0_s2[63], input0_s1[63], input0_s0[63]}), .c ({new_AGEMA_signal_3228, new_AGEMA_signal_3227, new_AGEMA_signal_3226, sbox_inst_15_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_t5_AND_U1 ( .a ({input0_s3[61], input0_s2[61], input0_s1[61], input0_s0[61]}), .b ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, new_AGEMA_signal_1843, sbox_inst_15_T3}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, new_AGEMA_signal_2617, sbox_inst_15_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_15_t6_AND_U1 ( .a ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, new_AGEMA_signal_1825, sbox_inst_15_L0}), .b ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, new_AGEMA_signal_1837, sbox_inst_15_T1}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, new_AGEMA_signal_2620, sbox_inst_15_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U15 ( .a ({new_AGEMA_signal_1872, new_AGEMA_signal_1871, new_AGEMA_signal_1870, sbox_inst_14_T2}), .b ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, new_AGEMA_signal_3763, sbox_inst_14_n20}), .c ({output0_s3[54], output0_s2[54], output0_s1[54], output0_s0[54]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U14 ( .a ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, new_AGEMA_signal_3235, sbox_inst_14_n19}), .b ({new_AGEMA_signal_3234, new_AGEMA_signal_3233, new_AGEMA_signal_3232, sbox_inst_14_n18}), .c ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, new_AGEMA_signal_3763, sbox_inst_14_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U13 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, sbox_inst_14_T1}), .b ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, new_AGEMA_signal_2632, sbox_inst_14_T5}), .c ({new_AGEMA_signal_3234, new_AGEMA_signal_3233, new_AGEMA_signal_3232, sbox_inst_14_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U11 ( .a ({input0_s3[57], input0_s2[57], input0_s1[57], input0_s0[57]}), .b ({new_AGEMA_signal_3240, new_AGEMA_signal_3239, new_AGEMA_signal_3238, sbox_inst_14_n16}), .c ({output0_s3[94], output0_s2[94], output0_s1[94], output0_s0[94]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U10 ( .a ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, new_AGEMA_signal_2626, sbox_inst_14_n15}), .b ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, new_AGEMA_signal_2632, sbox_inst_14_T5}), .c ({new_AGEMA_signal_3240, new_AGEMA_signal_3239, new_AGEMA_signal_3238, sbox_inst_14_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U9 ( .a ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, new_AGEMA_signal_2626, sbox_inst_14_n15}), .b ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, new_AGEMA_signal_3769, sbox_inst_14_n14}), .c ({output0_s3[134], output0_s2[134], output0_s1[134], output0_s0[134]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U8 ( .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, new_AGEMA_signal_2623, sbox_inst_14_n13}), .b ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, new_AGEMA_signal_3241, sbox_inst_14_n12}), .c ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, new_AGEMA_signal_3769, sbox_inst_14_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_U7 ( .a ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, new_AGEMA_signal_2635, sbox_inst_14_T6}), .b ({input0_s3[59], input0_s2[59], input0_s1[59], input0_s0[59]}), .c ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, new_AGEMA_signal_3241, sbox_inst_14_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_t5_AND_U1 ( .a ({input0_s3[57], input0_s2[57], input0_s1[57], input0_s0[57]}), .b ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, new_AGEMA_signal_1873, sbox_inst_14_T3}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, new_AGEMA_signal_2632, sbox_inst_14_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_14_t6_AND_U1 ( .a ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, new_AGEMA_signal_1855, sbox_inst_14_L0}), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, new_AGEMA_signal_1867, sbox_inst_14_T1}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, new_AGEMA_signal_2635, sbox_inst_14_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U15 ( .a ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, new_AGEMA_signal_1900, sbox_inst_13_T2}), .b ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, new_AGEMA_signal_3775, sbox_inst_13_n20}), .c ({output0_s3[53], output0_s2[53], output0_s1[53], output0_s0[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U14 ( .a ({new_AGEMA_signal_3252, new_AGEMA_signal_3251, new_AGEMA_signal_3250, sbox_inst_13_n19}), .b ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, new_AGEMA_signal_3247, sbox_inst_13_n18}), .c ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, new_AGEMA_signal_3775, sbox_inst_13_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U13 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, new_AGEMA_signal_1897, sbox_inst_13_T1}), .b ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, new_AGEMA_signal_2647, sbox_inst_13_T5}), .c ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, new_AGEMA_signal_3247, sbox_inst_13_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U11 ( .a ({input0_s3[53], input0_s2[53], input0_s1[53], input0_s0[53]}), .b ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, new_AGEMA_signal_3253, sbox_inst_13_n16}), .c ({output0_s3[93], output0_s2[93], output0_s1[93], output0_s0[93]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U10 ( .a ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, new_AGEMA_signal_2641, sbox_inst_13_n15}), .b ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, new_AGEMA_signal_2647, sbox_inst_13_T5}), .c ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, new_AGEMA_signal_3253, sbox_inst_13_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U9 ( .a ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, new_AGEMA_signal_2641, sbox_inst_13_n15}), .b ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, new_AGEMA_signal_3781, sbox_inst_13_n14}), .c ({output0_s3[133], output0_s2[133], output0_s1[133], output0_s0[133]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U8 ( .a ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, sbox_inst_13_n13}), .b ({new_AGEMA_signal_3258, new_AGEMA_signal_3257, new_AGEMA_signal_3256, sbox_inst_13_n12}), .c ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, new_AGEMA_signal_3781, sbox_inst_13_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_U7 ( .a ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, new_AGEMA_signal_2650, sbox_inst_13_T6}), .b ({input0_s3[55], input0_s2[55], input0_s1[55], input0_s0[55]}), .c ({new_AGEMA_signal_3258, new_AGEMA_signal_3257, new_AGEMA_signal_3256, sbox_inst_13_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_t5_AND_U1 ( .a ({input0_s3[53], input0_s2[53], input0_s1[53], input0_s0[53]}), .b ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, new_AGEMA_signal_1903, sbox_inst_13_T3}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, new_AGEMA_signal_2647, sbox_inst_13_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_13_t6_AND_U1 ( .a ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, new_AGEMA_signal_1885, sbox_inst_13_L0}), .b ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, new_AGEMA_signal_1897, sbox_inst_13_T1}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, new_AGEMA_signal_2650, sbox_inst_13_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U15 ( .a ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, new_AGEMA_signal_1930, sbox_inst_12_T2}), .b ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, new_AGEMA_signal_3787, sbox_inst_12_n20}), .c ({output0_s3[52], output0_s2[52], output0_s1[52], output0_s0[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U14 ( .a ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, new_AGEMA_signal_3265, sbox_inst_12_n19}), .b ({new_AGEMA_signal_3264, new_AGEMA_signal_3263, new_AGEMA_signal_3262, sbox_inst_12_n18}), .c ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, new_AGEMA_signal_3787, sbox_inst_12_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U13 ( .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, sbox_inst_12_T1}), .b ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, new_AGEMA_signal_2662, sbox_inst_12_T5}), .c ({new_AGEMA_signal_3264, new_AGEMA_signal_3263, new_AGEMA_signal_3262, sbox_inst_12_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U11 ( .a ({input0_s3[49], input0_s2[49], input0_s1[49], input0_s0[49]}), .b ({new_AGEMA_signal_3270, new_AGEMA_signal_3269, new_AGEMA_signal_3268, sbox_inst_12_n16}), .c ({output0_s3[92], output0_s2[92], output0_s1[92], output0_s0[92]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U10 ( .a ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, new_AGEMA_signal_2656, sbox_inst_12_n15}), .b ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, new_AGEMA_signal_2662, sbox_inst_12_T5}), .c ({new_AGEMA_signal_3270, new_AGEMA_signal_3269, new_AGEMA_signal_3268, sbox_inst_12_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U9 ( .a ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, new_AGEMA_signal_2656, sbox_inst_12_n15}), .b ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, new_AGEMA_signal_3793, sbox_inst_12_n14}), .c ({output0_s3[132], output0_s2[132], output0_s1[132], output0_s0[132]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U8 ( .a ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, new_AGEMA_signal_2653, sbox_inst_12_n13}), .b ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, new_AGEMA_signal_3271, sbox_inst_12_n12}), .c ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, new_AGEMA_signal_3793, sbox_inst_12_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_U7 ( .a ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, new_AGEMA_signal_2665, sbox_inst_12_T6}), .b ({input0_s3[51], input0_s2[51], input0_s1[51], input0_s0[51]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, new_AGEMA_signal_3271, sbox_inst_12_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_t5_AND_U1 ( .a ({input0_s3[49], input0_s2[49], input0_s1[49], input0_s0[49]}), .b ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, new_AGEMA_signal_1933, sbox_inst_12_T3}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, new_AGEMA_signal_2662, sbox_inst_12_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_12_t6_AND_U1 ( .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, new_AGEMA_signal_1915, sbox_inst_12_L0}), .b ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, new_AGEMA_signal_1927, sbox_inst_12_T1}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, new_AGEMA_signal_2665, sbox_inst_12_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U15 ( .a ({new_AGEMA_signal_1962, new_AGEMA_signal_1961, new_AGEMA_signal_1960, sbox_inst_11_T2}), .b ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, new_AGEMA_signal_3799, sbox_inst_11_n20}), .c ({output0_s3[51], output0_s2[51], output0_s1[51], output0_s0[51]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U14 ( .a ({new_AGEMA_signal_3282, new_AGEMA_signal_3281, new_AGEMA_signal_3280, sbox_inst_11_n19}), .b ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, new_AGEMA_signal_3277, sbox_inst_11_n18}), .c ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, new_AGEMA_signal_3799, sbox_inst_11_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U13 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, sbox_inst_11_T1}), .b ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, new_AGEMA_signal_2677, sbox_inst_11_T5}), .c ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, new_AGEMA_signal_3277, sbox_inst_11_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U11 ( .a ({input0_s3[45], input0_s2[45], input0_s1[45], input0_s0[45]}), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, new_AGEMA_signal_3283, sbox_inst_11_n16}), .c ({output0_s3[91], output0_s2[91], output0_s1[91], output0_s0[91]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U10 ( .a ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, new_AGEMA_signal_2671, sbox_inst_11_n15}), .b ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, new_AGEMA_signal_2677, sbox_inst_11_T5}), .c ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, new_AGEMA_signal_3283, sbox_inst_11_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U9 ( .a ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, new_AGEMA_signal_2671, sbox_inst_11_n15}), .b ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, new_AGEMA_signal_3805, sbox_inst_11_n14}), .c ({output0_s3[131], output0_s2[131], output0_s1[131], output0_s0[131]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U8 ( .a ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, new_AGEMA_signal_2668, sbox_inst_11_n13}), .b ({new_AGEMA_signal_3288, new_AGEMA_signal_3287, new_AGEMA_signal_3286, sbox_inst_11_n12}), .c ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, new_AGEMA_signal_3805, sbox_inst_11_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_U7 ( .a ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, new_AGEMA_signal_2680, sbox_inst_11_T6}), .b ({input0_s3[47], input0_s2[47], input0_s1[47], input0_s0[47]}), .c ({new_AGEMA_signal_3288, new_AGEMA_signal_3287, new_AGEMA_signal_3286, sbox_inst_11_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_t5_AND_U1 ( .a ({input0_s3[45], input0_s2[45], input0_s1[45], input0_s0[45]}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, new_AGEMA_signal_1963, sbox_inst_11_T3}), .clk (clk), .r ({Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, new_AGEMA_signal_2677, sbox_inst_11_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_11_t6_AND_U1 ( .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, new_AGEMA_signal_1945, sbox_inst_11_L0}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, new_AGEMA_signal_1957, sbox_inst_11_T1}), .clk (clk), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, new_AGEMA_signal_2680, sbox_inst_11_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U15 ( .a ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, new_AGEMA_signal_1990, sbox_inst_10_T2}), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, new_AGEMA_signal_3811, sbox_inst_10_n20}), .c ({output0_s3[50], output0_s2[50], output0_s1[50], output0_s0[50]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U14 ( .a ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, new_AGEMA_signal_3295, sbox_inst_10_n19}), .b ({new_AGEMA_signal_3294, new_AGEMA_signal_3293, new_AGEMA_signal_3292, sbox_inst_10_n18}), .c ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, new_AGEMA_signal_3811, sbox_inst_10_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U13 ( .a ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, new_AGEMA_signal_1987, sbox_inst_10_T1}), .b ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, new_AGEMA_signal_2692, sbox_inst_10_T5}), .c ({new_AGEMA_signal_3294, new_AGEMA_signal_3293, new_AGEMA_signal_3292, sbox_inst_10_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U11 ( .a ({input0_s3[41], input0_s2[41], input0_s1[41], input0_s0[41]}), .b ({new_AGEMA_signal_3300, new_AGEMA_signal_3299, new_AGEMA_signal_3298, sbox_inst_10_n16}), .c ({output0_s3[90], output0_s2[90], output0_s1[90], output0_s0[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U10 ( .a ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, sbox_inst_10_n15}), .b ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, new_AGEMA_signal_2692, sbox_inst_10_T5}), .c ({new_AGEMA_signal_3300, new_AGEMA_signal_3299, new_AGEMA_signal_3298, sbox_inst_10_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U9 ( .a ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, sbox_inst_10_n15}), .b ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, new_AGEMA_signal_3817, sbox_inst_10_n14}), .c ({output0_s3[130], output0_s2[130], output0_s1[130], output0_s0[130]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U8 ( .a ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, new_AGEMA_signal_2683, sbox_inst_10_n13}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, new_AGEMA_signal_3301, sbox_inst_10_n12}), .c ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, new_AGEMA_signal_3817, sbox_inst_10_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_U7 ( .a ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, new_AGEMA_signal_2695, sbox_inst_10_T6}), .b ({input0_s3[43], input0_s2[43], input0_s1[43], input0_s0[43]}), .c ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, new_AGEMA_signal_3301, sbox_inst_10_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_t5_AND_U1 ( .a ({input0_s3[41], input0_s2[41], input0_s1[41], input0_s0[41]}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, new_AGEMA_signal_1993, sbox_inst_10_T3}), .clk (clk), .r ({Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, new_AGEMA_signal_2692, sbox_inst_10_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_10_t6_AND_U1 ( .a ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, new_AGEMA_signal_1975, sbox_inst_10_L0}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, new_AGEMA_signal_1987, sbox_inst_10_T1}), .clk (clk), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, new_AGEMA_signal_2695, sbox_inst_10_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U15 ( .a ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, new_AGEMA_signal_2020, sbox_inst_9_T2}), .b ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, new_AGEMA_signal_3823, sbox_inst_9_n20}), .c ({output0_s3[49], output0_s2[49], output0_s1[49], output0_s0[49]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U14 ( .a ({new_AGEMA_signal_3312, new_AGEMA_signal_3311, new_AGEMA_signal_3310, sbox_inst_9_n19}), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, new_AGEMA_signal_3307, sbox_inst_9_n18}), .c ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, new_AGEMA_signal_3823, sbox_inst_9_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U13 ( .a ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, new_AGEMA_signal_2017, sbox_inst_9_T1}), .b ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, new_AGEMA_signal_2707, sbox_inst_9_T5}), .c ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, new_AGEMA_signal_3307, sbox_inst_9_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U11 ( .a ({input0_s3[37], input0_s2[37], input0_s1[37], input0_s0[37]}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, new_AGEMA_signal_3313, sbox_inst_9_n16}), .c ({output0_s3[89], output0_s2[89], output0_s1[89], output0_s0[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U10 ( .a ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, new_AGEMA_signal_2701, sbox_inst_9_n15}), .b ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, new_AGEMA_signal_2707, sbox_inst_9_T5}), .c ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, new_AGEMA_signal_3313, sbox_inst_9_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U9 ( .a ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, new_AGEMA_signal_2701, sbox_inst_9_n15}), .b ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, new_AGEMA_signal_3829, sbox_inst_9_n14}), .c ({output0_s3[129], output0_s2[129], output0_s1[129], output0_s0[129]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U8 ( .a ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, new_AGEMA_signal_2698, sbox_inst_9_n13}), .b ({new_AGEMA_signal_3318, new_AGEMA_signal_3317, new_AGEMA_signal_3316, sbox_inst_9_n12}), .c ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, new_AGEMA_signal_3829, sbox_inst_9_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_U7 ( .a ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, new_AGEMA_signal_2710, sbox_inst_9_T6}), .b ({input0_s3[39], input0_s2[39], input0_s1[39], input0_s0[39]}), .c ({new_AGEMA_signal_3318, new_AGEMA_signal_3317, new_AGEMA_signal_3316, sbox_inst_9_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_t5_AND_U1 ( .a ({input0_s3[37], input0_s2[37], input0_s1[37], input0_s0[37]}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, new_AGEMA_signal_2023, sbox_inst_9_T3}), .clk (clk), .r ({Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, new_AGEMA_signal_2707, sbox_inst_9_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_9_t6_AND_U1 ( .a ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, new_AGEMA_signal_2005, sbox_inst_9_L0}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, new_AGEMA_signal_2017, sbox_inst_9_T1}), .clk (clk), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, new_AGEMA_signal_2710, sbox_inst_9_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U15 ( .a ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, new_AGEMA_signal_2050, sbox_inst_8_T2}), .b ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, new_AGEMA_signal_3835, sbox_inst_8_n20}), .c ({output0_s3[48], output0_s2[48], output0_s1[48], output0_s0[48]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U14 ( .a ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, new_AGEMA_signal_3325, sbox_inst_8_n19}), .b ({new_AGEMA_signal_3324, new_AGEMA_signal_3323, new_AGEMA_signal_3322, sbox_inst_8_n18}), .c ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, new_AGEMA_signal_3835, sbox_inst_8_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U13 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, sbox_inst_8_T1}), .b ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, new_AGEMA_signal_2722, sbox_inst_8_T5}), .c ({new_AGEMA_signal_3324, new_AGEMA_signal_3323, new_AGEMA_signal_3322, sbox_inst_8_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U11 ( .a ({input0_s3[33], input0_s2[33], input0_s1[33], input0_s0[33]}), .b ({new_AGEMA_signal_3330, new_AGEMA_signal_3329, new_AGEMA_signal_3328, sbox_inst_8_n16}), .c ({output0_s3[88], output0_s2[88], output0_s1[88], output0_s0[88]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U10 ( .a ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, new_AGEMA_signal_2716, sbox_inst_8_n15}), .b ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, new_AGEMA_signal_2722, sbox_inst_8_T5}), .c ({new_AGEMA_signal_3330, new_AGEMA_signal_3329, new_AGEMA_signal_3328, sbox_inst_8_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U9 ( .a ({new_AGEMA_signal_2718, new_AGEMA_signal_2717, new_AGEMA_signal_2716, sbox_inst_8_n15}), .b ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, new_AGEMA_signal_3841, sbox_inst_8_n14}), .c ({output0_s3[128], output0_s2[128], output0_s1[128], output0_s0[128]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U8 ( .a ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, new_AGEMA_signal_2713, sbox_inst_8_n13}), .b ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, new_AGEMA_signal_3331, sbox_inst_8_n12}), .c ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, new_AGEMA_signal_3841, sbox_inst_8_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_U7 ( .a ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, new_AGEMA_signal_2725, sbox_inst_8_T6}), .b ({input0_s3[35], input0_s2[35], input0_s1[35], input0_s0[35]}), .c ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, new_AGEMA_signal_3331, sbox_inst_8_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_t5_AND_U1 ( .a ({input0_s3[33], input0_s2[33], input0_s1[33], input0_s0[33]}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, new_AGEMA_signal_2053, sbox_inst_8_T3}), .clk (clk), .r ({Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, new_AGEMA_signal_2722, sbox_inst_8_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_8_t6_AND_U1 ( .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, new_AGEMA_signal_2035, sbox_inst_8_L0}), .b ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, new_AGEMA_signal_2047, sbox_inst_8_T1}), .clk (clk), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, new_AGEMA_signal_2725, sbox_inst_8_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U15 ( .a ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, new_AGEMA_signal_2080, sbox_inst_7_T2}), .b ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, new_AGEMA_signal_3847, sbox_inst_7_n20}), .c ({output0_s3[47], output0_s2[47], output0_s1[47], output0_s0[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U14 ( .a ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, new_AGEMA_signal_3340, sbox_inst_7_n19}), .b ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, new_AGEMA_signal_3337, sbox_inst_7_n18}), .c ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, new_AGEMA_signal_3847, sbox_inst_7_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U13 ( .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, new_AGEMA_signal_2077, sbox_inst_7_T1}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, new_AGEMA_signal_2737, sbox_inst_7_T5}), .c ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, new_AGEMA_signal_3337, sbox_inst_7_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U11 ( .a ({input0_s3[29], input0_s2[29], input0_s1[29], input0_s0[29]}), .b ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, new_AGEMA_signal_3343, sbox_inst_7_n16}), .c ({output0_s3[87], output0_s2[87], output0_s1[87], output0_s0[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U10 ( .a ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, new_AGEMA_signal_2731, sbox_inst_7_n15}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, new_AGEMA_signal_2737, sbox_inst_7_T5}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, new_AGEMA_signal_3343, sbox_inst_7_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U9 ( .a ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, new_AGEMA_signal_2731, sbox_inst_7_n15}), .b ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, new_AGEMA_signal_3853, sbox_inst_7_n14}), .c ({output0_s3[127], output0_s2[127], output0_s1[127], output0_s0[127]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U8 ( .a ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, new_AGEMA_signal_2728, sbox_inst_7_n13}), .b ({new_AGEMA_signal_3348, new_AGEMA_signal_3347, new_AGEMA_signal_3346, sbox_inst_7_n12}), .c ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, new_AGEMA_signal_3853, sbox_inst_7_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_U7 ( .a ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, new_AGEMA_signal_2740, sbox_inst_7_T6}), .b ({input0_s3[31], input0_s2[31], input0_s1[31], input0_s0[31]}), .c ({new_AGEMA_signal_3348, new_AGEMA_signal_3347, new_AGEMA_signal_3346, sbox_inst_7_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_t5_AND_U1 ( .a ({input0_s3[29], input0_s2[29], input0_s1[29], input0_s0[29]}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, new_AGEMA_signal_2083, sbox_inst_7_T3}), .clk (clk), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, new_AGEMA_signal_2737, sbox_inst_7_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_7_t6_AND_U1 ( .a ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, new_AGEMA_signal_2065, sbox_inst_7_L0}), .b ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, new_AGEMA_signal_2077, sbox_inst_7_T1}), .clk (clk), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, new_AGEMA_signal_2740, sbox_inst_7_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U15 ( .a ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, new_AGEMA_signal_2110, sbox_inst_6_T2}), .b ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, new_AGEMA_signal_3859, sbox_inst_6_n20}), .c ({output0_s3[46], output0_s2[46], output0_s1[46], output0_s0[46]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U14 ( .a ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, new_AGEMA_signal_3355, sbox_inst_6_n19}), .b ({new_AGEMA_signal_3354, new_AGEMA_signal_3353, new_AGEMA_signal_3352, sbox_inst_6_n18}), .c ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, new_AGEMA_signal_3859, sbox_inst_6_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U13 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, sbox_inst_6_T1}), .b ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, new_AGEMA_signal_2752, sbox_inst_6_T5}), .c ({new_AGEMA_signal_3354, new_AGEMA_signal_3353, new_AGEMA_signal_3352, sbox_inst_6_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U11 ( .a ({input0_s3[25], input0_s2[25], input0_s1[25], input0_s0[25]}), .b ({new_AGEMA_signal_3360, new_AGEMA_signal_3359, new_AGEMA_signal_3358, sbox_inst_6_n16}), .c ({output0_s3[86], output0_s2[86], output0_s1[86], output0_s0[86]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U10 ( .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, new_AGEMA_signal_2746, sbox_inst_6_n15}), .b ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, new_AGEMA_signal_2752, sbox_inst_6_T5}), .c ({new_AGEMA_signal_3360, new_AGEMA_signal_3359, new_AGEMA_signal_3358, sbox_inst_6_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U9 ( .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, new_AGEMA_signal_2746, sbox_inst_6_n15}), .b ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, new_AGEMA_signal_3865, sbox_inst_6_n14}), .c ({output0_s3[126], output0_s2[126], output0_s1[126], output0_s0[126]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U8 ( .a ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, new_AGEMA_signal_2743, sbox_inst_6_n13}), .b ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, new_AGEMA_signal_3361, sbox_inst_6_n12}), .c ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, new_AGEMA_signal_3865, sbox_inst_6_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_U7 ( .a ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, new_AGEMA_signal_2755, sbox_inst_6_T6}), .b ({input0_s3[27], input0_s2[27], input0_s1[27], input0_s0[27]}), .c ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, new_AGEMA_signal_3361, sbox_inst_6_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_t5_AND_U1 ( .a ({input0_s3[25], input0_s2[25], input0_s1[25], input0_s0[25]}), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, new_AGEMA_signal_2113, sbox_inst_6_T3}), .clk (clk), .r ({Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_2754, new_AGEMA_signal_2753, new_AGEMA_signal_2752, sbox_inst_6_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_6_t6_AND_U1 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, new_AGEMA_signal_2095, sbox_inst_6_L0}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, new_AGEMA_signal_2107, sbox_inst_6_T1}), .clk (clk), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, new_AGEMA_signal_2755, sbox_inst_6_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U15 ( .a ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, new_AGEMA_signal_2140, sbox_inst_5_T2}), .b ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, new_AGEMA_signal_3871, sbox_inst_5_n20}), .c ({output0_s3[45], output0_s2[45], output0_s1[45], output0_s0[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U14 ( .a ({new_AGEMA_signal_3372, new_AGEMA_signal_3371, new_AGEMA_signal_3370, sbox_inst_5_n19}), .b ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, new_AGEMA_signal_3367, sbox_inst_5_n18}), .c ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, new_AGEMA_signal_3871, sbox_inst_5_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U13 ( .a ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, sbox_inst_5_T1}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, new_AGEMA_signal_2767, sbox_inst_5_T5}), .c ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, new_AGEMA_signal_3367, sbox_inst_5_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U11 ( .a ({input0_s3[21], input0_s2[21], input0_s1[21], input0_s0[21]}), .b ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, new_AGEMA_signal_3373, sbox_inst_5_n16}), .c ({output0_s3[85], output0_s2[85], output0_s1[85], output0_s0[85]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U10 ( .a ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, new_AGEMA_signal_2761, sbox_inst_5_n15}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, new_AGEMA_signal_2767, sbox_inst_5_T5}), .c ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, new_AGEMA_signal_3373, sbox_inst_5_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U9 ( .a ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, new_AGEMA_signal_2761, sbox_inst_5_n15}), .b ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, new_AGEMA_signal_3877, sbox_inst_5_n14}), .c ({output0_s3[125], output0_s2[125], output0_s1[125], output0_s0[125]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U8 ( .a ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, new_AGEMA_signal_2758, sbox_inst_5_n13}), .b ({new_AGEMA_signal_3378, new_AGEMA_signal_3377, new_AGEMA_signal_3376, sbox_inst_5_n12}), .c ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, new_AGEMA_signal_3877, sbox_inst_5_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_U7 ( .a ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, new_AGEMA_signal_2770, sbox_inst_5_T6}), .b ({input0_s3[23], input0_s2[23], input0_s1[23], input0_s0[23]}), .c ({new_AGEMA_signal_3378, new_AGEMA_signal_3377, new_AGEMA_signal_3376, sbox_inst_5_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_t5_AND_U1 ( .a ({input0_s3[21], input0_s2[21], input0_s1[21], input0_s0[21]}), .b ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, new_AGEMA_signal_2143, sbox_inst_5_T3}), .clk (clk), .r ({Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, new_AGEMA_signal_2767, sbox_inst_5_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_5_t6_AND_U1 ( .a ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, new_AGEMA_signal_2125, sbox_inst_5_L0}), .b ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, new_AGEMA_signal_2137, sbox_inst_5_T1}), .clk (clk), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, new_AGEMA_signal_2770, sbox_inst_5_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U15 ( .a ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, new_AGEMA_signal_2170, sbox_inst_4_T2}), .b ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, new_AGEMA_signal_3883, sbox_inst_4_n20}), .c ({output0_s3[44], output0_s2[44], output0_s1[44], output0_s0[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U14 ( .a ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, new_AGEMA_signal_3385, sbox_inst_4_n19}), .b ({new_AGEMA_signal_3384, new_AGEMA_signal_3383, new_AGEMA_signal_3382, sbox_inst_4_n18}), .c ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, new_AGEMA_signal_3883, sbox_inst_4_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U13 ( .a ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, sbox_inst_4_T1}), .b ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, new_AGEMA_signal_2782, sbox_inst_4_T5}), .c ({new_AGEMA_signal_3384, new_AGEMA_signal_3383, new_AGEMA_signal_3382, sbox_inst_4_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U11 ( .a ({input0_s3[17], input0_s2[17], input0_s1[17], input0_s0[17]}), .b ({new_AGEMA_signal_3390, new_AGEMA_signal_3389, new_AGEMA_signal_3388, sbox_inst_4_n16}), .c ({output0_s3[84], output0_s2[84], output0_s1[84], output0_s0[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U10 ( .a ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, new_AGEMA_signal_2776, sbox_inst_4_n15}), .b ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, new_AGEMA_signal_2782, sbox_inst_4_T5}), .c ({new_AGEMA_signal_3390, new_AGEMA_signal_3389, new_AGEMA_signal_3388, sbox_inst_4_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U9 ( .a ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, new_AGEMA_signal_2776, sbox_inst_4_n15}), .b ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, new_AGEMA_signal_3889, sbox_inst_4_n14}), .c ({output0_s3[124], output0_s2[124], output0_s1[124], output0_s0[124]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U8 ( .a ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, new_AGEMA_signal_2773, sbox_inst_4_n13}), .b ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, new_AGEMA_signal_3391, sbox_inst_4_n12}), .c ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, new_AGEMA_signal_3889, sbox_inst_4_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_U7 ( .a ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, new_AGEMA_signal_2785, sbox_inst_4_T6}), .b ({input0_s3[19], input0_s2[19], input0_s1[19], input0_s0[19]}), .c ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, new_AGEMA_signal_3391, sbox_inst_4_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_t5_AND_U1 ( .a ({input0_s3[17], input0_s2[17], input0_s1[17], input0_s0[17]}), .b ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, new_AGEMA_signal_2173, sbox_inst_4_T3}), .clk (clk), .r ({Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, new_AGEMA_signal_2782, sbox_inst_4_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_4_t6_AND_U1 ( .a ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, new_AGEMA_signal_2155, sbox_inst_4_L0}), .b ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, new_AGEMA_signal_2167, sbox_inst_4_T1}), .clk (clk), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, new_AGEMA_signal_2785, sbox_inst_4_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U15 ( .a ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, new_AGEMA_signal_2200, sbox_inst_3_T2}), .b ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, new_AGEMA_signal_3895, sbox_inst_3_n20}), .c ({output0_s3[43], output0_s2[43], output0_s1[43], output0_s0[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U14 ( .a ({new_AGEMA_signal_3402, new_AGEMA_signal_3401, new_AGEMA_signal_3400, sbox_inst_3_n19}), .b ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, new_AGEMA_signal_3397, sbox_inst_3_n18}), .c ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, new_AGEMA_signal_3895, sbox_inst_3_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U13 ( .a ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, new_AGEMA_signal_2197, sbox_inst_3_T1}), .b ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, new_AGEMA_signal_2797, sbox_inst_3_T5}), .c ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, new_AGEMA_signal_3397, sbox_inst_3_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U11 ( .a ({input0_s3[13], input0_s2[13], input0_s1[13], input0_s0[13]}), .b ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, new_AGEMA_signal_3403, sbox_inst_3_n16}), .c ({output0_s3[83], output0_s2[83], output0_s1[83], output0_s0[83]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U10 ( .a ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, new_AGEMA_signal_2791, sbox_inst_3_n15}), .b ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, new_AGEMA_signal_2797, sbox_inst_3_T5}), .c ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, new_AGEMA_signal_3403, sbox_inst_3_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U9 ( .a ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, new_AGEMA_signal_2791, sbox_inst_3_n15}), .b ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, new_AGEMA_signal_3901, sbox_inst_3_n14}), .c ({output0_s3[123], output0_s2[123], output0_s1[123], output0_s0[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U8 ( .a ({new_AGEMA_signal_2790, new_AGEMA_signal_2789, new_AGEMA_signal_2788, sbox_inst_3_n13}), .b ({new_AGEMA_signal_3408, new_AGEMA_signal_3407, new_AGEMA_signal_3406, sbox_inst_3_n12}), .c ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, new_AGEMA_signal_3901, sbox_inst_3_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_U7 ( .a ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, new_AGEMA_signal_2800, sbox_inst_3_T6}), .b ({input0_s3[15], input0_s2[15], input0_s1[15], input0_s0[15]}), .c ({new_AGEMA_signal_3408, new_AGEMA_signal_3407, new_AGEMA_signal_3406, sbox_inst_3_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_t5_AND_U1 ( .a ({input0_s3[13], input0_s2[13], input0_s1[13], input0_s0[13]}), .b ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, new_AGEMA_signal_2203, sbox_inst_3_T3}), .clk (clk), .r ({Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, new_AGEMA_signal_2797, sbox_inst_3_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_3_t6_AND_U1 ( .a ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, new_AGEMA_signal_2185, sbox_inst_3_L0}), .b ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, new_AGEMA_signal_2197, sbox_inst_3_T1}), .clk (clk), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, new_AGEMA_signal_2800, sbox_inst_3_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U15 ( .a ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, new_AGEMA_signal_2230, sbox_inst_2_T2}), .b ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, new_AGEMA_signal_3907, sbox_inst_2_n20}), .c ({output0_s3[42], output0_s2[42], output0_s1[42], output0_s0[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U14 ( .a ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, new_AGEMA_signal_3415, sbox_inst_2_n19}), .b ({new_AGEMA_signal_3414, new_AGEMA_signal_3413, new_AGEMA_signal_3412, sbox_inst_2_n18}), .c ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, new_AGEMA_signal_3907, sbox_inst_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U13 ( .a ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, new_AGEMA_signal_2227, sbox_inst_2_T1}), .b ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, new_AGEMA_signal_2812, sbox_inst_2_T5}), .c ({new_AGEMA_signal_3414, new_AGEMA_signal_3413, new_AGEMA_signal_3412, sbox_inst_2_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U11 ( .a ({input0_s3[9], input0_s2[9], input0_s1[9], input0_s0[9]}), .b ({new_AGEMA_signal_3420, new_AGEMA_signal_3419, new_AGEMA_signal_3418, sbox_inst_2_n16}), .c ({output0_s3[82], output0_s2[82], output0_s1[82], output0_s0[82]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U10 ( .a ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, new_AGEMA_signal_2806, sbox_inst_2_n15}), .b ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, new_AGEMA_signal_2812, sbox_inst_2_T5}), .c ({new_AGEMA_signal_3420, new_AGEMA_signal_3419, new_AGEMA_signal_3418, sbox_inst_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U9 ( .a ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, new_AGEMA_signal_2806, sbox_inst_2_n15}), .b ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, new_AGEMA_signal_3913, sbox_inst_2_n14}), .c ({output0_s3[122], output0_s2[122], output0_s1[122], output0_s0[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U8 ( .a ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, new_AGEMA_signal_2803, sbox_inst_2_n13}), .b ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, new_AGEMA_signal_3421, sbox_inst_2_n12}), .c ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, new_AGEMA_signal_3913, sbox_inst_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_U7 ( .a ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, new_AGEMA_signal_2815, sbox_inst_2_T6}), .b ({input0_s3[11], input0_s2[11], input0_s1[11], input0_s0[11]}), .c ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, new_AGEMA_signal_3421, sbox_inst_2_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_t5_AND_U1 ( .a ({input0_s3[9], input0_s2[9], input0_s1[9], input0_s0[9]}), .b ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, new_AGEMA_signal_2233, sbox_inst_2_T3}), .clk (clk), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, new_AGEMA_signal_2812, sbox_inst_2_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_2_t6_AND_U1 ( .a ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, new_AGEMA_signal_2215, sbox_inst_2_L0}), .b ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, new_AGEMA_signal_2227, sbox_inst_2_T1}), .clk (clk), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, new_AGEMA_signal_2815, sbox_inst_2_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U15 ( .a ({new_AGEMA_signal_2832, new_AGEMA_signal_2831, new_AGEMA_signal_2830, sbox_inst_1_T2}), .b ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, new_AGEMA_signal_4189, sbox_inst_1_n20}), .c ({output0_s3[41], output0_s2[41], output0_s1[41], output0_s0[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U14 ( .a ({new_AGEMA_signal_3924, new_AGEMA_signal_3923, new_AGEMA_signal_3922, sbox_inst_1_n19}), .b ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, new_AGEMA_signal_3919, sbox_inst_1_n18}), .c ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, new_AGEMA_signal_4189, sbox_inst_1_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U13 ( .a ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, new_AGEMA_signal_2827, sbox_inst_1_T1}), .b ({new_AGEMA_signal_3438, new_AGEMA_signal_3437, new_AGEMA_signal_3436, sbox_inst_1_T5}), .c ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, new_AGEMA_signal_3919, sbox_inst_1_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U11 ( .a ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, input_array_5}), .b ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, new_AGEMA_signal_3925, sbox_inst_1_n16}), .c ({output0_s3[81], output0_s2[81], output0_s1[81], output0_s0[81]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U10 ( .a ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, new_AGEMA_signal_3430, sbox_inst_1_n15}), .b ({new_AGEMA_signal_3438, new_AGEMA_signal_3437, new_AGEMA_signal_3436, sbox_inst_1_T5}), .c ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, new_AGEMA_signal_3925, sbox_inst_1_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U9 ( .a ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, new_AGEMA_signal_3430, sbox_inst_1_n15}), .b ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, new_AGEMA_signal_4195, sbox_inst_1_n14}), .c ({output0_s3[121], output0_s2[121], output0_s1[121], output0_s0[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U8 ( .a ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, new_AGEMA_signal_3427, sbox_inst_1_n13}), .b ({new_AGEMA_signal_3930, new_AGEMA_signal_3929, new_AGEMA_signal_3928, sbox_inst_1_n12}), .c ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, new_AGEMA_signal_4195, sbox_inst_1_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_U7 ( .a ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, new_AGEMA_signal_3439, sbox_inst_1_T6}), .b ({input0_s3[7], input0_s2[7], input0_s1[7], input0_s0[7]}), .c ({new_AGEMA_signal_3930, new_AGEMA_signal_3929, new_AGEMA_signal_3928, sbox_inst_1_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_t5_AND_U1 ( .a ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, new_AGEMA_signal_1096, input_array_5}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, new_AGEMA_signal_2833, sbox_inst_1_T3}), .clk (clk), .r ({Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({new_AGEMA_signal_3438, new_AGEMA_signal_3437, new_AGEMA_signal_3436, sbox_inst_1_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_1_t6_AND_U1 ( .a ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, new_AGEMA_signal_2818, sbox_inst_1_L0}), .b ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, new_AGEMA_signal_2827, sbox_inst_1_T1}), .clk (clk), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, new_AGEMA_signal_3439, sbox_inst_1_T6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U15 ( .a ({new_AGEMA_signal_2850, new_AGEMA_signal_2849, new_AGEMA_signal_2848, sbox_inst_0_T2}), .b ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, new_AGEMA_signal_4201, sbox_inst_0_n20}), .c ({output0_s3[40], output0_s2[40], output0_s1[40], output0_s0[40]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U14 ( .a ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, new_AGEMA_signal_3937, sbox_inst_0_n19}), .b ({new_AGEMA_signal_3936, new_AGEMA_signal_3935, new_AGEMA_signal_3934, sbox_inst_0_n18}), .c ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, new_AGEMA_signal_4201, sbox_inst_0_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U13 ( .a ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, new_AGEMA_signal_2845, sbox_inst_0_T1}), .b ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, new_AGEMA_signal_3451, sbox_inst_0_T5}), .c ({new_AGEMA_signal_3936, new_AGEMA_signal_3935, new_AGEMA_signal_3934, sbox_inst_0_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U11 ( .a ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, input_array_1}), .b ({new_AGEMA_signal_3942, new_AGEMA_signal_3941, new_AGEMA_signal_3940, sbox_inst_0_n16}), .c ({output0_s3[80], output0_s2[80], output0_s1[80], output0_s0[80]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U10 ( .a ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, new_AGEMA_signal_3445, sbox_inst_0_n15}), .b ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, new_AGEMA_signal_3451, sbox_inst_0_T5}), .c ({new_AGEMA_signal_3942, new_AGEMA_signal_3941, new_AGEMA_signal_3940, sbox_inst_0_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U9 ( .a ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, new_AGEMA_signal_3445, sbox_inst_0_n15}), .b ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, new_AGEMA_signal_4207, sbox_inst_0_n14}), .c ({output0_s3[120], output0_s2[120], output0_s1[120], output0_s0[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U8 ( .a ({new_AGEMA_signal_3444, new_AGEMA_signal_3443, new_AGEMA_signal_3442, sbox_inst_0_n13}), .b ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, new_AGEMA_signal_3943, sbox_inst_0_n12}), .c ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, new_AGEMA_signal_4207, sbox_inst_0_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_U7 ( .a ({new_AGEMA_signal_3456, new_AGEMA_signal_3455, new_AGEMA_signal_3454, sbox_inst_0_T6}), .b ({new_AGEMA_signal_1116, new_AGEMA_signal_1115, new_AGEMA_signal_1114, input_array_3}), .c ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, new_AGEMA_signal_3943, sbox_inst_0_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_t5_AND_U1 ( .a ({new_AGEMA_signal_1080, new_AGEMA_signal_1079, new_AGEMA_signal_1078, input_array_1}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, new_AGEMA_signal_2851, sbox_inst_0_T3}), .clk (clk), .r ({Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, new_AGEMA_signal_3451, sbox_inst_0_T5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) sbox_inst_0_t6_AND_U1 ( .a ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, new_AGEMA_signal_2839, sbox_inst_0_L0}), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, new_AGEMA_signal_2845, sbox_inst_0_T1}), .clk (clk), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({new_AGEMA_signal_3456, new_AGEMA_signal_3455, new_AGEMA_signal_3454, sbox_inst_0_T6}) ) ;

endmodule
