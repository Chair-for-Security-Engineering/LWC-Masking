/* modified netlist. Source: module elephant_perm in file ./test/elephant_perm.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module elephant_perm_HPC2_ClockGating_d2 (input0_s0, lfsr, rev_lfsr, clk, input0_s1, input0_s2, Fresh, /*rst,*/ output0_s0, output0_s1, output0_s2/*, Synch*/);
    input [159:0] input0_s0 ;
    input [6:0] lfsr ;
    input [6:0] rev_lfsr ;
    input clk ;
    input [159:0] input0_s1 ;
    input [159:0] input0_s2 ;
    //input rst ;
    input [839:0] Fresh ;
    output [159:0] output0_s0 ;
    output [159:0] output0_s1 ;
    output [159:0] output0_s2 ;
    //output Synch ;
    wire input_array_6 ;
    wire input_array_5 ;
    wire input_array_4 ;
    wire input_array_3 ;
    wire input_array_2 ;
    wire input_array_1 ;
    wire input_array_0 ;
    wire sbox_inst_39_n20 ;
    wire sbox_inst_39_n19 ;
    wire sbox_inst_39_n18 ;
    wire sbox_inst_39_n17 ;
    wire sbox_inst_39_n16 ;
    wire sbox_inst_39_n15 ;
    wire sbox_inst_39_n14 ;
    wire sbox_inst_39_n13 ;
    wire sbox_inst_39_n12 ;
    wire sbox_inst_39_n11 ;
    wire sbox_inst_39_T6 ;
    wire sbox_inst_39_L0 ;
    wire sbox_inst_39_T5 ;
    wire sbox_inst_39_T4 ;
    wire sbox_inst_39_T3 ;
    wire sbox_inst_39_T2 ;
    wire sbox_inst_39_T1 ;
    wire sbox_inst_39_T0 ;
    wire sbox_inst_38_n20 ;
    wire sbox_inst_38_n19 ;
    wire sbox_inst_38_n18 ;
    wire sbox_inst_38_n17 ;
    wire sbox_inst_38_n16 ;
    wire sbox_inst_38_n15 ;
    wire sbox_inst_38_n14 ;
    wire sbox_inst_38_n13 ;
    wire sbox_inst_38_n12 ;
    wire sbox_inst_38_n11 ;
    wire sbox_inst_38_T6 ;
    wire sbox_inst_38_L0 ;
    wire sbox_inst_38_T5 ;
    wire sbox_inst_38_T4 ;
    wire sbox_inst_38_T3 ;
    wire sbox_inst_38_T2 ;
    wire sbox_inst_38_T1 ;
    wire sbox_inst_38_T0 ;
    wire sbox_inst_37_n20 ;
    wire sbox_inst_37_n19 ;
    wire sbox_inst_37_n18 ;
    wire sbox_inst_37_n17 ;
    wire sbox_inst_37_n16 ;
    wire sbox_inst_37_n15 ;
    wire sbox_inst_37_n14 ;
    wire sbox_inst_37_n13 ;
    wire sbox_inst_37_n12 ;
    wire sbox_inst_37_n11 ;
    wire sbox_inst_37_T6 ;
    wire sbox_inst_37_L0 ;
    wire sbox_inst_37_T5 ;
    wire sbox_inst_37_T4 ;
    wire sbox_inst_37_T3 ;
    wire sbox_inst_37_T2 ;
    wire sbox_inst_37_T1 ;
    wire sbox_inst_37_T0 ;
    wire sbox_inst_36_n20 ;
    wire sbox_inst_36_n19 ;
    wire sbox_inst_36_n18 ;
    wire sbox_inst_36_n17 ;
    wire sbox_inst_36_n16 ;
    wire sbox_inst_36_n15 ;
    wire sbox_inst_36_n14 ;
    wire sbox_inst_36_n13 ;
    wire sbox_inst_36_n12 ;
    wire sbox_inst_36_n11 ;
    wire sbox_inst_36_T6 ;
    wire sbox_inst_36_L0 ;
    wire sbox_inst_36_T5 ;
    wire sbox_inst_36_T4 ;
    wire sbox_inst_36_T3 ;
    wire sbox_inst_36_T2 ;
    wire sbox_inst_36_T1 ;
    wire sbox_inst_36_T0 ;
    wire sbox_inst_35_n20 ;
    wire sbox_inst_35_n19 ;
    wire sbox_inst_35_n18 ;
    wire sbox_inst_35_n17 ;
    wire sbox_inst_35_n16 ;
    wire sbox_inst_35_n15 ;
    wire sbox_inst_35_n14 ;
    wire sbox_inst_35_n13 ;
    wire sbox_inst_35_n12 ;
    wire sbox_inst_35_n11 ;
    wire sbox_inst_35_T6 ;
    wire sbox_inst_35_L0 ;
    wire sbox_inst_35_T5 ;
    wire sbox_inst_35_T4 ;
    wire sbox_inst_35_T3 ;
    wire sbox_inst_35_T2 ;
    wire sbox_inst_35_T1 ;
    wire sbox_inst_35_T0 ;
    wire sbox_inst_34_n20 ;
    wire sbox_inst_34_n19 ;
    wire sbox_inst_34_n18 ;
    wire sbox_inst_34_n17 ;
    wire sbox_inst_34_n16 ;
    wire sbox_inst_34_n15 ;
    wire sbox_inst_34_n14 ;
    wire sbox_inst_34_n13 ;
    wire sbox_inst_34_n12 ;
    wire sbox_inst_34_n11 ;
    wire sbox_inst_34_T6 ;
    wire sbox_inst_34_L0 ;
    wire sbox_inst_34_T5 ;
    wire sbox_inst_34_T4 ;
    wire sbox_inst_34_T3 ;
    wire sbox_inst_34_T2 ;
    wire sbox_inst_34_T1 ;
    wire sbox_inst_34_T0 ;
    wire sbox_inst_33_n20 ;
    wire sbox_inst_33_n19 ;
    wire sbox_inst_33_n18 ;
    wire sbox_inst_33_n17 ;
    wire sbox_inst_33_n16 ;
    wire sbox_inst_33_n15 ;
    wire sbox_inst_33_n14 ;
    wire sbox_inst_33_n13 ;
    wire sbox_inst_33_n12 ;
    wire sbox_inst_33_n11 ;
    wire sbox_inst_33_T6 ;
    wire sbox_inst_33_L0 ;
    wire sbox_inst_33_T5 ;
    wire sbox_inst_33_T4 ;
    wire sbox_inst_33_T3 ;
    wire sbox_inst_33_T2 ;
    wire sbox_inst_33_T1 ;
    wire sbox_inst_33_T0 ;
    wire sbox_inst_32_n20 ;
    wire sbox_inst_32_n19 ;
    wire sbox_inst_32_n18 ;
    wire sbox_inst_32_n17 ;
    wire sbox_inst_32_n16 ;
    wire sbox_inst_32_n15 ;
    wire sbox_inst_32_n14 ;
    wire sbox_inst_32_n13 ;
    wire sbox_inst_32_n12 ;
    wire sbox_inst_32_n11 ;
    wire sbox_inst_32_T6 ;
    wire sbox_inst_32_L0 ;
    wire sbox_inst_32_T5 ;
    wire sbox_inst_32_T4 ;
    wire sbox_inst_32_T3 ;
    wire sbox_inst_32_T2 ;
    wire sbox_inst_32_T1 ;
    wire sbox_inst_32_T0 ;
    wire sbox_inst_31_n20 ;
    wire sbox_inst_31_n19 ;
    wire sbox_inst_31_n18 ;
    wire sbox_inst_31_n17 ;
    wire sbox_inst_31_n16 ;
    wire sbox_inst_31_n15 ;
    wire sbox_inst_31_n14 ;
    wire sbox_inst_31_n13 ;
    wire sbox_inst_31_n12 ;
    wire sbox_inst_31_n11 ;
    wire sbox_inst_31_T6 ;
    wire sbox_inst_31_L0 ;
    wire sbox_inst_31_T5 ;
    wire sbox_inst_31_T4 ;
    wire sbox_inst_31_T3 ;
    wire sbox_inst_31_T2 ;
    wire sbox_inst_31_T1 ;
    wire sbox_inst_31_T0 ;
    wire sbox_inst_30_n20 ;
    wire sbox_inst_30_n19 ;
    wire sbox_inst_30_n18 ;
    wire sbox_inst_30_n17 ;
    wire sbox_inst_30_n16 ;
    wire sbox_inst_30_n15 ;
    wire sbox_inst_30_n14 ;
    wire sbox_inst_30_n13 ;
    wire sbox_inst_30_n12 ;
    wire sbox_inst_30_n11 ;
    wire sbox_inst_30_T6 ;
    wire sbox_inst_30_L0 ;
    wire sbox_inst_30_T5 ;
    wire sbox_inst_30_T4 ;
    wire sbox_inst_30_T3 ;
    wire sbox_inst_30_T2 ;
    wire sbox_inst_30_T1 ;
    wire sbox_inst_30_T0 ;
    wire sbox_inst_29_n20 ;
    wire sbox_inst_29_n19 ;
    wire sbox_inst_29_n18 ;
    wire sbox_inst_29_n17 ;
    wire sbox_inst_29_n16 ;
    wire sbox_inst_29_n15 ;
    wire sbox_inst_29_n14 ;
    wire sbox_inst_29_n13 ;
    wire sbox_inst_29_n12 ;
    wire sbox_inst_29_n11 ;
    wire sbox_inst_29_T6 ;
    wire sbox_inst_29_L0 ;
    wire sbox_inst_29_T5 ;
    wire sbox_inst_29_T4 ;
    wire sbox_inst_29_T3 ;
    wire sbox_inst_29_T2 ;
    wire sbox_inst_29_T1 ;
    wire sbox_inst_29_T0 ;
    wire sbox_inst_28_n20 ;
    wire sbox_inst_28_n19 ;
    wire sbox_inst_28_n18 ;
    wire sbox_inst_28_n17 ;
    wire sbox_inst_28_n16 ;
    wire sbox_inst_28_n15 ;
    wire sbox_inst_28_n14 ;
    wire sbox_inst_28_n13 ;
    wire sbox_inst_28_n12 ;
    wire sbox_inst_28_n11 ;
    wire sbox_inst_28_T6 ;
    wire sbox_inst_28_L0 ;
    wire sbox_inst_28_T5 ;
    wire sbox_inst_28_T4 ;
    wire sbox_inst_28_T3 ;
    wire sbox_inst_28_T2 ;
    wire sbox_inst_28_T1 ;
    wire sbox_inst_28_T0 ;
    wire sbox_inst_27_n20 ;
    wire sbox_inst_27_n19 ;
    wire sbox_inst_27_n18 ;
    wire sbox_inst_27_n17 ;
    wire sbox_inst_27_n16 ;
    wire sbox_inst_27_n15 ;
    wire sbox_inst_27_n14 ;
    wire sbox_inst_27_n13 ;
    wire sbox_inst_27_n12 ;
    wire sbox_inst_27_n11 ;
    wire sbox_inst_27_T6 ;
    wire sbox_inst_27_L0 ;
    wire sbox_inst_27_T5 ;
    wire sbox_inst_27_T4 ;
    wire sbox_inst_27_T3 ;
    wire sbox_inst_27_T2 ;
    wire sbox_inst_27_T1 ;
    wire sbox_inst_27_T0 ;
    wire sbox_inst_26_n20 ;
    wire sbox_inst_26_n19 ;
    wire sbox_inst_26_n18 ;
    wire sbox_inst_26_n17 ;
    wire sbox_inst_26_n16 ;
    wire sbox_inst_26_n15 ;
    wire sbox_inst_26_n14 ;
    wire sbox_inst_26_n13 ;
    wire sbox_inst_26_n12 ;
    wire sbox_inst_26_n11 ;
    wire sbox_inst_26_T6 ;
    wire sbox_inst_26_L0 ;
    wire sbox_inst_26_T5 ;
    wire sbox_inst_26_T4 ;
    wire sbox_inst_26_T3 ;
    wire sbox_inst_26_T2 ;
    wire sbox_inst_26_T1 ;
    wire sbox_inst_26_T0 ;
    wire sbox_inst_25_n20 ;
    wire sbox_inst_25_n19 ;
    wire sbox_inst_25_n18 ;
    wire sbox_inst_25_n17 ;
    wire sbox_inst_25_n16 ;
    wire sbox_inst_25_n15 ;
    wire sbox_inst_25_n14 ;
    wire sbox_inst_25_n13 ;
    wire sbox_inst_25_n12 ;
    wire sbox_inst_25_n11 ;
    wire sbox_inst_25_T6 ;
    wire sbox_inst_25_L0 ;
    wire sbox_inst_25_T5 ;
    wire sbox_inst_25_T4 ;
    wire sbox_inst_25_T3 ;
    wire sbox_inst_25_T2 ;
    wire sbox_inst_25_T1 ;
    wire sbox_inst_25_T0 ;
    wire sbox_inst_24_n20 ;
    wire sbox_inst_24_n19 ;
    wire sbox_inst_24_n18 ;
    wire sbox_inst_24_n17 ;
    wire sbox_inst_24_n16 ;
    wire sbox_inst_24_n15 ;
    wire sbox_inst_24_n14 ;
    wire sbox_inst_24_n13 ;
    wire sbox_inst_24_n12 ;
    wire sbox_inst_24_n11 ;
    wire sbox_inst_24_T6 ;
    wire sbox_inst_24_L0 ;
    wire sbox_inst_24_T5 ;
    wire sbox_inst_24_T4 ;
    wire sbox_inst_24_T3 ;
    wire sbox_inst_24_T2 ;
    wire sbox_inst_24_T1 ;
    wire sbox_inst_24_T0 ;
    wire sbox_inst_23_n20 ;
    wire sbox_inst_23_n19 ;
    wire sbox_inst_23_n18 ;
    wire sbox_inst_23_n17 ;
    wire sbox_inst_23_n16 ;
    wire sbox_inst_23_n15 ;
    wire sbox_inst_23_n14 ;
    wire sbox_inst_23_n13 ;
    wire sbox_inst_23_n12 ;
    wire sbox_inst_23_n11 ;
    wire sbox_inst_23_T6 ;
    wire sbox_inst_23_L0 ;
    wire sbox_inst_23_T5 ;
    wire sbox_inst_23_T4 ;
    wire sbox_inst_23_T3 ;
    wire sbox_inst_23_T2 ;
    wire sbox_inst_23_T1 ;
    wire sbox_inst_23_T0 ;
    wire sbox_inst_22_n20 ;
    wire sbox_inst_22_n19 ;
    wire sbox_inst_22_n18 ;
    wire sbox_inst_22_n17 ;
    wire sbox_inst_22_n16 ;
    wire sbox_inst_22_n15 ;
    wire sbox_inst_22_n14 ;
    wire sbox_inst_22_n13 ;
    wire sbox_inst_22_n12 ;
    wire sbox_inst_22_n11 ;
    wire sbox_inst_22_T6 ;
    wire sbox_inst_22_L0 ;
    wire sbox_inst_22_T5 ;
    wire sbox_inst_22_T4 ;
    wire sbox_inst_22_T3 ;
    wire sbox_inst_22_T2 ;
    wire sbox_inst_22_T1 ;
    wire sbox_inst_22_T0 ;
    wire sbox_inst_21_n20 ;
    wire sbox_inst_21_n19 ;
    wire sbox_inst_21_n18 ;
    wire sbox_inst_21_n17 ;
    wire sbox_inst_21_n16 ;
    wire sbox_inst_21_n15 ;
    wire sbox_inst_21_n14 ;
    wire sbox_inst_21_n13 ;
    wire sbox_inst_21_n12 ;
    wire sbox_inst_21_n11 ;
    wire sbox_inst_21_T6 ;
    wire sbox_inst_21_L0 ;
    wire sbox_inst_21_T5 ;
    wire sbox_inst_21_T4 ;
    wire sbox_inst_21_T3 ;
    wire sbox_inst_21_T2 ;
    wire sbox_inst_21_T1 ;
    wire sbox_inst_21_T0 ;
    wire sbox_inst_20_n20 ;
    wire sbox_inst_20_n19 ;
    wire sbox_inst_20_n18 ;
    wire sbox_inst_20_n17 ;
    wire sbox_inst_20_n16 ;
    wire sbox_inst_20_n15 ;
    wire sbox_inst_20_n14 ;
    wire sbox_inst_20_n13 ;
    wire sbox_inst_20_n12 ;
    wire sbox_inst_20_n11 ;
    wire sbox_inst_20_T6 ;
    wire sbox_inst_20_L0 ;
    wire sbox_inst_20_T5 ;
    wire sbox_inst_20_T4 ;
    wire sbox_inst_20_T3 ;
    wire sbox_inst_20_T2 ;
    wire sbox_inst_20_T1 ;
    wire sbox_inst_20_T0 ;
    wire sbox_inst_19_n20 ;
    wire sbox_inst_19_n19 ;
    wire sbox_inst_19_n18 ;
    wire sbox_inst_19_n17 ;
    wire sbox_inst_19_n16 ;
    wire sbox_inst_19_n15 ;
    wire sbox_inst_19_n14 ;
    wire sbox_inst_19_n13 ;
    wire sbox_inst_19_n12 ;
    wire sbox_inst_19_n11 ;
    wire sbox_inst_19_T6 ;
    wire sbox_inst_19_L0 ;
    wire sbox_inst_19_T5 ;
    wire sbox_inst_19_T4 ;
    wire sbox_inst_19_T3 ;
    wire sbox_inst_19_T2 ;
    wire sbox_inst_19_T1 ;
    wire sbox_inst_19_T0 ;
    wire sbox_inst_18_n20 ;
    wire sbox_inst_18_n19 ;
    wire sbox_inst_18_n18 ;
    wire sbox_inst_18_n17 ;
    wire sbox_inst_18_n16 ;
    wire sbox_inst_18_n15 ;
    wire sbox_inst_18_n14 ;
    wire sbox_inst_18_n13 ;
    wire sbox_inst_18_n12 ;
    wire sbox_inst_18_n11 ;
    wire sbox_inst_18_T6 ;
    wire sbox_inst_18_L0 ;
    wire sbox_inst_18_T5 ;
    wire sbox_inst_18_T4 ;
    wire sbox_inst_18_T3 ;
    wire sbox_inst_18_T2 ;
    wire sbox_inst_18_T1 ;
    wire sbox_inst_18_T0 ;
    wire sbox_inst_17_n20 ;
    wire sbox_inst_17_n19 ;
    wire sbox_inst_17_n18 ;
    wire sbox_inst_17_n17 ;
    wire sbox_inst_17_n16 ;
    wire sbox_inst_17_n15 ;
    wire sbox_inst_17_n14 ;
    wire sbox_inst_17_n13 ;
    wire sbox_inst_17_n12 ;
    wire sbox_inst_17_n11 ;
    wire sbox_inst_17_T6 ;
    wire sbox_inst_17_L0 ;
    wire sbox_inst_17_T5 ;
    wire sbox_inst_17_T4 ;
    wire sbox_inst_17_T3 ;
    wire sbox_inst_17_T2 ;
    wire sbox_inst_17_T1 ;
    wire sbox_inst_17_T0 ;
    wire sbox_inst_16_n20 ;
    wire sbox_inst_16_n19 ;
    wire sbox_inst_16_n18 ;
    wire sbox_inst_16_n17 ;
    wire sbox_inst_16_n16 ;
    wire sbox_inst_16_n15 ;
    wire sbox_inst_16_n14 ;
    wire sbox_inst_16_n13 ;
    wire sbox_inst_16_n12 ;
    wire sbox_inst_16_n11 ;
    wire sbox_inst_16_T6 ;
    wire sbox_inst_16_L0 ;
    wire sbox_inst_16_T5 ;
    wire sbox_inst_16_T4 ;
    wire sbox_inst_16_T3 ;
    wire sbox_inst_16_T2 ;
    wire sbox_inst_16_T1 ;
    wire sbox_inst_16_T0 ;
    wire sbox_inst_15_n20 ;
    wire sbox_inst_15_n19 ;
    wire sbox_inst_15_n18 ;
    wire sbox_inst_15_n17 ;
    wire sbox_inst_15_n16 ;
    wire sbox_inst_15_n15 ;
    wire sbox_inst_15_n14 ;
    wire sbox_inst_15_n13 ;
    wire sbox_inst_15_n12 ;
    wire sbox_inst_15_n11 ;
    wire sbox_inst_15_T6 ;
    wire sbox_inst_15_L0 ;
    wire sbox_inst_15_T5 ;
    wire sbox_inst_15_T4 ;
    wire sbox_inst_15_T3 ;
    wire sbox_inst_15_T2 ;
    wire sbox_inst_15_T1 ;
    wire sbox_inst_15_T0 ;
    wire sbox_inst_14_n20 ;
    wire sbox_inst_14_n19 ;
    wire sbox_inst_14_n18 ;
    wire sbox_inst_14_n17 ;
    wire sbox_inst_14_n16 ;
    wire sbox_inst_14_n15 ;
    wire sbox_inst_14_n14 ;
    wire sbox_inst_14_n13 ;
    wire sbox_inst_14_n12 ;
    wire sbox_inst_14_n11 ;
    wire sbox_inst_14_T6 ;
    wire sbox_inst_14_L0 ;
    wire sbox_inst_14_T5 ;
    wire sbox_inst_14_T4 ;
    wire sbox_inst_14_T3 ;
    wire sbox_inst_14_T2 ;
    wire sbox_inst_14_T1 ;
    wire sbox_inst_14_T0 ;
    wire sbox_inst_13_n20 ;
    wire sbox_inst_13_n19 ;
    wire sbox_inst_13_n18 ;
    wire sbox_inst_13_n17 ;
    wire sbox_inst_13_n16 ;
    wire sbox_inst_13_n15 ;
    wire sbox_inst_13_n14 ;
    wire sbox_inst_13_n13 ;
    wire sbox_inst_13_n12 ;
    wire sbox_inst_13_n11 ;
    wire sbox_inst_13_T6 ;
    wire sbox_inst_13_L0 ;
    wire sbox_inst_13_T5 ;
    wire sbox_inst_13_T4 ;
    wire sbox_inst_13_T3 ;
    wire sbox_inst_13_T2 ;
    wire sbox_inst_13_T1 ;
    wire sbox_inst_13_T0 ;
    wire sbox_inst_12_n20 ;
    wire sbox_inst_12_n19 ;
    wire sbox_inst_12_n18 ;
    wire sbox_inst_12_n17 ;
    wire sbox_inst_12_n16 ;
    wire sbox_inst_12_n15 ;
    wire sbox_inst_12_n14 ;
    wire sbox_inst_12_n13 ;
    wire sbox_inst_12_n12 ;
    wire sbox_inst_12_n11 ;
    wire sbox_inst_12_T6 ;
    wire sbox_inst_12_L0 ;
    wire sbox_inst_12_T5 ;
    wire sbox_inst_12_T4 ;
    wire sbox_inst_12_T3 ;
    wire sbox_inst_12_T2 ;
    wire sbox_inst_12_T1 ;
    wire sbox_inst_12_T0 ;
    wire sbox_inst_11_n20 ;
    wire sbox_inst_11_n19 ;
    wire sbox_inst_11_n18 ;
    wire sbox_inst_11_n17 ;
    wire sbox_inst_11_n16 ;
    wire sbox_inst_11_n15 ;
    wire sbox_inst_11_n14 ;
    wire sbox_inst_11_n13 ;
    wire sbox_inst_11_n12 ;
    wire sbox_inst_11_n11 ;
    wire sbox_inst_11_T6 ;
    wire sbox_inst_11_L0 ;
    wire sbox_inst_11_T5 ;
    wire sbox_inst_11_T4 ;
    wire sbox_inst_11_T3 ;
    wire sbox_inst_11_T2 ;
    wire sbox_inst_11_T1 ;
    wire sbox_inst_11_T0 ;
    wire sbox_inst_10_n20 ;
    wire sbox_inst_10_n19 ;
    wire sbox_inst_10_n18 ;
    wire sbox_inst_10_n17 ;
    wire sbox_inst_10_n16 ;
    wire sbox_inst_10_n15 ;
    wire sbox_inst_10_n14 ;
    wire sbox_inst_10_n13 ;
    wire sbox_inst_10_n12 ;
    wire sbox_inst_10_n11 ;
    wire sbox_inst_10_T6 ;
    wire sbox_inst_10_L0 ;
    wire sbox_inst_10_T5 ;
    wire sbox_inst_10_T4 ;
    wire sbox_inst_10_T3 ;
    wire sbox_inst_10_T2 ;
    wire sbox_inst_10_T1 ;
    wire sbox_inst_10_T0 ;
    wire sbox_inst_9_n20 ;
    wire sbox_inst_9_n19 ;
    wire sbox_inst_9_n18 ;
    wire sbox_inst_9_n17 ;
    wire sbox_inst_9_n16 ;
    wire sbox_inst_9_n15 ;
    wire sbox_inst_9_n14 ;
    wire sbox_inst_9_n13 ;
    wire sbox_inst_9_n12 ;
    wire sbox_inst_9_n11 ;
    wire sbox_inst_9_T6 ;
    wire sbox_inst_9_L0 ;
    wire sbox_inst_9_T5 ;
    wire sbox_inst_9_T4 ;
    wire sbox_inst_9_T3 ;
    wire sbox_inst_9_T2 ;
    wire sbox_inst_9_T1 ;
    wire sbox_inst_9_T0 ;
    wire sbox_inst_8_n20 ;
    wire sbox_inst_8_n19 ;
    wire sbox_inst_8_n18 ;
    wire sbox_inst_8_n17 ;
    wire sbox_inst_8_n16 ;
    wire sbox_inst_8_n15 ;
    wire sbox_inst_8_n14 ;
    wire sbox_inst_8_n13 ;
    wire sbox_inst_8_n12 ;
    wire sbox_inst_8_n11 ;
    wire sbox_inst_8_T6 ;
    wire sbox_inst_8_L0 ;
    wire sbox_inst_8_T5 ;
    wire sbox_inst_8_T4 ;
    wire sbox_inst_8_T3 ;
    wire sbox_inst_8_T2 ;
    wire sbox_inst_8_T1 ;
    wire sbox_inst_8_T0 ;
    wire sbox_inst_7_n20 ;
    wire sbox_inst_7_n19 ;
    wire sbox_inst_7_n18 ;
    wire sbox_inst_7_n17 ;
    wire sbox_inst_7_n16 ;
    wire sbox_inst_7_n15 ;
    wire sbox_inst_7_n14 ;
    wire sbox_inst_7_n13 ;
    wire sbox_inst_7_n12 ;
    wire sbox_inst_7_n11 ;
    wire sbox_inst_7_T6 ;
    wire sbox_inst_7_L0 ;
    wire sbox_inst_7_T5 ;
    wire sbox_inst_7_T4 ;
    wire sbox_inst_7_T3 ;
    wire sbox_inst_7_T2 ;
    wire sbox_inst_7_T1 ;
    wire sbox_inst_7_T0 ;
    wire sbox_inst_6_n20 ;
    wire sbox_inst_6_n19 ;
    wire sbox_inst_6_n18 ;
    wire sbox_inst_6_n17 ;
    wire sbox_inst_6_n16 ;
    wire sbox_inst_6_n15 ;
    wire sbox_inst_6_n14 ;
    wire sbox_inst_6_n13 ;
    wire sbox_inst_6_n12 ;
    wire sbox_inst_6_n11 ;
    wire sbox_inst_6_T6 ;
    wire sbox_inst_6_L0 ;
    wire sbox_inst_6_T5 ;
    wire sbox_inst_6_T4 ;
    wire sbox_inst_6_T3 ;
    wire sbox_inst_6_T2 ;
    wire sbox_inst_6_T1 ;
    wire sbox_inst_6_T0 ;
    wire sbox_inst_5_n20 ;
    wire sbox_inst_5_n19 ;
    wire sbox_inst_5_n18 ;
    wire sbox_inst_5_n17 ;
    wire sbox_inst_5_n16 ;
    wire sbox_inst_5_n15 ;
    wire sbox_inst_5_n14 ;
    wire sbox_inst_5_n13 ;
    wire sbox_inst_5_n12 ;
    wire sbox_inst_5_n11 ;
    wire sbox_inst_5_T6 ;
    wire sbox_inst_5_L0 ;
    wire sbox_inst_5_T5 ;
    wire sbox_inst_5_T4 ;
    wire sbox_inst_5_T3 ;
    wire sbox_inst_5_T2 ;
    wire sbox_inst_5_T1 ;
    wire sbox_inst_5_T0 ;
    wire sbox_inst_4_n20 ;
    wire sbox_inst_4_n19 ;
    wire sbox_inst_4_n18 ;
    wire sbox_inst_4_n17 ;
    wire sbox_inst_4_n16 ;
    wire sbox_inst_4_n15 ;
    wire sbox_inst_4_n14 ;
    wire sbox_inst_4_n13 ;
    wire sbox_inst_4_n12 ;
    wire sbox_inst_4_n11 ;
    wire sbox_inst_4_T6 ;
    wire sbox_inst_4_L0 ;
    wire sbox_inst_4_T5 ;
    wire sbox_inst_4_T4 ;
    wire sbox_inst_4_T3 ;
    wire sbox_inst_4_T2 ;
    wire sbox_inst_4_T1 ;
    wire sbox_inst_4_T0 ;
    wire sbox_inst_3_n20 ;
    wire sbox_inst_3_n19 ;
    wire sbox_inst_3_n18 ;
    wire sbox_inst_3_n17 ;
    wire sbox_inst_3_n16 ;
    wire sbox_inst_3_n15 ;
    wire sbox_inst_3_n14 ;
    wire sbox_inst_3_n13 ;
    wire sbox_inst_3_n12 ;
    wire sbox_inst_3_n11 ;
    wire sbox_inst_3_T6 ;
    wire sbox_inst_3_L0 ;
    wire sbox_inst_3_T5 ;
    wire sbox_inst_3_T4 ;
    wire sbox_inst_3_T3 ;
    wire sbox_inst_3_T2 ;
    wire sbox_inst_3_T1 ;
    wire sbox_inst_3_T0 ;
    wire sbox_inst_2_n20 ;
    wire sbox_inst_2_n19 ;
    wire sbox_inst_2_n18 ;
    wire sbox_inst_2_n17 ;
    wire sbox_inst_2_n16 ;
    wire sbox_inst_2_n15 ;
    wire sbox_inst_2_n14 ;
    wire sbox_inst_2_n13 ;
    wire sbox_inst_2_n12 ;
    wire sbox_inst_2_n11 ;
    wire sbox_inst_2_T6 ;
    wire sbox_inst_2_L0 ;
    wire sbox_inst_2_T5 ;
    wire sbox_inst_2_T4 ;
    wire sbox_inst_2_T3 ;
    wire sbox_inst_2_T2 ;
    wire sbox_inst_2_T1 ;
    wire sbox_inst_2_T0 ;
    wire sbox_inst_1_n20 ;
    wire sbox_inst_1_n19 ;
    wire sbox_inst_1_n18 ;
    wire sbox_inst_1_n17 ;
    wire sbox_inst_1_n16 ;
    wire sbox_inst_1_n15 ;
    wire sbox_inst_1_n14 ;
    wire sbox_inst_1_n13 ;
    wire sbox_inst_1_n12 ;
    wire sbox_inst_1_n11 ;
    wire sbox_inst_1_T6 ;
    wire sbox_inst_1_L0 ;
    wire sbox_inst_1_T5 ;
    wire sbox_inst_1_T4 ;
    wire sbox_inst_1_T3 ;
    wire sbox_inst_1_T2 ;
    wire sbox_inst_1_T1 ;
    wire sbox_inst_1_T0 ;
    wire sbox_inst_0_n20 ;
    wire sbox_inst_0_n19 ;
    wire sbox_inst_0_n18 ;
    wire sbox_inst_0_n17 ;
    wire sbox_inst_0_n16 ;
    wire sbox_inst_0_n15 ;
    wire sbox_inst_0_n14 ;
    wire sbox_inst_0_n13 ;
    wire sbox_inst_0_n12 ;
    wire sbox_inst_0_n11 ;
    wire sbox_inst_0_T6 ;
    wire sbox_inst_0_L0 ;
    wire sbox_inst_0_T5 ;
    wire sbox_inst_0_T4 ;
    wire sbox_inst_0_T3 ;
    wire sbox_inst_0_T2 ;
    wire sbox_inst_0_T1 ;
    wire sbox_inst_0_T0 ;
    wire [159:153] input_array ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    //wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) U29 ( .a ({input0_s2[1], input0_s1[1], input0_s0[1]}), .b ({1'b0, 1'b0, lfsr[1]}), .c ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, input_array_1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U30 ( .a ({input0_s2[157], input0_s1[157], input0_s0[157]}), .b ({1'b0, 1'b0, rev_lfsr[4]}), .c ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, input_array[157]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U31 ( .a ({input0_s2[153], input0_s1[153], input0_s0[153]}), .b ({1'b0, 1'b0, rev_lfsr[0]}), .c ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, input_array[153]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U32 ( .a ({input0_s2[5], input0_s1[5], input0_s0[5]}), .b ({1'b0, 1'b0, lfsr[5]}), .c ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, input_array_5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U33 ( .a ({input0_s2[6], input0_s1[6], input0_s0[6]}), .b ({1'b0, 1'b0, lfsr[6]}), .c ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, input_array_6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U34 ( .a ({input0_s2[4], input0_s1[4], input0_s0[4]}), .b ({1'b0, 1'b0, lfsr[4]}), .c ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, input_array_4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U35 ( .a ({input0_s2[3], input0_s1[3], input0_s0[3]}), .b ({1'b0, 1'b0, lfsr[3]}), .c ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, input_array_3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U36 ( .a ({input0_s2[2], input0_s1[2], input0_s0[2]}), .b ({1'b0, 1'b0, lfsr[2]}), .c ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, input_array_2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U37 ( .a ({input0_s2[0], input0_s1[0], input0_s0[0]}), .b ({1'b0, 1'b0, lfsr[0]}), .c ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, input_array_0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U38 ( .a ({input0_s2[159], input0_s1[159], input0_s0[159]}), .b ({1'b0, 1'b0, rev_lfsr[6]}), .c ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, input_array[159]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U39 ( .a ({input0_s2[158], input0_s1[158], input0_s0[158]}), .b ({1'b0, 1'b0, rev_lfsr[5]}), .c ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, input_array[158]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U40 ( .a ({input0_s2[156], input0_s1[156], input0_s0[156]}), .b ({1'b0, 1'b0, rev_lfsr[3]}), .c ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, input_array[156]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U41 ( .a ({input0_s2[155], input0_s1[155], input0_s0[155]}), .b ({1'b0, 1'b0, rev_lfsr[2]}), .c ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, input_array[155]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U42 ( .a ({input0_s2[154], input0_s1[154], input0_s0[154]}), .b ({1'b0, 1'b0, rev_lfsr[1]}), .c ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, input_array[154]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U1 ( .a ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, input_array[158]}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, input_array[157]}), .c ({new_AGEMA_signal_1852, new_AGEMA_signal_1851, sbox_inst_39_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U1 ( .a ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, input_array[154]}), .b ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, input_array[153]}), .c ({new_AGEMA_signal_1864, new_AGEMA_signal_1863, sbox_inst_38_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U1 ( .a ({input0_s2[150], input0_s1[150], input0_s0[150]}), .b ({input0_s2[149], input0_s1[149], input0_s0[149]}), .c ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, sbox_inst_37_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U1 ( .a ({input0_s2[146], input0_s1[146], input0_s0[146]}), .b ({input0_s2[145], input0_s1[145], input0_s0[145]}), .c ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, sbox_inst_36_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U1 ( .a ({input0_s2[142], input0_s1[142], input0_s0[142]}), .b ({input0_s2[141], input0_s1[141], input0_s0[141]}), .c ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, sbox_inst_35_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U1 ( .a ({input0_s2[138], input0_s1[138], input0_s0[138]}), .b ({input0_s2[137], input0_s1[137], input0_s0[137]}), .c ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, sbox_inst_34_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U1 ( .a ({input0_s2[134], input0_s1[134], input0_s0[134]}), .b ({input0_s2[133], input0_s1[133], input0_s0[133]}), .c ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, sbox_inst_33_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U1 ( .a ({input0_s2[130], input0_s1[130], input0_s0[130]}), .b ({input0_s2[129], input0_s1[129], input0_s0[129]}), .c ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, sbox_inst_32_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U1 ( .a ({input0_s2[126], input0_s1[126], input0_s0[126]}), .b ({input0_s2[125], input0_s1[125], input0_s0[125]}), .c ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, sbox_inst_31_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U1 ( .a ({input0_s2[122], input0_s1[122], input0_s0[122]}), .b ({input0_s2[121], input0_s1[121], input0_s0[121]}), .c ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, sbox_inst_30_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U1 ( .a ({input0_s2[118], input0_s1[118], input0_s0[118]}), .b ({input0_s2[117], input0_s1[117], input0_s0[117]}), .c ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, sbox_inst_29_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U1 ( .a ({input0_s2[114], input0_s1[114], input0_s0[114]}), .b ({input0_s2[113], input0_s1[113], input0_s0[113]}), .c ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, sbox_inst_28_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U1 ( .a ({input0_s2[110], input0_s1[110], input0_s0[110]}), .b ({input0_s2[109], input0_s1[109], input0_s0[109]}), .c ({new_AGEMA_signal_1336, new_AGEMA_signal_1335, sbox_inst_27_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U1 ( .a ({input0_s2[106], input0_s1[106], input0_s0[106]}), .b ({input0_s2[105], input0_s1[105], input0_s0[105]}), .c ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, sbox_inst_26_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U1 ( .a ({input0_s2[102], input0_s1[102], input0_s0[102]}), .b ({input0_s2[101], input0_s1[101], input0_s0[101]}), .c ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, sbox_inst_25_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U1 ( .a ({input0_s2[98], input0_s1[98], input0_s0[98]}), .b ({input0_s2[97], input0_s1[97], input0_s0[97]}), .c ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, sbox_inst_24_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U1 ( .a ({input0_s2[94], input0_s1[94], input0_s0[94]}), .b ({input0_s2[93], input0_s1[93], input0_s0[93]}), .c ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, sbox_inst_23_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U1 ( .a ({input0_s2[90], input0_s1[90], input0_s0[90]}), .b ({input0_s2[89], input0_s1[89], input0_s0[89]}), .c ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, sbox_inst_22_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U1 ( .a ({input0_s2[86], input0_s1[86], input0_s0[86]}), .b ({input0_s2[85], input0_s1[85], input0_s0[85]}), .c ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, sbox_inst_21_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U1 ( .a ({input0_s2[82], input0_s1[82], input0_s0[82]}), .b ({input0_s2[81], input0_s1[81], input0_s0[81]}), .c ({new_AGEMA_signal_1476, new_AGEMA_signal_1475, sbox_inst_20_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U1 ( .a ({input0_s2[78], input0_s1[78], input0_s0[78]}), .b ({input0_s2[77], input0_s1[77], input0_s0[77]}), .c ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, sbox_inst_19_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U1 ( .a ({input0_s2[74], input0_s1[74], input0_s0[74]}), .b ({input0_s2[73], input0_s1[73], input0_s0[73]}), .c ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, sbox_inst_18_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U1 ( .a ({input0_s2[70], input0_s1[70], input0_s0[70]}), .b ({input0_s2[69], input0_s1[69], input0_s0[69]}), .c ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, sbox_inst_17_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U1 ( .a ({input0_s2[66], input0_s1[66], input0_s0[66]}), .b ({input0_s2[65], input0_s1[65], input0_s0[65]}), .c ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, sbox_inst_16_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U1 ( .a ({input0_s2[62], input0_s1[62], input0_s0[62]}), .b ({input0_s2[61], input0_s1[61], input0_s0[61]}), .c ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, sbox_inst_15_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U1 ( .a ({input0_s2[58], input0_s1[58], input0_s0[58]}), .b ({input0_s2[57], input0_s1[57], input0_s0[57]}), .c ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, sbox_inst_14_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U1 ( .a ({input0_s2[54], input0_s1[54], input0_s0[54]}), .b ({input0_s2[53], input0_s1[53], input0_s0[53]}), .c ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, sbox_inst_13_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U1 ( .a ({input0_s2[50], input0_s1[50], input0_s0[50]}), .b ({input0_s2[49], input0_s1[49], input0_s0[49]}), .c ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, sbox_inst_12_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U1 ( .a ({input0_s2[46], input0_s1[46], input0_s0[46]}), .b ({input0_s2[45], input0_s1[45], input0_s0[45]}), .c ({new_AGEMA_signal_1656, new_AGEMA_signal_1655, sbox_inst_11_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U1 ( .a ({input0_s2[42], input0_s1[42], input0_s0[42]}), .b ({input0_s2[41], input0_s1[41], input0_s0[41]}), .c ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, sbox_inst_10_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U1 ( .a ({input0_s2[38], input0_s1[38], input0_s0[38]}), .b ({input0_s2[37], input0_s1[37], input0_s0[37]}), .c ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, sbox_inst_9_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U1 ( .a ({input0_s2[34], input0_s1[34], input0_s0[34]}), .b ({input0_s2[33], input0_s1[33], input0_s0[33]}), .c ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, sbox_inst_8_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U1 ( .a ({input0_s2[30], input0_s1[30], input0_s0[30]}), .b ({input0_s2[29], input0_s1[29], input0_s0[29]}), .c ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, sbox_inst_7_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U1 ( .a ({input0_s2[26], input0_s1[26], input0_s0[26]}), .b ({input0_s2[25], input0_s1[25], input0_s0[25]}), .c ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, sbox_inst_6_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U1 ( .a ({input0_s2[22], input0_s1[22], input0_s0[22]}), .b ({input0_s2[21], input0_s1[21], input0_s0[21]}), .c ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, sbox_inst_5_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U1 ( .a ({input0_s2[18], input0_s1[18], input0_s0[18]}), .b ({input0_s2[17], input0_s1[17], input0_s0[17]}), .c ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, sbox_inst_4_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U1 ( .a ({input0_s2[14], input0_s1[14], input0_s0[14]}), .b ({input0_s2[13], input0_s1[13], input0_s0[13]}), .c ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, sbox_inst_3_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U1 ( .a ({input0_s2[10], input0_s1[10], input0_s0[10]}), .b ({input0_s2[9], input0_s1[9], input0_s0[9]}), .c ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, sbox_inst_2_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U1 ( .a ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, input_array_6}), .b ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, input_array_5}), .c ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, sbox_inst_1_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U1 ( .a ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, input_array_2}), .b ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, input_array_1}), .c ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, sbox_inst_0_L0}) ) ;
    //ClockGatingController #(4) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U12 ( .a ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, sbox_inst_39_T3}), .b ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, sbox_inst_39_n17}), .c ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, sbox_inst_39_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U6 ( .a ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, sbox_inst_39_T4}), .b ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, sbox_inst_39_T2}), .c ({new_AGEMA_signal_2264, new_AGEMA_signal_2263, sbox_inst_39_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U5 ( .a ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, sbox_inst_39_T1}), .b ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, input_array[158]}), .c ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, sbox_inst_39_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U4 ( .a ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, sbox_inst_39_n11}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, input_array[157]}), .c ({output0_s2[39], output0_s1[39], output0_s0[39]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U3 ( .a ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, input_array[159]}), .b ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, sbox_inst_39_n17}), .c ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, sbox_inst_39_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U2 ( .a ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, input_array[156]}), .b ({new_AGEMA_signal_1854, new_AGEMA_signal_1853, sbox_inst_39_T0}), .c ({new_AGEMA_signal_2268, new_AGEMA_signal_2267, sbox_inst_39_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_t0_AND_U1 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, input_array[157]}), .b ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, input_array[158]}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1854, new_AGEMA_signal_1853, sbox_inst_39_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_t1_AND_U1 ( .a ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, input_array[156]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, input_array[159]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, sbox_inst_39_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_t2_AND_U1 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, input_array[157]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, input_array[159]}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, sbox_inst_39_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_t3_AND_U1 ( .a ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, input_array[158]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, input_array[159]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, sbox_inst_39_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_t4_AND_U1 ( .a ({new_AGEMA_signal_1122, new_AGEMA_signal_1121, input_array[156]}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, input_array[157]}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, sbox_inst_39_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U12 ( .a ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, sbox_inst_38_T3}), .b ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, sbox_inst_38_n17}), .c ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, sbox_inst_38_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U6 ( .a ({new_AGEMA_signal_1876, new_AGEMA_signal_1875, sbox_inst_38_T4}), .b ({new_AGEMA_signal_1872, new_AGEMA_signal_1871, sbox_inst_38_T2}), .c ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, sbox_inst_38_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U5 ( .a ({new_AGEMA_signal_1870, new_AGEMA_signal_1869, sbox_inst_38_T1}), .b ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, input_array[154]}), .c ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, sbox_inst_38_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U4 ( .a ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, sbox_inst_38_n11}), .b ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, input_array[153]}), .c ({output0_s2[38], output0_s1[38], output0_s0[38]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U3 ( .a ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, input_array[155]}), .b ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, sbox_inst_38_n17}), .c ({new_AGEMA_signal_2682, new_AGEMA_signal_2681, sbox_inst_38_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U2 ( .a ({input0_s2[152], input0_s1[152], input0_s0[152]}), .b ({new_AGEMA_signal_1866, new_AGEMA_signal_1865, sbox_inst_38_T0}), .c ({new_AGEMA_signal_2278, new_AGEMA_signal_2277, sbox_inst_38_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_t0_AND_U1 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, input_array[153]}), .b ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, input_array[154]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_1866, new_AGEMA_signal_1865, sbox_inst_38_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_t1_AND_U1 ( .a ({input0_s2[152], input0_s1[152], input0_s0[152]}), .b ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, input_array[155]}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1870, new_AGEMA_signal_1869, sbox_inst_38_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_t2_AND_U1 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, input_array[153]}), .b ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, input_array[155]}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_1872, new_AGEMA_signal_1871, sbox_inst_38_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_t3_AND_U1 ( .a ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, input_array[154]}), .b ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, input_array[155]}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, sbox_inst_38_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_t4_AND_U1 ( .a ({input0_s2[152], input0_s1[152], input0_s0[152]}), .b ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, input_array[153]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_1876, new_AGEMA_signal_1875, sbox_inst_38_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U12 ( .a ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, sbox_inst_37_T3}), .b ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, sbox_inst_37_n17}), .c ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, sbox_inst_37_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U6 ( .a ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, sbox_inst_37_T4}), .b ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, sbox_inst_37_T2}), .c ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, sbox_inst_37_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U5 ( .a ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, sbox_inst_37_T1}), .b ({input0_s2[150], input0_s1[150], input0_s0[150]}), .c ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, sbox_inst_37_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U4 ( .a ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, sbox_inst_37_n11}), .b ({input0_s2[149], input0_s1[149], input0_s0[149]}), .c ({output0_s2[37], output0_s1[37], output0_s0[37]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U3 ( .a ({input0_s2[151], input0_s1[151], input0_s0[151]}), .b ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, sbox_inst_37_n17}), .c ({new_AGEMA_signal_2292, new_AGEMA_signal_2291, sbox_inst_37_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U2 ( .a ({input0_s2[148], input0_s1[148], input0_s0[148]}), .b ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, sbox_inst_37_T0}), .c ({new_AGEMA_signal_1882, new_AGEMA_signal_1881, sbox_inst_37_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_t0_AND_U1 ( .a ({input0_s2[149], input0_s1[149], input0_s0[149]}), .b ({input0_s2[150], input0_s1[150], input0_s0[150]}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, sbox_inst_37_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_t1_AND_U1 ( .a ({input0_s2[148], input0_s1[148], input0_s0[148]}), .b ({input0_s2[151], input0_s1[151], input0_s0[151]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, sbox_inst_37_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_t2_AND_U1 ( .a ({input0_s2[149], input0_s1[149], input0_s0[149]}), .b ({input0_s2[151], input0_s1[151], input0_s0[151]}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, sbox_inst_37_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_t3_AND_U1 ( .a ({input0_s2[150], input0_s1[150], input0_s0[150]}), .b ({input0_s2[151], input0_s1[151], input0_s0[151]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, sbox_inst_37_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_t4_AND_U1 ( .a ({input0_s2[148], input0_s1[148], input0_s0[148]}), .b ({input0_s2[149], input0_s1[149], input0_s0[149]}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1150, new_AGEMA_signal_1149, sbox_inst_37_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U12 ( .a ({new_AGEMA_signal_1168, new_AGEMA_signal_1167, sbox_inst_36_T3}), .b ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, sbox_inst_36_n17}), .c ({new_AGEMA_signal_2296, new_AGEMA_signal_2295, sbox_inst_36_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U6 ( .a ({new_AGEMA_signal_1170, new_AGEMA_signal_1169, sbox_inst_36_T4}), .b ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, sbox_inst_36_T2}), .c ({new_AGEMA_signal_1888, new_AGEMA_signal_1887, sbox_inst_36_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U5 ( .a ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, sbox_inst_36_T1}), .b ({input0_s2[146], input0_s1[146], input0_s0[146]}), .c ({new_AGEMA_signal_1890, new_AGEMA_signal_1889, sbox_inst_36_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U4 ( .a ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, sbox_inst_36_n11}), .b ({input0_s2[145], input0_s1[145], input0_s0[145]}), .c ({output0_s2[36], output0_s1[36], output0_s0[36]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U3 ( .a ({input0_s2[147], input0_s1[147], input0_s0[147]}), .b ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, sbox_inst_36_n17}), .c ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, sbox_inst_36_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U2 ( .a ({input0_s2[144], input0_s1[144], input0_s0[144]}), .b ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, sbox_inst_36_T0}), .c ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, sbox_inst_36_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_t0_AND_U1 ( .a ({input0_s2[145], input0_s1[145], input0_s0[145]}), .b ({input0_s2[146], input0_s1[146], input0_s0[146]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_1158, new_AGEMA_signal_1157, sbox_inst_36_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_t1_AND_U1 ( .a ({input0_s2[144], input0_s1[144], input0_s0[144]}), .b ({input0_s2[147], input0_s1[147], input0_s0[147]}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, sbox_inst_36_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_t2_AND_U1 ( .a ({input0_s2[145], input0_s1[145], input0_s0[145]}), .b ({input0_s2[147], input0_s1[147], input0_s0[147]}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, sbox_inst_36_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_t3_AND_U1 ( .a ({input0_s2[146], input0_s1[146], input0_s0[146]}), .b ({input0_s2[147], input0_s1[147], input0_s0[147]}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1168, new_AGEMA_signal_1167, sbox_inst_36_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_t4_AND_U1 ( .a ({input0_s2[144], input0_s1[144], input0_s0[144]}), .b ({input0_s2[145], input0_s1[145], input0_s0[145]}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_1170, new_AGEMA_signal_1169, sbox_inst_36_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U12 ( .a ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, sbox_inst_35_T3}), .b ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, sbox_inst_35_n17}), .c ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, sbox_inst_35_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U6 ( .a ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, sbox_inst_35_T4}), .b ({new_AGEMA_signal_1186, new_AGEMA_signal_1185, sbox_inst_35_T2}), .c ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, sbox_inst_35_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U5 ( .a ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, sbox_inst_35_T1}), .b ({input0_s2[142], input0_s1[142], input0_s0[142]}), .c ({new_AGEMA_signal_1900, new_AGEMA_signal_1899, sbox_inst_35_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U4 ( .a ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, sbox_inst_35_n11}), .b ({input0_s2[141], input0_s1[141], input0_s0[141]}), .c ({output0_s2[35], output0_s1[35], output0_s0[35]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U3 ( .a ({input0_s2[143], input0_s1[143], input0_s0[143]}), .b ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, sbox_inst_35_n17}), .c ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, sbox_inst_35_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U2 ( .a ({input0_s2[140], input0_s1[140], input0_s0[140]}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, sbox_inst_35_T0}), .c ({new_AGEMA_signal_1902, new_AGEMA_signal_1901, sbox_inst_35_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_t0_AND_U1 ( .a ({input0_s2[141], input0_s1[141], input0_s0[141]}), .b ({input0_s2[142], input0_s1[142], input0_s0[142]}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, sbox_inst_35_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_t1_AND_U1 ( .a ({input0_s2[140], input0_s1[140], input0_s0[140]}), .b ({input0_s2[143], input0_s1[143], input0_s0[143]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, sbox_inst_35_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_t2_AND_U1 ( .a ({input0_s2[141], input0_s1[141], input0_s0[141]}), .b ({input0_s2[143], input0_s1[143], input0_s0[143]}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1186, new_AGEMA_signal_1185, sbox_inst_35_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_t3_AND_U1 ( .a ({input0_s2[142], input0_s1[142], input0_s0[142]}), .b ({input0_s2[143], input0_s1[143], input0_s0[143]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, sbox_inst_35_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_t4_AND_U1 ( .a ({input0_s2[140], input0_s1[140], input0_s0[140]}), .b ({input0_s2[141], input0_s1[141], input0_s0[141]}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, sbox_inst_35_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U12 ( .a ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, sbox_inst_34_T3}), .b ({new_AGEMA_signal_1912, new_AGEMA_signal_1911, sbox_inst_34_n17}), .c ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, sbox_inst_34_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U6 ( .a ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, sbox_inst_34_T4}), .b ({new_AGEMA_signal_1206, new_AGEMA_signal_1205, sbox_inst_34_T2}), .c ({new_AGEMA_signal_1908, new_AGEMA_signal_1907, sbox_inst_34_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U5 ( .a ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, sbox_inst_34_T1}), .b ({input0_s2[138], input0_s1[138], input0_s0[138]}), .c ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, sbox_inst_34_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U4 ( .a ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, sbox_inst_34_n11}), .b ({input0_s2[137], input0_s1[137], input0_s0[137]}), .c ({output0_s2[34], output0_s1[34], output0_s0[34]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U3 ( .a ({input0_s2[139], input0_s1[139], input0_s0[139]}), .b ({new_AGEMA_signal_1912, new_AGEMA_signal_1911, sbox_inst_34_n17}), .c ({new_AGEMA_signal_2322, new_AGEMA_signal_2321, sbox_inst_34_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U2 ( .a ({input0_s2[136], input0_s1[136], input0_s0[136]}), .b ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, sbox_inst_34_T0}), .c ({new_AGEMA_signal_1912, new_AGEMA_signal_1911, sbox_inst_34_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_t0_AND_U1 ( .a ({input0_s2[137], input0_s1[137], input0_s0[137]}), .b ({input0_s2[138], input0_s1[138], input0_s0[138]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_1198, new_AGEMA_signal_1197, sbox_inst_34_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_t1_AND_U1 ( .a ({input0_s2[136], input0_s1[136], input0_s0[136]}), .b ({input0_s2[139], input0_s1[139], input0_s0[139]}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, sbox_inst_34_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_t2_AND_U1 ( .a ({input0_s2[137], input0_s1[137], input0_s0[137]}), .b ({input0_s2[139], input0_s1[139], input0_s0[139]}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_1206, new_AGEMA_signal_1205, sbox_inst_34_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_t3_AND_U1 ( .a ({input0_s2[138], input0_s1[138], input0_s0[138]}), .b ({input0_s2[139], input0_s1[139], input0_s0[139]}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, sbox_inst_34_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_t4_AND_U1 ( .a ({input0_s2[136], input0_s1[136], input0_s0[136]}), .b ({input0_s2[137], input0_s1[137], input0_s0[137]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, sbox_inst_34_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U12 ( .a ({new_AGEMA_signal_1228, new_AGEMA_signal_1227, sbox_inst_33_T3}), .b ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, sbox_inst_33_n17}), .c ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, sbox_inst_33_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U6 ( .a ({new_AGEMA_signal_1230, new_AGEMA_signal_1229, sbox_inst_33_T4}), .b ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, sbox_inst_33_T2}), .c ({new_AGEMA_signal_1918, new_AGEMA_signal_1917, sbox_inst_33_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U5 ( .a ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, sbox_inst_33_T1}), .b ({input0_s2[134], input0_s1[134], input0_s0[134]}), .c ({new_AGEMA_signal_1920, new_AGEMA_signal_1919, sbox_inst_33_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U4 ( .a ({new_AGEMA_signal_2332, new_AGEMA_signal_2331, sbox_inst_33_n11}), .b ({input0_s2[133], input0_s1[133], input0_s0[133]}), .c ({output0_s2[33], output0_s1[33], output0_s0[33]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U3 ( .a ({input0_s2[135], input0_s1[135], input0_s0[135]}), .b ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, sbox_inst_33_n17}), .c ({new_AGEMA_signal_2332, new_AGEMA_signal_2331, sbox_inst_33_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U2 ( .a ({input0_s2[132], input0_s1[132], input0_s0[132]}), .b ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, sbox_inst_33_T0}), .c ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, sbox_inst_33_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_t0_AND_U1 ( .a ({input0_s2[133], input0_s1[133], input0_s0[133]}), .b ({input0_s2[134], input0_s1[134], input0_s0[134]}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1218, new_AGEMA_signal_1217, sbox_inst_33_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_t1_AND_U1 ( .a ({input0_s2[132], input0_s1[132], input0_s0[132]}), .b ({input0_s2[135], input0_s1[135], input0_s0[135]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, sbox_inst_33_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_t2_AND_U1 ( .a ({input0_s2[133], input0_s1[133], input0_s0[133]}), .b ({input0_s2[135], input0_s1[135], input0_s0[135]}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, sbox_inst_33_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_t3_AND_U1 ( .a ({input0_s2[134], input0_s1[134], input0_s0[134]}), .b ({input0_s2[135], input0_s1[135], input0_s0[135]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_1228, new_AGEMA_signal_1227, sbox_inst_33_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_t4_AND_U1 ( .a ({input0_s2[132], input0_s1[132], input0_s0[132]}), .b ({input0_s2[133], input0_s1[133], input0_s0[133]}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1230, new_AGEMA_signal_1229, sbox_inst_33_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U12 ( .a ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, sbox_inst_32_T3}), .b ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, sbox_inst_32_n17}), .c ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, sbox_inst_32_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U6 ( .a ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, sbox_inst_32_T4}), .b ({new_AGEMA_signal_1246, new_AGEMA_signal_1245, sbox_inst_32_T2}), .c ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, sbox_inst_32_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U5 ( .a ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, sbox_inst_32_T1}), .b ({input0_s2[130], input0_s1[130], input0_s0[130]}), .c ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, sbox_inst_32_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U4 ( .a ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, sbox_inst_32_n11}), .b ({input0_s2[129], input0_s1[129], input0_s0[129]}), .c ({output0_s2[32], output0_s1[32], output0_s0[32]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U3 ( .a ({input0_s2[131], input0_s1[131], input0_s0[131]}), .b ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, sbox_inst_32_n17}), .c ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, sbox_inst_32_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U2 ( .a ({input0_s2[128], input0_s1[128], input0_s0[128]}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, sbox_inst_32_T0}), .c ({new_AGEMA_signal_1932, new_AGEMA_signal_1931, sbox_inst_32_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_t0_AND_U1 ( .a ({input0_s2[129], input0_s1[129], input0_s0[129]}), .b ({input0_s2[130], input0_s1[130], input0_s0[130]}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, sbox_inst_32_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_t1_AND_U1 ( .a ({input0_s2[128], input0_s1[128], input0_s0[128]}), .b ({input0_s2[131], input0_s1[131], input0_s0[131]}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, sbox_inst_32_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_t2_AND_U1 ( .a ({input0_s2[129], input0_s1[129], input0_s0[129]}), .b ({input0_s2[131], input0_s1[131], input0_s0[131]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_1246, new_AGEMA_signal_1245, sbox_inst_32_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_t3_AND_U1 ( .a ({input0_s2[130], input0_s1[130], input0_s0[130]}), .b ({input0_s2[131], input0_s1[131], input0_s0[131]}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, sbox_inst_32_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_t4_AND_U1 ( .a ({input0_s2[128], input0_s1[128], input0_s0[128]}), .b ({input0_s2[129], input0_s1[129], input0_s0[129]}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, sbox_inst_32_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U12 ( .a ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, sbox_inst_31_T3}), .b ({new_AGEMA_signal_1942, new_AGEMA_signal_1941, sbox_inst_31_n17}), .c ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, sbox_inst_31_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U6 ( .a ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, sbox_inst_31_T4}), .b ({new_AGEMA_signal_1266, new_AGEMA_signal_1265, sbox_inst_31_T2}), .c ({new_AGEMA_signal_1938, new_AGEMA_signal_1937, sbox_inst_31_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U5 ( .a ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, sbox_inst_31_T1}), .b ({input0_s2[126], input0_s1[126], input0_s0[126]}), .c ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, sbox_inst_31_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U4 ( .a ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, sbox_inst_31_n11}), .b ({input0_s2[125], input0_s1[125], input0_s0[125]}), .c ({output0_s2[31], output0_s1[31], output0_s0[31]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U3 ( .a ({input0_s2[127], input0_s1[127], input0_s0[127]}), .b ({new_AGEMA_signal_1942, new_AGEMA_signal_1941, sbox_inst_31_n17}), .c ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, sbox_inst_31_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U2 ( .a ({input0_s2[124], input0_s1[124], input0_s0[124]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, sbox_inst_31_T0}), .c ({new_AGEMA_signal_1942, new_AGEMA_signal_1941, sbox_inst_31_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_t0_AND_U1 ( .a ({input0_s2[125], input0_s1[125], input0_s0[125]}), .b ({input0_s2[126], input0_s1[126], input0_s0[126]}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, sbox_inst_31_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_t1_AND_U1 ( .a ({input0_s2[124], input0_s1[124], input0_s0[124]}), .b ({input0_s2[127], input0_s1[127], input0_s0[127]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, sbox_inst_31_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_t2_AND_U1 ( .a ({input0_s2[125], input0_s1[125], input0_s0[125]}), .b ({input0_s2[127], input0_s1[127], input0_s0[127]}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1266, new_AGEMA_signal_1265, sbox_inst_31_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_t3_AND_U1 ( .a ({input0_s2[126], input0_s1[126], input0_s0[126]}), .b ({input0_s2[127], input0_s1[127], input0_s0[127]}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, sbox_inst_31_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_t4_AND_U1 ( .a ({input0_s2[124], input0_s1[124], input0_s0[124]}), .b ({input0_s2[125], input0_s1[125], input0_s0[125]}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1270, new_AGEMA_signal_1269, sbox_inst_31_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U12 ( .a ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, sbox_inst_30_T3}), .b ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, sbox_inst_30_n17}), .c ({new_AGEMA_signal_2356, new_AGEMA_signal_2355, sbox_inst_30_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U6 ( .a ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, sbox_inst_30_T4}), .b ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, sbox_inst_30_T2}), .c ({new_AGEMA_signal_1948, new_AGEMA_signal_1947, sbox_inst_30_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U5 ( .a ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, sbox_inst_30_T1}), .b ({input0_s2[122], input0_s1[122], input0_s0[122]}), .c ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, sbox_inst_30_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U4 ( .a ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, sbox_inst_30_n11}), .b ({input0_s2[121], input0_s1[121], input0_s0[121]}), .c ({output0_s2[30], output0_s1[30], output0_s0[30]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U3 ( .a ({input0_s2[123], input0_s1[123], input0_s0[123]}), .b ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, sbox_inst_30_n17}), .c ({new_AGEMA_signal_2362, new_AGEMA_signal_2361, sbox_inst_30_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U2 ( .a ({input0_s2[120], input0_s1[120], input0_s0[120]}), .b ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, sbox_inst_30_T0}), .c ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, sbox_inst_30_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_t0_AND_U1 ( .a ({input0_s2[121], input0_s1[121], input0_s0[121]}), .b ({input0_s2[122], input0_s1[122], input0_s0[122]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_1278, new_AGEMA_signal_1277, sbox_inst_30_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_t1_AND_U1 ( .a ({input0_s2[120], input0_s1[120], input0_s0[120]}), .b ({input0_s2[123], input0_s1[123], input0_s0[123]}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, sbox_inst_30_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_t2_AND_U1 ( .a ({input0_s2[121], input0_s1[121], input0_s0[121]}), .b ({input0_s2[123], input0_s1[123], input0_s0[123]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, sbox_inst_30_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_t3_AND_U1 ( .a ({input0_s2[122], input0_s1[122], input0_s0[122]}), .b ({input0_s2[123], input0_s1[123], input0_s0[123]}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, sbox_inst_30_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_t4_AND_U1 ( .a ({input0_s2[120], input0_s1[120], input0_s0[120]}), .b ({input0_s2[121], input0_s1[121], input0_s0[121]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_1290, new_AGEMA_signal_1289, sbox_inst_30_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U12 ( .a ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, sbox_inst_29_T3}), .b ({new_AGEMA_signal_1962, new_AGEMA_signal_1961, sbox_inst_29_n17}), .c ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, sbox_inst_29_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U6 ( .a ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, sbox_inst_29_T4}), .b ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, sbox_inst_29_T2}), .c ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, sbox_inst_29_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U5 ( .a ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, sbox_inst_29_T1}), .b ({input0_s2[118], input0_s1[118], input0_s0[118]}), .c ({new_AGEMA_signal_1960, new_AGEMA_signal_1959, sbox_inst_29_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U4 ( .a ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, sbox_inst_29_n11}), .b ({input0_s2[117], input0_s1[117], input0_s0[117]}), .c ({output0_s2[29], output0_s1[29], output0_s0[29]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U3 ( .a ({input0_s2[119], input0_s1[119], input0_s0[119]}), .b ({new_AGEMA_signal_1962, new_AGEMA_signal_1961, sbox_inst_29_n17}), .c ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, sbox_inst_29_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U2 ( .a ({input0_s2[116], input0_s1[116], input0_s0[116]}), .b ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, sbox_inst_29_T0}), .c ({new_AGEMA_signal_1962, new_AGEMA_signal_1961, sbox_inst_29_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_t0_AND_U1 ( .a ({input0_s2[117], input0_s1[117], input0_s0[117]}), .b ({input0_s2[118], input0_s1[118], input0_s0[118]}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, sbox_inst_29_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_t1_AND_U1 ( .a ({input0_s2[116], input0_s1[116], input0_s0[116]}), .b ({input0_s2[119], input0_s1[119], input0_s0[119]}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, sbox_inst_29_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_t2_AND_U1 ( .a ({input0_s2[117], input0_s1[117], input0_s0[117]}), .b ({input0_s2[119], input0_s1[119], input0_s0[119]}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, sbox_inst_29_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_t3_AND_U1 ( .a ({input0_s2[118], input0_s1[118], input0_s0[118]}), .b ({input0_s2[119], input0_s1[119], input0_s0[119]}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, sbox_inst_29_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_t4_AND_U1 ( .a ({input0_s2[116], input0_s1[116], input0_s0[116]}), .b ({input0_s2[117], input0_s1[117], input0_s0[117]}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, sbox_inst_29_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U12 ( .a ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, sbox_inst_28_T3}), .b ({new_AGEMA_signal_1972, new_AGEMA_signal_1971, sbox_inst_28_n17}), .c ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, sbox_inst_28_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U6 ( .a ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, sbox_inst_28_T4}), .b ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, sbox_inst_28_T2}), .c ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, sbox_inst_28_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U5 ( .a ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, sbox_inst_28_T1}), .b ({input0_s2[114], input0_s1[114], input0_s0[114]}), .c ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, sbox_inst_28_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U4 ( .a ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, sbox_inst_28_n11}), .b ({input0_s2[113], input0_s1[113], input0_s0[113]}), .c ({output0_s2[28], output0_s1[28], output0_s0[28]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U3 ( .a ({input0_s2[115], input0_s1[115], input0_s0[115]}), .b ({new_AGEMA_signal_1972, new_AGEMA_signal_1971, sbox_inst_28_n17}), .c ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, sbox_inst_28_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U2 ( .a ({input0_s2[112], input0_s1[112], input0_s0[112]}), .b ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, sbox_inst_28_T0}), .c ({new_AGEMA_signal_1972, new_AGEMA_signal_1971, sbox_inst_28_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_t0_AND_U1 ( .a ({input0_s2[113], input0_s1[113], input0_s0[113]}), .b ({input0_s2[114], input0_s1[114], input0_s0[114]}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_1318, new_AGEMA_signal_1317, sbox_inst_28_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_t1_AND_U1 ( .a ({input0_s2[112], input0_s1[112], input0_s0[112]}), .b ({input0_s2[115], input0_s1[115], input0_s0[115]}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, sbox_inst_28_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_t2_AND_U1 ( .a ({input0_s2[113], input0_s1[113], input0_s0[113]}), .b ({input0_s2[115], input0_s1[115], input0_s0[115]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, sbox_inst_28_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_t3_AND_U1 ( .a ({input0_s2[114], input0_s1[114], input0_s0[114]}), .b ({input0_s2[115], input0_s1[115], input0_s0[115]}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, sbox_inst_28_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_t4_AND_U1 ( .a ({input0_s2[112], input0_s1[112], input0_s0[112]}), .b ({input0_s2[113], input0_s1[113], input0_s0[113]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, sbox_inst_28_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U12 ( .a ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, sbox_inst_27_T3}), .b ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, sbox_inst_27_n17}), .c ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, sbox_inst_27_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U6 ( .a ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, sbox_inst_27_T4}), .b ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, sbox_inst_27_T2}), .c ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, sbox_inst_27_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U5 ( .a ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, sbox_inst_27_T1}), .b ({input0_s2[110], input0_s1[110], input0_s0[110]}), .c ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, sbox_inst_27_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U4 ( .a ({new_AGEMA_signal_2392, new_AGEMA_signal_2391, sbox_inst_27_n11}), .b ({input0_s2[109], input0_s1[109], input0_s0[109]}), .c ({output0_s2[27], output0_s1[27], output0_s0[27]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U3 ( .a ({input0_s2[111], input0_s1[111], input0_s0[111]}), .b ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, sbox_inst_27_n17}), .c ({new_AGEMA_signal_2392, new_AGEMA_signal_2391, sbox_inst_27_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U2 ( .a ({input0_s2[108], input0_s1[108], input0_s0[108]}), .b ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, sbox_inst_27_T0}), .c ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, sbox_inst_27_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_t0_AND_U1 ( .a ({input0_s2[109], input0_s1[109], input0_s0[109]}), .b ({input0_s2[110], input0_s1[110], input0_s0[110]}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1338, new_AGEMA_signal_1337, sbox_inst_27_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_t1_AND_U1 ( .a ({input0_s2[108], input0_s1[108], input0_s0[108]}), .b ({input0_s2[111], input0_s1[111], input0_s0[111]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, sbox_inst_27_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_t2_AND_U1 ( .a ({input0_s2[109], input0_s1[109], input0_s0[109]}), .b ({input0_s2[111], input0_s1[111], input0_s0[111]}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, sbox_inst_27_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_t3_AND_U1 ( .a ({input0_s2[110], input0_s1[110], input0_s0[110]}), .b ({input0_s2[111], input0_s1[111], input0_s0[111]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, sbox_inst_27_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_t4_AND_U1 ( .a ({input0_s2[108], input0_s1[108], input0_s0[108]}), .b ({input0_s2[109], input0_s1[109], input0_s0[109]}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1350, new_AGEMA_signal_1349, sbox_inst_27_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U12 ( .a ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, sbox_inst_26_T3}), .b ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, sbox_inst_26_n17}), .c ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, sbox_inst_26_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U6 ( .a ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, sbox_inst_26_T4}), .b ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, sbox_inst_26_T2}), .c ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, sbox_inst_26_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U5 ( .a ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, sbox_inst_26_T1}), .b ({input0_s2[106], input0_s1[106], input0_s0[106]}), .c ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, sbox_inst_26_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U4 ( .a ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, sbox_inst_26_n11}), .b ({input0_s2[105], input0_s1[105], input0_s0[105]}), .c ({output0_s2[26], output0_s1[26], output0_s0[26]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U3 ( .a ({input0_s2[107], input0_s1[107], input0_s0[107]}), .b ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, sbox_inst_26_n17}), .c ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, sbox_inst_26_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U2 ( .a ({input0_s2[104], input0_s1[104], input0_s0[104]}), .b ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, sbox_inst_26_T0}), .c ({new_AGEMA_signal_1992, new_AGEMA_signal_1991, sbox_inst_26_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_t0_AND_U1 ( .a ({input0_s2[105], input0_s1[105], input0_s0[105]}), .b ({input0_s2[106], input0_s1[106], input0_s0[106]}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, sbox_inst_26_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_t1_AND_U1 ( .a ({input0_s2[104], input0_s1[104], input0_s0[104]}), .b ({input0_s2[107], input0_s1[107], input0_s0[107]}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, sbox_inst_26_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_t2_AND_U1 ( .a ({input0_s2[105], input0_s1[105], input0_s0[105]}), .b ({input0_s2[107], input0_s1[107], input0_s0[107]}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, sbox_inst_26_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_t3_AND_U1 ( .a ({input0_s2[106], input0_s1[106], input0_s0[106]}), .b ({input0_s2[107], input0_s1[107], input0_s0[107]}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, sbox_inst_26_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_t4_AND_U1 ( .a ({input0_s2[104], input0_s1[104], input0_s0[104]}), .b ({input0_s2[105], input0_s1[105], input0_s0[105]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, sbox_inst_26_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U12 ( .a ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, sbox_inst_25_T3}), .b ({new_AGEMA_signal_2002, new_AGEMA_signal_2001, sbox_inst_25_n17}), .c ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, sbox_inst_25_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U6 ( .a ({new_AGEMA_signal_1390, new_AGEMA_signal_1389, sbox_inst_25_T4}), .b ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, sbox_inst_25_T2}), .c ({new_AGEMA_signal_1998, new_AGEMA_signal_1997, sbox_inst_25_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U5 ( .a ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, sbox_inst_25_T1}), .b ({input0_s2[102], input0_s1[102], input0_s0[102]}), .c ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, sbox_inst_25_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U4 ( .a ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, sbox_inst_25_n11}), .b ({input0_s2[101], input0_s1[101], input0_s0[101]}), .c ({output0_s2[25], output0_s1[25], output0_s0[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U3 ( .a ({input0_s2[103], input0_s1[103], input0_s0[103]}), .b ({new_AGEMA_signal_2002, new_AGEMA_signal_2001, sbox_inst_25_n17}), .c ({new_AGEMA_signal_2412, new_AGEMA_signal_2411, sbox_inst_25_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U2 ( .a ({input0_s2[100], input0_s1[100], input0_s0[100]}), .b ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, sbox_inst_25_T0}), .c ({new_AGEMA_signal_2002, new_AGEMA_signal_2001, sbox_inst_25_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_t0_AND_U1 ( .a ({input0_s2[101], input0_s1[101], input0_s0[101]}), .b ({input0_s2[102], input0_s1[102], input0_s0[102]}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, sbox_inst_25_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_t1_AND_U1 ( .a ({input0_s2[100], input0_s1[100], input0_s0[100]}), .b ({input0_s2[103], input0_s1[103], input0_s0[103]}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, sbox_inst_25_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_t2_AND_U1 ( .a ({input0_s2[101], input0_s1[101], input0_s0[101]}), .b ({input0_s2[103], input0_s1[103], input0_s0[103]}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, sbox_inst_25_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_t3_AND_U1 ( .a ({input0_s2[102], input0_s1[102], input0_s0[102]}), .b ({input0_s2[103], input0_s1[103], input0_s0[103]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, sbox_inst_25_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_t4_AND_U1 ( .a ({input0_s2[100], input0_s1[100], input0_s0[100]}), .b ({input0_s2[101], input0_s1[101], input0_s0[101]}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1390, new_AGEMA_signal_1389, sbox_inst_25_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U12 ( .a ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, sbox_inst_24_T3}), .b ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, sbox_inst_24_n17}), .c ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, sbox_inst_24_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U6 ( .a ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, sbox_inst_24_T4}), .b ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, sbox_inst_24_T2}), .c ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, sbox_inst_24_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U5 ( .a ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, sbox_inst_24_T1}), .b ({input0_s2[98], input0_s1[98], input0_s0[98]}), .c ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, sbox_inst_24_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U4 ( .a ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, sbox_inst_24_n11}), .b ({input0_s2[97], input0_s1[97], input0_s0[97]}), .c ({output0_s2[24], output0_s1[24], output0_s0[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U3 ( .a ({input0_s2[99], input0_s1[99], input0_s0[99]}), .b ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, sbox_inst_24_n17}), .c ({new_AGEMA_signal_2422, new_AGEMA_signal_2421, sbox_inst_24_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U2 ( .a ({input0_s2[96], input0_s1[96], input0_s0[96]}), .b ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, sbox_inst_24_T0}), .c ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, sbox_inst_24_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_t0_AND_U1 ( .a ({input0_s2[97], input0_s1[97], input0_s0[97]}), .b ({input0_s2[98], input0_s1[98], input0_s0[98]}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_1398, new_AGEMA_signal_1397, sbox_inst_24_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_t1_AND_U1 ( .a ({input0_s2[96], input0_s1[96], input0_s0[96]}), .b ({input0_s2[99], input0_s1[99], input0_s0[99]}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, sbox_inst_24_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_t2_AND_U1 ( .a ({input0_s2[97], input0_s1[97], input0_s0[97]}), .b ({input0_s2[99], input0_s1[99], input0_s0[99]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, sbox_inst_24_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_t3_AND_U1 ( .a ({input0_s2[98], input0_s1[98], input0_s0[98]}), .b ({input0_s2[99], input0_s1[99], input0_s0[99]}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, sbox_inst_24_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_t4_AND_U1 ( .a ({input0_s2[96], input0_s1[96], input0_s0[96]}), .b ({input0_s2[97], input0_s1[97], input0_s0[97]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_1410, new_AGEMA_signal_1409, sbox_inst_24_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U12 ( .a ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, sbox_inst_23_T3}), .b ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, sbox_inst_23_n17}), .c ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, sbox_inst_23_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U6 ( .a ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, sbox_inst_23_T4}), .b ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, sbox_inst_23_T2}), .c ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, sbox_inst_23_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U5 ( .a ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, sbox_inst_23_T1}), .b ({input0_s2[94], input0_s1[94], input0_s0[94]}), .c ({new_AGEMA_signal_2020, new_AGEMA_signal_2019, sbox_inst_23_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U4 ( .a ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, sbox_inst_23_n11}), .b ({input0_s2[93], input0_s1[93], input0_s0[93]}), .c ({output0_s2[23], output0_s1[23], output0_s0[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U3 ( .a ({input0_s2[95], input0_s1[95], input0_s0[95]}), .b ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, sbox_inst_23_n17}), .c ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, sbox_inst_23_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U2 ( .a ({input0_s2[92], input0_s1[92], input0_s0[92]}), .b ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, sbox_inst_23_T0}), .c ({new_AGEMA_signal_2022, new_AGEMA_signal_2021, sbox_inst_23_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_t0_AND_U1 ( .a ({input0_s2[93], input0_s1[93], input0_s0[93]}), .b ({input0_s2[94], input0_s1[94], input0_s0[94]}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, sbox_inst_23_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_t1_AND_U1 ( .a ({input0_s2[92], input0_s1[92], input0_s0[92]}), .b ({input0_s2[95], input0_s1[95], input0_s0[95]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, sbox_inst_23_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_t2_AND_U1 ( .a ({input0_s2[93], input0_s1[93], input0_s0[93]}), .b ({input0_s2[95], input0_s1[95], input0_s0[95]}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, sbox_inst_23_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_t3_AND_U1 ( .a ({input0_s2[94], input0_s1[94], input0_s0[94]}), .b ({input0_s2[95], input0_s1[95], input0_s0[95]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, sbox_inst_23_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_t4_AND_U1 ( .a ({input0_s2[92], input0_s1[92], input0_s0[92]}), .b ({input0_s2[93], input0_s1[93], input0_s0[93]}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, sbox_inst_23_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U12 ( .a ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, sbox_inst_22_T3}), .b ({new_AGEMA_signal_2032, new_AGEMA_signal_2031, sbox_inst_22_n17}), .c ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, sbox_inst_22_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U6 ( .a ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, sbox_inst_22_T4}), .b ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, sbox_inst_22_T2}), .c ({new_AGEMA_signal_2028, new_AGEMA_signal_2027, sbox_inst_22_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U5 ( .a ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, sbox_inst_22_T1}), .b ({input0_s2[90], input0_s1[90], input0_s0[90]}), .c ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, sbox_inst_22_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U4 ( .a ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, sbox_inst_22_n11}), .b ({input0_s2[89], input0_s1[89], input0_s0[89]}), .c ({output0_s2[22], output0_s1[22], output0_s0[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U3 ( .a ({input0_s2[91], input0_s1[91], input0_s0[91]}), .b ({new_AGEMA_signal_2032, new_AGEMA_signal_2031, sbox_inst_22_n17}), .c ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, sbox_inst_22_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U2 ( .a ({input0_s2[88], input0_s1[88], input0_s0[88]}), .b ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, sbox_inst_22_T0}), .c ({new_AGEMA_signal_2032, new_AGEMA_signal_2031, sbox_inst_22_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_t0_AND_U1 ( .a ({input0_s2[89], input0_s1[89], input0_s0[89]}), .b ({input0_s2[90], input0_s1[90], input0_s0[90]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, sbox_inst_22_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_t1_AND_U1 ( .a ({input0_s2[88], input0_s1[88], input0_s0[88]}), .b ({input0_s2[91], input0_s1[91], input0_s0[91]}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, sbox_inst_22_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_t2_AND_U1 ( .a ({input0_s2[89], input0_s1[89], input0_s0[89]}), .b ({input0_s2[91], input0_s1[91], input0_s0[91]}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, sbox_inst_22_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_t3_AND_U1 ( .a ({input0_s2[90], input0_s1[90], input0_s0[90]}), .b ({input0_s2[91], input0_s1[91], input0_s0[91]}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, sbox_inst_22_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_t4_AND_U1 ( .a ({input0_s2[88], input0_s1[88], input0_s0[88]}), .b ({input0_s2[89], input0_s1[89], input0_s0[89]}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, sbox_inst_22_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U12 ( .a ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, sbox_inst_21_T3}), .b ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, sbox_inst_21_n17}), .c ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, sbox_inst_21_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U6 ( .a ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, sbox_inst_21_T4}), .b ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, sbox_inst_21_T2}), .c ({new_AGEMA_signal_2038, new_AGEMA_signal_2037, sbox_inst_21_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U5 ( .a ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, sbox_inst_21_T1}), .b ({input0_s2[86], input0_s1[86], input0_s0[86]}), .c ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, sbox_inst_21_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U4 ( .a ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, sbox_inst_21_n11}), .b ({input0_s2[85], input0_s1[85], input0_s0[85]}), .c ({output0_s2[21], output0_s1[21], output0_s0[21]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U3 ( .a ({input0_s2[87], input0_s1[87], input0_s0[87]}), .b ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, sbox_inst_21_n17}), .c ({new_AGEMA_signal_2452, new_AGEMA_signal_2451, sbox_inst_21_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U2 ( .a ({input0_s2[84], input0_s1[84], input0_s0[84]}), .b ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, sbox_inst_21_T0}), .c ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, sbox_inst_21_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_t0_AND_U1 ( .a ({input0_s2[85], input0_s1[85], input0_s0[85]}), .b ({input0_s2[86], input0_s1[86], input0_s0[86]}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1458, new_AGEMA_signal_1457, sbox_inst_21_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_t1_AND_U1 ( .a ({input0_s2[84], input0_s1[84], input0_s0[84]}), .b ({input0_s2[87], input0_s1[87], input0_s0[87]}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, sbox_inst_21_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_t2_AND_U1 ( .a ({input0_s2[85], input0_s1[85], input0_s0[85]}), .b ({input0_s2[87], input0_s1[87], input0_s0[87]}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, sbox_inst_21_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_t3_AND_U1 ( .a ({input0_s2[86], input0_s1[86], input0_s0[86]}), .b ({input0_s2[87], input0_s1[87], input0_s0[87]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, sbox_inst_21_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_t4_AND_U1 ( .a ({input0_s2[84], input0_s1[84], input0_s0[84]}), .b ({input0_s2[85], input0_s1[85], input0_s0[85]}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1470, new_AGEMA_signal_1469, sbox_inst_21_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U12 ( .a ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, sbox_inst_20_T3}), .b ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, sbox_inst_20_n17}), .c ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, sbox_inst_20_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U6 ( .a ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, sbox_inst_20_T4}), .b ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, sbox_inst_20_T2}), .c ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, sbox_inst_20_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U5 ( .a ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, sbox_inst_20_T1}), .b ({input0_s2[82], input0_s1[82], input0_s0[82]}), .c ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, sbox_inst_20_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U4 ( .a ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, sbox_inst_20_n11}), .b ({input0_s2[81], input0_s1[81], input0_s0[81]}), .c ({output0_s2[20], output0_s1[20], output0_s0[20]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U3 ( .a ({input0_s2[83], input0_s1[83], input0_s0[83]}), .b ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, sbox_inst_20_n17}), .c ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, sbox_inst_20_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U2 ( .a ({input0_s2[80], input0_s1[80], input0_s0[80]}), .b ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, sbox_inst_20_T0}), .c ({new_AGEMA_signal_2052, new_AGEMA_signal_2051, sbox_inst_20_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_t0_AND_U1 ( .a ({input0_s2[81], input0_s1[81], input0_s0[81]}), .b ({input0_s2[82], input0_s1[82], input0_s0[82]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, sbox_inst_20_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_t1_AND_U1 ( .a ({input0_s2[80], input0_s1[80], input0_s0[80]}), .b ({input0_s2[83], input0_s1[83], input0_s0[83]}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, sbox_inst_20_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_t2_AND_U1 ( .a ({input0_s2[81], input0_s1[81], input0_s0[81]}), .b ({input0_s2[83], input0_s1[83], input0_s0[83]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, sbox_inst_20_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_t3_AND_U1 ( .a ({input0_s2[82], input0_s1[82], input0_s0[82]}), .b ({input0_s2[83], input0_s1[83], input0_s0[83]}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, sbox_inst_20_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_t4_AND_U1 ( .a ({input0_s2[80], input0_s1[80], input0_s0[80]}), .b ({input0_s2[81], input0_s1[81], input0_s0[81]}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, sbox_inst_20_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U12 ( .a ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, sbox_inst_19_T3}), .b ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, sbox_inst_19_n17}), .c ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, sbox_inst_19_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U6 ( .a ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, sbox_inst_19_T4}), .b ({new_AGEMA_signal_1506, new_AGEMA_signal_1505, sbox_inst_19_T2}), .c ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, sbox_inst_19_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U5 ( .a ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, sbox_inst_19_T1}), .b ({input0_s2[78], input0_s1[78], input0_s0[78]}), .c ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, sbox_inst_19_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U4 ( .a ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, sbox_inst_19_n11}), .b ({input0_s2[77], input0_s1[77], input0_s0[77]}), .c ({output0_s2[19], output0_s1[19], output0_s0[19]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U3 ( .a ({input0_s2[79], input0_s1[79], input0_s0[79]}), .b ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, sbox_inst_19_n17}), .c ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, sbox_inst_19_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U2 ( .a ({input0_s2[76], input0_s1[76], input0_s0[76]}), .b ({new_AGEMA_signal_1498, new_AGEMA_signal_1497, sbox_inst_19_T0}), .c ({new_AGEMA_signal_2062, new_AGEMA_signal_2061, sbox_inst_19_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_t0_AND_U1 ( .a ({input0_s2[77], input0_s1[77], input0_s0[77]}), .b ({input0_s2[78], input0_s1[78], input0_s0[78]}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1498, new_AGEMA_signal_1497, sbox_inst_19_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_t1_AND_U1 ( .a ({input0_s2[76], input0_s1[76], input0_s0[76]}), .b ({input0_s2[79], input0_s1[79], input0_s0[79]}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, sbox_inst_19_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_t2_AND_U1 ( .a ({input0_s2[77], input0_s1[77], input0_s0[77]}), .b ({input0_s2[79], input0_s1[79], input0_s0[79]}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1506, new_AGEMA_signal_1505, sbox_inst_19_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_t3_AND_U1 ( .a ({input0_s2[78], input0_s1[78], input0_s0[78]}), .b ({input0_s2[79], input0_s1[79], input0_s0[79]}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, sbox_inst_19_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_t4_AND_U1 ( .a ({input0_s2[76], input0_s1[76], input0_s0[76]}), .b ({input0_s2[77], input0_s1[77], input0_s0[77]}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, sbox_inst_19_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U12 ( .a ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, sbox_inst_18_T3}), .b ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, sbox_inst_18_n17}), .c ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, sbox_inst_18_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U6 ( .a ({new_AGEMA_signal_1530, new_AGEMA_signal_1529, sbox_inst_18_T4}), .b ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, sbox_inst_18_T2}), .c ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, sbox_inst_18_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U5 ( .a ({new_AGEMA_signal_1524, new_AGEMA_signal_1523, sbox_inst_18_T1}), .b ({input0_s2[74], input0_s1[74], input0_s0[74]}), .c ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, sbox_inst_18_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U4 ( .a ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, sbox_inst_18_n11}), .b ({input0_s2[73], input0_s1[73], input0_s0[73]}), .c ({output0_s2[18], output0_s1[18], output0_s0[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U3 ( .a ({input0_s2[75], input0_s1[75], input0_s0[75]}), .b ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, sbox_inst_18_n17}), .c ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, sbox_inst_18_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U2 ( .a ({input0_s2[72], input0_s1[72], input0_s0[72]}), .b ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, sbox_inst_18_T0}), .c ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, sbox_inst_18_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_t0_AND_U1 ( .a ({input0_s2[73], input0_s1[73], input0_s0[73]}), .b ({input0_s2[74], input0_s1[74], input0_s0[74]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_1518, new_AGEMA_signal_1517, sbox_inst_18_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_t1_AND_U1 ( .a ({input0_s2[72], input0_s1[72], input0_s0[72]}), .b ({input0_s2[75], input0_s1[75], input0_s0[75]}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1524, new_AGEMA_signal_1523, sbox_inst_18_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_t2_AND_U1 ( .a ({input0_s2[73], input0_s1[73], input0_s0[73]}), .b ({input0_s2[75], input0_s1[75], input0_s0[75]}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, sbox_inst_18_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_t3_AND_U1 ( .a ({input0_s2[74], input0_s1[74], input0_s0[74]}), .b ({input0_s2[75], input0_s1[75], input0_s0[75]}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, sbox_inst_18_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_t4_AND_U1 ( .a ({input0_s2[72], input0_s1[72], input0_s0[72]}), .b ({input0_s2[73], input0_s1[73], input0_s0[73]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_1530, new_AGEMA_signal_1529, sbox_inst_18_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U12 ( .a ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, sbox_inst_17_T3}), .b ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, sbox_inst_17_n17}), .c ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, sbox_inst_17_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U6 ( .a ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, sbox_inst_17_T4}), .b ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, sbox_inst_17_T2}), .c ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, sbox_inst_17_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U5 ( .a ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, sbox_inst_17_T1}), .b ({input0_s2[70], input0_s1[70], input0_s0[70]}), .c ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, sbox_inst_17_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U4 ( .a ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, sbox_inst_17_n11}), .b ({input0_s2[69], input0_s1[69], input0_s0[69]}), .c ({output0_s2[17], output0_s1[17], output0_s0[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U3 ( .a ({input0_s2[71], input0_s1[71], input0_s0[71]}), .b ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, sbox_inst_17_n17}), .c ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, sbox_inst_17_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U2 ( .a ({input0_s2[68], input0_s1[68], input0_s0[68]}), .b ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, sbox_inst_17_T0}), .c ({new_AGEMA_signal_2082, new_AGEMA_signal_2081, sbox_inst_17_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_t0_AND_U1 ( .a ({input0_s2[69], input0_s1[69], input0_s0[69]}), .b ({input0_s2[70], input0_s1[70], input0_s0[70]}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, sbox_inst_17_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_t1_AND_U1 ( .a ({input0_s2[68], input0_s1[68], input0_s0[68]}), .b ({input0_s2[71], input0_s1[71], input0_s0[71]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, sbox_inst_17_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_t2_AND_U1 ( .a ({input0_s2[69], input0_s1[69], input0_s0[69]}), .b ({input0_s2[71], input0_s1[71], input0_s0[71]}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, sbox_inst_17_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_t3_AND_U1 ( .a ({input0_s2[70], input0_s1[70], input0_s0[70]}), .b ({input0_s2[71], input0_s1[71], input0_s0[71]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, sbox_inst_17_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_t4_AND_U1 ( .a ({input0_s2[68], input0_s1[68], input0_s0[68]}), .b ({input0_s2[69], input0_s1[69], input0_s0[69]}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, sbox_inst_17_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U12 ( .a ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, sbox_inst_16_T3}), .b ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, sbox_inst_16_n17}), .c ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, sbox_inst_16_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U6 ( .a ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, sbox_inst_16_T4}), .b ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, sbox_inst_16_T2}), .c ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, sbox_inst_16_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U5 ( .a ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, sbox_inst_16_T1}), .b ({input0_s2[66], input0_s1[66], input0_s0[66]}), .c ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, sbox_inst_16_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U4 ( .a ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, sbox_inst_16_n11}), .b ({input0_s2[65], input0_s1[65], input0_s0[65]}), .c ({output0_s2[16], output0_s1[16], output0_s0[16]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U3 ( .a ({input0_s2[67], input0_s1[67], input0_s0[67]}), .b ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, sbox_inst_16_n17}), .c ({new_AGEMA_signal_2502, new_AGEMA_signal_2501, sbox_inst_16_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U2 ( .a ({input0_s2[64], input0_s1[64], input0_s0[64]}), .b ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, sbox_inst_16_T0}), .c ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, sbox_inst_16_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_t0_AND_U1 ( .a ({input0_s2[65], input0_s1[65], input0_s0[65]}), .b ({input0_s2[66], input0_s1[66], input0_s0[66]}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, sbox_inst_16_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_t1_AND_U1 ( .a ({input0_s2[64], input0_s1[64], input0_s0[64]}), .b ({input0_s2[67], input0_s1[67], input0_s0[67]}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, sbox_inst_16_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_t2_AND_U1 ( .a ({input0_s2[65], input0_s1[65], input0_s0[65]}), .b ({input0_s2[67], input0_s1[67], input0_s0[67]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, sbox_inst_16_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_t3_AND_U1 ( .a ({input0_s2[66], input0_s1[66], input0_s0[66]}), .b ({input0_s2[67], input0_s1[67], input0_s0[67]}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, sbox_inst_16_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_t4_AND_U1 ( .a ({input0_s2[64], input0_s1[64], input0_s0[64]}), .b ({input0_s2[65], input0_s1[65], input0_s0[65]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, sbox_inst_16_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U12 ( .a ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, sbox_inst_15_T3}), .b ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, sbox_inst_15_n17}), .c ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, sbox_inst_15_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U6 ( .a ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, sbox_inst_15_T4}), .b ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, sbox_inst_15_T2}), .c ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, sbox_inst_15_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U5 ( .a ({new_AGEMA_signal_1584, new_AGEMA_signal_1583, sbox_inst_15_T1}), .b ({input0_s2[62], input0_s1[62], input0_s0[62]}), .c ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, sbox_inst_15_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U4 ( .a ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, sbox_inst_15_n11}), .b ({input0_s2[61], input0_s1[61], input0_s0[61]}), .c ({output0_s2[15], output0_s1[15], output0_s0[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U3 ( .a ({input0_s2[63], input0_s1[63], input0_s0[63]}), .b ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, sbox_inst_15_n17}), .c ({new_AGEMA_signal_2512, new_AGEMA_signal_2511, sbox_inst_15_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U2 ( .a ({input0_s2[60], input0_s1[60], input0_s0[60]}), .b ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, sbox_inst_15_T0}), .c ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, sbox_inst_15_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_t0_AND_U1 ( .a ({input0_s2[61], input0_s1[61], input0_s0[61]}), .b ({input0_s2[62], input0_s1[62], input0_s0[62]}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1578, new_AGEMA_signal_1577, sbox_inst_15_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_t1_AND_U1 ( .a ({input0_s2[60], input0_s1[60], input0_s0[60]}), .b ({input0_s2[63], input0_s1[63], input0_s0[63]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_1584, new_AGEMA_signal_1583, sbox_inst_15_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_t2_AND_U1 ( .a ({input0_s2[61], input0_s1[61], input0_s0[61]}), .b ({input0_s2[63], input0_s1[63], input0_s0[63]}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, sbox_inst_15_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_t3_AND_U1 ( .a ({input0_s2[62], input0_s1[62], input0_s0[62]}), .b ({input0_s2[63], input0_s1[63], input0_s0[63]}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, sbox_inst_15_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_t4_AND_U1 ( .a ({input0_s2[60], input0_s1[60], input0_s0[60]}), .b ({input0_s2[61], input0_s1[61], input0_s0[61]}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1590, new_AGEMA_signal_1589, sbox_inst_15_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U12 ( .a ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, sbox_inst_14_T3}), .b ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, sbox_inst_14_n17}), .c ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, sbox_inst_14_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U6 ( .a ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, sbox_inst_14_T4}), .b ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, sbox_inst_14_T2}), .c ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, sbox_inst_14_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U5 ( .a ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, sbox_inst_14_T1}), .b ({input0_s2[58], input0_s1[58], input0_s0[58]}), .c ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, sbox_inst_14_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U4 ( .a ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, sbox_inst_14_n11}), .b ({input0_s2[57], input0_s1[57], input0_s0[57]}), .c ({output0_s2[14], output0_s1[14], output0_s0[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U3 ( .a ({input0_s2[59], input0_s1[59], input0_s0[59]}), .b ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, sbox_inst_14_n17}), .c ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, sbox_inst_14_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U2 ( .a ({input0_s2[56], input0_s1[56], input0_s0[56]}), .b ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, sbox_inst_14_T0}), .c ({new_AGEMA_signal_2112, new_AGEMA_signal_2111, sbox_inst_14_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_t0_AND_U1 ( .a ({input0_s2[57], input0_s1[57], input0_s0[57]}), .b ({input0_s2[58], input0_s1[58], input0_s0[58]}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, sbox_inst_14_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_t1_AND_U1 ( .a ({input0_s2[56], input0_s1[56], input0_s0[56]}), .b ({input0_s2[59], input0_s1[59], input0_s0[59]}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, sbox_inst_14_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_t2_AND_U1 ( .a ({input0_s2[57], input0_s1[57], input0_s0[57]}), .b ({input0_s2[59], input0_s1[59], input0_s0[59]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, sbox_inst_14_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_t3_AND_U1 ( .a ({input0_s2[58], input0_s1[58], input0_s0[58]}), .b ({input0_s2[59], input0_s1[59], input0_s0[59]}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, sbox_inst_14_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_t4_AND_U1 ( .a ({input0_s2[56], input0_s1[56], input0_s0[56]}), .b ({input0_s2[57], input0_s1[57], input0_s0[57]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, sbox_inst_14_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U12 ( .a ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, sbox_inst_13_T3}), .b ({new_AGEMA_signal_2122, new_AGEMA_signal_2121, sbox_inst_13_n17}), .c ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, sbox_inst_13_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U6 ( .a ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, sbox_inst_13_T4}), .b ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, sbox_inst_13_T2}), .c ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, sbox_inst_13_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U5 ( .a ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, sbox_inst_13_T1}), .b ({input0_s2[54], input0_s1[54], input0_s0[54]}), .c ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, sbox_inst_13_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U4 ( .a ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, sbox_inst_13_n11}), .b ({input0_s2[53], input0_s1[53], input0_s0[53]}), .c ({output0_s2[13], output0_s1[13], output0_s0[13]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U3 ( .a ({input0_s2[55], input0_s1[55], input0_s0[55]}), .b ({new_AGEMA_signal_2122, new_AGEMA_signal_2121, sbox_inst_13_n17}), .c ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, sbox_inst_13_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U2 ( .a ({input0_s2[52], input0_s1[52], input0_s0[52]}), .b ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, sbox_inst_13_T0}), .c ({new_AGEMA_signal_2122, new_AGEMA_signal_2121, sbox_inst_13_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_t0_AND_U1 ( .a ({input0_s2[53], input0_s1[53], input0_s0[53]}), .b ({input0_s2[54], input0_s1[54], input0_s0[54]}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, sbox_inst_13_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_t1_AND_U1 ( .a ({input0_s2[52], input0_s1[52], input0_s0[52]}), .b ({input0_s2[55], input0_s1[55], input0_s0[55]}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, sbox_inst_13_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_t2_AND_U1 ( .a ({input0_s2[53], input0_s1[53], input0_s0[53]}), .b ({input0_s2[55], input0_s1[55], input0_s0[55]}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, sbox_inst_13_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_t3_AND_U1 ( .a ({input0_s2[54], input0_s1[54], input0_s0[54]}), .b ({input0_s2[55], input0_s1[55], input0_s0[55]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, sbox_inst_13_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_t4_AND_U1 ( .a ({input0_s2[52], input0_s1[52], input0_s0[52]}), .b ({input0_s2[53], input0_s1[53], input0_s0[53]}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, sbox_inst_13_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U12 ( .a ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, sbox_inst_12_T3}), .b ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, sbox_inst_12_n17}), .c ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, sbox_inst_12_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U6 ( .a ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, sbox_inst_12_T4}), .b ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, sbox_inst_12_T2}), .c ({new_AGEMA_signal_2128, new_AGEMA_signal_2127, sbox_inst_12_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U5 ( .a ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, sbox_inst_12_T1}), .b ({input0_s2[50], input0_s1[50], input0_s0[50]}), .c ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, sbox_inst_12_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U4 ( .a ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, sbox_inst_12_n11}), .b ({input0_s2[49], input0_s1[49], input0_s0[49]}), .c ({output0_s2[12], output0_s1[12], output0_s0[12]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U3 ( .a ({input0_s2[51], input0_s1[51], input0_s0[51]}), .b ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, sbox_inst_12_n17}), .c ({new_AGEMA_signal_2542, new_AGEMA_signal_2541, sbox_inst_12_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U2 ( .a ({input0_s2[48], input0_s1[48], input0_s0[48]}), .b ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, sbox_inst_12_T0}), .c ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, sbox_inst_12_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_t0_AND_U1 ( .a ({input0_s2[49], input0_s1[49], input0_s0[49]}), .b ({input0_s2[50], input0_s1[50], input0_s0[50]}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_1638, new_AGEMA_signal_1637, sbox_inst_12_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_t1_AND_U1 ( .a ({input0_s2[48], input0_s1[48], input0_s0[48]}), .b ({input0_s2[51], input0_s1[51], input0_s0[51]}), .clk (clk), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, sbox_inst_12_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_t2_AND_U1 ( .a ({input0_s2[49], input0_s1[49], input0_s0[49]}), .b ({input0_s2[51], input0_s1[51], input0_s0[51]}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, sbox_inst_12_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_t3_AND_U1 ( .a ({input0_s2[50], input0_s1[50], input0_s0[50]}), .b ({input0_s2[51], input0_s1[51], input0_s0[51]}), .clk (clk), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, sbox_inst_12_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_t4_AND_U1 ( .a ({input0_s2[48], input0_s1[48], input0_s0[48]}), .b ({input0_s2[49], input0_s1[49], input0_s0[49]}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_1650, new_AGEMA_signal_1649, sbox_inst_12_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U12 ( .a ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, sbox_inst_11_T3}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, sbox_inst_11_n17}), .c ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, sbox_inst_11_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U6 ( .a ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, sbox_inst_11_T4}), .b ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, sbox_inst_11_T2}), .c ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, sbox_inst_11_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U5 ( .a ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, sbox_inst_11_T1}), .b ({input0_s2[46], input0_s1[46], input0_s0[46]}), .c ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, sbox_inst_11_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U4 ( .a ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, sbox_inst_11_n11}), .b ({input0_s2[45], input0_s1[45], input0_s0[45]}), .c ({output0_s2[11], output0_s1[11], output0_s0[11]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U3 ( .a ({input0_s2[47], input0_s1[47], input0_s0[47]}), .b ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, sbox_inst_11_n17}), .c ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, sbox_inst_11_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U2 ( .a ({input0_s2[44], input0_s1[44], input0_s0[44]}), .b ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, sbox_inst_11_T0}), .c ({new_AGEMA_signal_2142, new_AGEMA_signal_2141, sbox_inst_11_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_t0_AND_U1 ( .a ({input0_s2[45], input0_s1[45], input0_s0[45]}), .b ({input0_s2[46], input0_s1[46], input0_s0[46]}), .clk (clk), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, sbox_inst_11_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_t1_AND_U1 ( .a ({input0_s2[44], input0_s1[44], input0_s0[44]}), .b ({input0_s2[47], input0_s1[47], input0_s0[47]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, sbox_inst_11_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_t2_AND_U1 ( .a ({input0_s2[45], input0_s1[45], input0_s0[45]}), .b ({input0_s2[47], input0_s1[47], input0_s0[47]}), .clk (clk), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, sbox_inst_11_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_t3_AND_U1 ( .a ({input0_s2[46], input0_s1[46], input0_s0[46]}), .b ({input0_s2[47], input0_s1[47], input0_s0[47]}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, sbox_inst_11_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_t4_AND_U1 ( .a ({input0_s2[44], input0_s1[44], input0_s0[44]}), .b ({input0_s2[45], input0_s1[45], input0_s0[45]}), .clk (clk), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, sbox_inst_11_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U12 ( .a ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, sbox_inst_10_T3}), .b ({new_AGEMA_signal_2152, new_AGEMA_signal_2151, sbox_inst_10_n17}), .c ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, sbox_inst_10_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U6 ( .a ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, sbox_inst_10_T4}), .b ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, sbox_inst_10_T2}), .c ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, sbox_inst_10_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U5 ( .a ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, sbox_inst_10_T1}), .b ({input0_s2[42], input0_s1[42], input0_s0[42]}), .c ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, sbox_inst_10_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U4 ( .a ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, sbox_inst_10_n11}), .b ({input0_s2[41], input0_s1[41], input0_s0[41]}), .c ({output0_s2[10], output0_s1[10], output0_s0[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U3 ( .a ({input0_s2[43], input0_s1[43], input0_s0[43]}), .b ({new_AGEMA_signal_2152, new_AGEMA_signal_2151, sbox_inst_10_n17}), .c ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, sbox_inst_10_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U2 ( .a ({input0_s2[40], input0_s1[40], input0_s0[40]}), .b ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, sbox_inst_10_T0}), .c ({new_AGEMA_signal_2152, new_AGEMA_signal_2151, sbox_inst_10_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_t0_AND_U1 ( .a ({input0_s2[41], input0_s1[41], input0_s0[41]}), .b ({input0_s2[42], input0_s1[42], input0_s0[42]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, sbox_inst_10_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_t1_AND_U1 ( .a ({input0_s2[40], input0_s1[40], input0_s0[40]}), .b ({input0_s2[43], input0_s1[43], input0_s0[43]}), .clk (clk), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, sbox_inst_10_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_t2_AND_U1 ( .a ({input0_s2[41], input0_s1[41], input0_s0[41]}), .b ({input0_s2[43], input0_s1[43], input0_s0[43]}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, sbox_inst_10_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_t3_AND_U1 ( .a ({input0_s2[42], input0_s1[42], input0_s0[42]}), .b ({input0_s2[43], input0_s1[43], input0_s0[43]}), .clk (clk), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, sbox_inst_10_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_t4_AND_U1 ( .a ({input0_s2[40], input0_s1[40], input0_s0[40]}), .b ({input0_s2[41], input0_s1[41], input0_s0[41]}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, sbox_inst_10_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U12 ( .a ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, sbox_inst_9_T3}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, sbox_inst_9_n17}), .c ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, sbox_inst_9_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U6 ( .a ({new_AGEMA_signal_1710, new_AGEMA_signal_1709, sbox_inst_9_T4}), .b ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, sbox_inst_9_T2}), .c ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, sbox_inst_9_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U5 ( .a ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, sbox_inst_9_T1}), .b ({input0_s2[38], input0_s1[38], input0_s0[38]}), .c ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, sbox_inst_9_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U4 ( .a ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, sbox_inst_9_n11}), .b ({input0_s2[37], input0_s1[37], input0_s0[37]}), .c ({output0_s2[9], output0_s1[9], output0_s0[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U3 ( .a ({input0_s2[39], input0_s1[39], input0_s0[39]}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, sbox_inst_9_n17}), .c ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, sbox_inst_9_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U2 ( .a ({input0_s2[36], input0_s1[36], input0_s0[36]}), .b ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, sbox_inst_9_T0}), .c ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, sbox_inst_9_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_t0_AND_U1 ( .a ({input0_s2[37], input0_s1[37], input0_s0[37]}), .b ({input0_s2[38], input0_s1[38], input0_s0[38]}), .clk (clk), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1698, new_AGEMA_signal_1697, sbox_inst_9_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_t1_AND_U1 ( .a ({input0_s2[36], input0_s1[36], input0_s0[36]}), .b ({input0_s2[39], input0_s1[39], input0_s0[39]}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, sbox_inst_9_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_t2_AND_U1 ( .a ({input0_s2[37], input0_s1[37], input0_s0[37]}), .b ({input0_s2[39], input0_s1[39], input0_s0[39]}), .clk (clk), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, sbox_inst_9_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_t3_AND_U1 ( .a ({input0_s2[38], input0_s1[38], input0_s0[38]}), .b ({input0_s2[39], input0_s1[39], input0_s0[39]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, sbox_inst_9_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_t4_AND_U1 ( .a ({input0_s2[36], input0_s1[36], input0_s0[36]}), .b ({input0_s2[37], input0_s1[37], input0_s0[37]}), .clk (clk), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1710, new_AGEMA_signal_1709, sbox_inst_9_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U12 ( .a ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, sbox_inst_8_T3}), .b ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, sbox_inst_8_n17}), .c ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, sbox_inst_8_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U6 ( .a ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, sbox_inst_8_T4}), .b ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, sbox_inst_8_T2}), .c ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, sbox_inst_8_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U5 ( .a ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, sbox_inst_8_T1}), .b ({input0_s2[34], input0_s1[34], input0_s0[34]}), .c ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, sbox_inst_8_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U4 ( .a ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, sbox_inst_8_n11}), .b ({input0_s2[33], input0_s1[33], input0_s0[33]}), .c ({output0_s2[8], output0_s1[8], output0_s0[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U3 ( .a ({input0_s2[35], input0_s1[35], input0_s0[35]}), .b ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, sbox_inst_8_n17}), .c ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, sbox_inst_8_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U2 ( .a ({input0_s2[32], input0_s1[32], input0_s0[32]}), .b ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, sbox_inst_8_T0}), .c ({new_AGEMA_signal_2172, new_AGEMA_signal_2171, sbox_inst_8_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_t0_AND_U1 ( .a ({input0_s2[33], input0_s1[33], input0_s0[33]}), .b ({input0_s2[34], input0_s1[34], input0_s0[34]}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, sbox_inst_8_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_t1_AND_U1 ( .a ({input0_s2[32], input0_s1[32], input0_s0[32]}), .b ({input0_s2[35], input0_s1[35], input0_s0[35]}), .clk (clk), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, sbox_inst_8_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_t2_AND_U1 ( .a ({input0_s2[33], input0_s1[33], input0_s0[33]}), .b ({input0_s2[35], input0_s1[35], input0_s0[35]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, sbox_inst_8_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_t3_AND_U1 ( .a ({input0_s2[34], input0_s1[34], input0_s0[34]}), .b ({input0_s2[35], input0_s1[35], input0_s0[35]}), .clk (clk), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, sbox_inst_8_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_t4_AND_U1 ( .a ({input0_s2[32], input0_s1[32], input0_s0[32]}), .b ({input0_s2[33], input0_s1[33], input0_s0[33]}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, sbox_inst_8_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U12 ( .a ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, sbox_inst_7_T3}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, sbox_inst_7_n17}), .c ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, sbox_inst_7_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U6 ( .a ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, sbox_inst_7_T4}), .b ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, sbox_inst_7_T2}), .c ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, sbox_inst_7_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U5 ( .a ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, sbox_inst_7_T1}), .b ({input0_s2[30], input0_s1[30], input0_s0[30]}), .c ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, sbox_inst_7_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U4 ( .a ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, sbox_inst_7_n11}), .b ({input0_s2[29], input0_s1[29], input0_s0[29]}), .c ({output0_s2[7], output0_s1[7], output0_s0[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U3 ( .a ({input0_s2[31], input0_s1[31], input0_s0[31]}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, sbox_inst_7_n17}), .c ({new_AGEMA_signal_2592, new_AGEMA_signal_2591, sbox_inst_7_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U2 ( .a ({input0_s2[28], input0_s1[28], input0_s0[28]}), .b ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, sbox_inst_7_T0}), .c ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, sbox_inst_7_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_t0_AND_U1 ( .a ({input0_s2[29], input0_s1[29], input0_s0[29]}), .b ({input0_s2[30], input0_s1[30], input0_s0[30]}), .clk (clk), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1738, new_AGEMA_signal_1737, sbox_inst_7_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_t1_AND_U1 ( .a ({input0_s2[28], input0_s1[28], input0_s0[28]}), .b ({input0_s2[31], input0_s1[31], input0_s0[31]}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, sbox_inst_7_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_t2_AND_U1 ( .a ({input0_s2[29], input0_s1[29], input0_s0[29]}), .b ({input0_s2[31], input0_s1[31], input0_s0[31]}), .clk (clk), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, sbox_inst_7_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_t3_AND_U1 ( .a ({input0_s2[30], input0_s1[30], input0_s0[30]}), .b ({input0_s2[31], input0_s1[31], input0_s0[31]}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, sbox_inst_7_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_t4_AND_U1 ( .a ({input0_s2[28], input0_s1[28], input0_s0[28]}), .b ({input0_s2[29], input0_s1[29], input0_s0[29]}), .clk (clk), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1750, new_AGEMA_signal_1749, sbox_inst_7_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U12 ( .a ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, sbox_inst_6_T3}), .b ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, sbox_inst_6_n17}), .c ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, sbox_inst_6_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U6 ( .a ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, sbox_inst_6_T4}), .b ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, sbox_inst_6_T2}), .c ({new_AGEMA_signal_2188, new_AGEMA_signal_2187, sbox_inst_6_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U5 ( .a ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, sbox_inst_6_T1}), .b ({input0_s2[26], input0_s1[26], input0_s0[26]}), .c ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, sbox_inst_6_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U4 ( .a ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, sbox_inst_6_n11}), .b ({input0_s2[25], input0_s1[25], input0_s0[25]}), .c ({output0_s2[6], output0_s1[6], output0_s0[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U3 ( .a ({input0_s2[27], input0_s1[27], input0_s0[27]}), .b ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, sbox_inst_6_n17}), .c ({new_AGEMA_signal_2602, new_AGEMA_signal_2601, sbox_inst_6_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U2 ( .a ({input0_s2[24], input0_s1[24], input0_s0[24]}), .b ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, sbox_inst_6_T0}), .c ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, sbox_inst_6_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_t0_AND_U1 ( .a ({input0_s2[25], input0_s1[25], input0_s0[25]}), .b ({input0_s2[26], input0_s1[26], input0_s0[26]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_1758, new_AGEMA_signal_1757, sbox_inst_6_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_t1_AND_U1 ( .a ({input0_s2[24], input0_s1[24], input0_s0[24]}), .b ({input0_s2[27], input0_s1[27], input0_s0[27]}), .clk (clk), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, sbox_inst_6_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_t2_AND_U1 ( .a ({input0_s2[25], input0_s1[25], input0_s0[25]}), .b ({input0_s2[27], input0_s1[27], input0_s0[27]}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, sbox_inst_6_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_t3_AND_U1 ( .a ({input0_s2[26], input0_s1[26], input0_s0[26]}), .b ({input0_s2[27], input0_s1[27], input0_s0[27]}), .clk (clk), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, sbox_inst_6_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_t4_AND_U1 ( .a ({input0_s2[24], input0_s1[24], input0_s0[24]}), .b ({input0_s2[25], input0_s1[25], input0_s0[25]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_1770, new_AGEMA_signal_1769, sbox_inst_6_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U12 ( .a ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, sbox_inst_5_T3}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, sbox_inst_5_n17}), .c ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, sbox_inst_5_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U6 ( .a ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, sbox_inst_5_T4}), .b ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, sbox_inst_5_T2}), .c ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, sbox_inst_5_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U5 ( .a ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, sbox_inst_5_T1}), .b ({input0_s2[22], input0_s1[22], input0_s0[22]}), .c ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, sbox_inst_5_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U4 ( .a ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, sbox_inst_5_n11}), .b ({input0_s2[21], input0_s1[21], input0_s0[21]}), .c ({output0_s2[5], output0_s1[5], output0_s0[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U3 ( .a ({input0_s2[23], input0_s1[23], input0_s0[23]}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, sbox_inst_5_n17}), .c ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, sbox_inst_5_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U2 ( .a ({input0_s2[20], input0_s1[20], input0_s0[20]}), .b ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, sbox_inst_5_T0}), .c ({new_AGEMA_signal_2202, new_AGEMA_signal_2201, sbox_inst_5_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_t0_AND_U1 ( .a ({input0_s2[21], input0_s1[21], input0_s0[21]}), .b ({input0_s2[22], input0_s1[22], input0_s0[22]}), .clk (clk), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, sbox_inst_5_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_t1_AND_U1 ( .a ({input0_s2[20], input0_s1[20], input0_s0[20]}), .b ({input0_s2[23], input0_s1[23], input0_s0[23]}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, sbox_inst_5_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_t2_AND_U1 ( .a ({input0_s2[21], input0_s1[21], input0_s0[21]}), .b ({input0_s2[23], input0_s1[23], input0_s0[23]}), .clk (clk), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, sbox_inst_5_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_t3_AND_U1 ( .a ({input0_s2[22], input0_s1[22], input0_s0[22]}), .b ({input0_s2[23], input0_s1[23], input0_s0[23]}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, sbox_inst_5_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_t4_AND_U1 ( .a ({input0_s2[20], input0_s1[20], input0_s0[20]}), .b ({input0_s2[21], input0_s1[21], input0_s0[21]}), .clk (clk), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, sbox_inst_5_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U12 ( .a ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, sbox_inst_4_T3}), .b ({new_AGEMA_signal_2212, new_AGEMA_signal_2211, sbox_inst_4_n17}), .c ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, sbox_inst_4_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U6 ( .a ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, sbox_inst_4_T4}), .b ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, sbox_inst_4_T2}), .c ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, sbox_inst_4_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U5 ( .a ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, sbox_inst_4_T1}), .b ({input0_s2[18], input0_s1[18], input0_s0[18]}), .c ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, sbox_inst_4_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U4 ( .a ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, sbox_inst_4_n11}), .b ({input0_s2[17], input0_s1[17], input0_s0[17]}), .c ({output0_s2[4], output0_s1[4], output0_s0[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U3 ( .a ({input0_s2[19], input0_s1[19], input0_s0[19]}), .b ({new_AGEMA_signal_2212, new_AGEMA_signal_2211, sbox_inst_4_n17}), .c ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, sbox_inst_4_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U2 ( .a ({input0_s2[16], input0_s1[16], input0_s0[16]}), .b ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, sbox_inst_4_T0}), .c ({new_AGEMA_signal_2212, new_AGEMA_signal_2211, sbox_inst_4_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_t0_AND_U1 ( .a ({input0_s2[17], input0_s1[17], input0_s0[17]}), .b ({input0_s2[18], input0_s1[18], input0_s0[18]}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, sbox_inst_4_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_t1_AND_U1 ( .a ({input0_s2[16], input0_s1[16], input0_s0[16]}), .b ({input0_s2[19], input0_s1[19], input0_s0[19]}), .clk (clk), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, sbox_inst_4_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_t2_AND_U1 ( .a ({input0_s2[17], input0_s1[17], input0_s0[17]}), .b ({input0_s2[19], input0_s1[19], input0_s0[19]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, sbox_inst_4_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_t3_AND_U1 ( .a ({input0_s2[18], input0_s1[18], input0_s0[18]}), .b ({input0_s2[19], input0_s1[19], input0_s0[19]}), .clk (clk), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, sbox_inst_4_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_t4_AND_U1 ( .a ({input0_s2[16], input0_s1[16], input0_s0[16]}), .b ({input0_s2[17], input0_s1[17], input0_s0[17]}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_1810, new_AGEMA_signal_1809, sbox_inst_4_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U12 ( .a ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, sbox_inst_3_T3}), .b ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, sbox_inst_3_n17}), .c ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, sbox_inst_3_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U6 ( .a ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, sbox_inst_3_T4}), .b ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, sbox_inst_3_T2}), .c ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, sbox_inst_3_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U5 ( .a ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, sbox_inst_3_T1}), .b ({input0_s2[14], input0_s1[14], input0_s0[14]}), .c ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, sbox_inst_3_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U4 ( .a ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, sbox_inst_3_n11}), .b ({input0_s2[13], input0_s1[13], input0_s0[13]}), .c ({output0_s2[3], output0_s1[3], output0_s0[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U3 ( .a ({input0_s2[15], input0_s1[15], input0_s0[15]}), .b ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, sbox_inst_3_n17}), .c ({new_AGEMA_signal_2632, new_AGEMA_signal_2631, sbox_inst_3_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U2 ( .a ({input0_s2[12], input0_s1[12], input0_s0[12]}), .b ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, sbox_inst_3_T0}), .c ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, sbox_inst_3_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_t0_AND_U1 ( .a ({input0_s2[13], input0_s1[13], input0_s0[13]}), .b ({input0_s2[14], input0_s1[14], input0_s0[14]}), .clk (clk), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1818, new_AGEMA_signal_1817, sbox_inst_3_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_t1_AND_U1 ( .a ({input0_s2[12], input0_s1[12], input0_s0[12]}), .b ({input0_s2[15], input0_s1[15], input0_s0[15]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, sbox_inst_3_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_t2_AND_U1 ( .a ({input0_s2[13], input0_s1[13], input0_s0[13]}), .b ({input0_s2[15], input0_s1[15], input0_s0[15]}), .clk (clk), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, sbox_inst_3_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_t3_AND_U1 ( .a ({input0_s2[14], input0_s1[14], input0_s0[14]}), .b ({input0_s2[15], input0_s1[15], input0_s0[15]}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, sbox_inst_3_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_t4_AND_U1 ( .a ({input0_s2[12], input0_s1[12], input0_s0[12]}), .b ({input0_s2[13], input0_s1[13], input0_s0[13]}), .clk (clk), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1830, new_AGEMA_signal_1829, sbox_inst_3_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U12 ( .a ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, sbox_inst_2_T3}), .b ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, sbox_inst_2_n17}), .c ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, sbox_inst_2_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U6 ( .a ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, sbox_inst_2_T4}), .b ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, sbox_inst_2_T2}), .c ({new_AGEMA_signal_2228, new_AGEMA_signal_2227, sbox_inst_2_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U5 ( .a ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, sbox_inst_2_T1}), .b ({input0_s2[10], input0_s1[10], input0_s0[10]}), .c ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, sbox_inst_2_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U4 ( .a ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, sbox_inst_2_n11}), .b ({input0_s2[9], input0_s1[9], input0_s0[9]}), .c ({output0_s2[2], output0_s1[2], output0_s0[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U3 ( .a ({input0_s2[11], input0_s1[11], input0_s0[11]}), .b ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, sbox_inst_2_n17}), .c ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, sbox_inst_2_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U2 ( .a ({input0_s2[8], input0_s1[8], input0_s0[8]}), .b ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, sbox_inst_2_T0}), .c ({new_AGEMA_signal_2232, new_AGEMA_signal_2231, sbox_inst_2_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_t0_AND_U1 ( .a ({input0_s2[9], input0_s1[9], input0_s0[9]}), .b ({input0_s2[10], input0_s1[10], input0_s0[10]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, sbox_inst_2_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_t1_AND_U1 ( .a ({input0_s2[8], input0_s1[8], input0_s0[8]}), .b ({input0_s2[11], input0_s1[11], input0_s0[11]}), .clk (clk), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, sbox_inst_2_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_t2_AND_U1 ( .a ({input0_s2[9], input0_s1[9], input0_s0[9]}), .b ({input0_s2[11], input0_s1[11], input0_s0[11]}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, sbox_inst_2_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_t3_AND_U1 ( .a ({input0_s2[10], input0_s1[10], input0_s0[10]}), .b ({input0_s2[11], input0_s1[11], input0_s0[11]}), .clk (clk), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, sbox_inst_2_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_t4_AND_U1 ( .a ({input0_s2[8], input0_s1[8], input0_s0[8]}), .b ({input0_s2[9], input0_s1[9], input0_s0[9]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, sbox_inst_2_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U12 ( .a ({new_AGEMA_signal_2248, new_AGEMA_signal_2247, sbox_inst_1_T3}), .b ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, sbox_inst_1_n17}), .c ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, sbox_inst_1_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U6 ( .a ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, sbox_inst_1_T4}), .b ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, sbox_inst_1_T2}), .c ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, sbox_inst_1_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U5 ( .a ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, sbox_inst_1_T1}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, input_array_6}), .c ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, sbox_inst_1_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U4 ( .a ({new_AGEMA_signal_2980, new_AGEMA_signal_2979, sbox_inst_1_n11}), .b ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, input_array_5}), .c ({output0_s2[1], output0_s1[1], output0_s0[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U3 ( .a ({input0_s2[7], input0_s1[7], input0_s0[7]}), .b ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, sbox_inst_1_n17}), .c ({new_AGEMA_signal_2980, new_AGEMA_signal_2979, sbox_inst_1_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U2 ( .a ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, input_array_4}), .b ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, sbox_inst_1_T0}), .c ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, sbox_inst_1_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_t0_AND_U1 ( .a ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, input_array_5}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, input_array_6}), .clk (clk), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, sbox_inst_1_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_t1_AND_U1 ( .a ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, input_array_4}), .b ({input0_s2[7], input0_s1[7], input0_s0[7]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, sbox_inst_1_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_t2_AND_U1 ( .a ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, input_array_5}), .b ({input0_s2[7], input0_s1[7], input0_s0[7]}), .clk (clk), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, sbox_inst_1_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_t3_AND_U1 ( .a ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, input_array_6}), .b ({input0_s2[7], input0_s1[7], input0_s0[7]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({new_AGEMA_signal_2248, new_AGEMA_signal_2247, sbox_inst_1_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_t4_AND_U1 ( .a ({new_AGEMA_signal_1098, new_AGEMA_signal_1097, input_array_4}), .b ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, input_array_5}), .clk (clk), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_2250, new_AGEMA_signal_2249, sbox_inst_1_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U12 ( .a ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, sbox_inst_0_T3}), .b ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, sbox_inst_0_n17}), .c ({new_AGEMA_signal_2984, new_AGEMA_signal_2983, sbox_inst_0_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U6 ( .a ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, sbox_inst_0_T4}), .b ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, sbox_inst_0_T2}), .c ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, sbox_inst_0_n13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U5 ( .a ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, sbox_inst_0_T1}), .b ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, input_array_2}), .c ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, sbox_inst_0_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U4 ( .a ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, sbox_inst_0_n11}), .b ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, input_array_1}), .c ({output0_s2[0], output0_s1[0], output0_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U3 ( .a ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, input_array_3}), .b ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, sbox_inst_0_n17}), .c ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, sbox_inst_0_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U2 ( .a ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, input_array_0}), .b ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, sbox_inst_0_T0}), .c ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, sbox_inst_0_n17}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_t0_AND_U1 ( .a ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, input_array_1}), .b ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, input_array_2}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, sbox_inst_0_T0}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_t1_AND_U1 ( .a ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, input_array_0}), .b ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, input_array_3}), .clk (clk), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, sbox_inst_0_T1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_t2_AND_U1 ( .a ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, input_array_1}), .b ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, input_array_3}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, sbox_inst_0_T2}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_t3_AND_U1 ( .a ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, input_array_2}), .b ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, input_array_3}), .clk (clk), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, sbox_inst_0_T3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_t4_AND_U1 ( .a ({new_AGEMA_signal_1110, new_AGEMA_signal_1109, input_array_0}), .b ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, input_array_1}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({new_AGEMA_signal_2262, new_AGEMA_signal_2261, sbox_inst_0_T4}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U15 ( .a ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, sbox_inst_39_T2}), .b ({new_AGEMA_signal_2992, new_AGEMA_signal_2991, sbox_inst_39_n20}), .c ({output0_s2[79], output0_s1[79], output0_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U14 ( .a ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, sbox_inst_39_n19}), .b ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, sbox_inst_39_n18}), .c ({new_AGEMA_signal_2992, new_AGEMA_signal_2991, sbox_inst_39_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U13 ( .a ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, sbox_inst_39_T1}), .b ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, sbox_inst_39_T5}), .c ({new_AGEMA_signal_2664, new_AGEMA_signal_2663, sbox_inst_39_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U11 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, input_array[157]}), .b ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, sbox_inst_39_n16}), .c ({output0_s2[119], output0_s1[119], output0_s0[119]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U10 ( .a ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, sbox_inst_39_n15}), .b ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, sbox_inst_39_T5}), .c ({new_AGEMA_signal_2668, new_AGEMA_signal_2667, sbox_inst_39_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U9 ( .a ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, sbox_inst_39_n15}), .b ({new_AGEMA_signal_2996, new_AGEMA_signal_2995, sbox_inst_39_n14}), .c ({output0_s2[159], output0_s1[159], output0_s0[159]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U8 ( .a ({new_AGEMA_signal_2264, new_AGEMA_signal_2263, sbox_inst_39_n13}), .b ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, sbox_inst_39_n12}), .c ({new_AGEMA_signal_2996, new_AGEMA_signal_2995, sbox_inst_39_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_U7 ( .a ({new_AGEMA_signal_2272, new_AGEMA_signal_2271, sbox_inst_39_T6}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, input_array[159]}), .c ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, sbox_inst_39_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_t5_AND_U1 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, input_array[157]}), .b ({new_AGEMA_signal_1860, new_AGEMA_signal_1859, sbox_inst_39_T3}), .clk (clk), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, sbox_inst_39_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_39_t6_AND_U1 ( .a ({new_AGEMA_signal_1852, new_AGEMA_signal_1851, sbox_inst_39_L0}), .b ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, sbox_inst_39_T1}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({new_AGEMA_signal_2272, new_AGEMA_signal_2271, sbox_inst_39_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U15 ( .a ({new_AGEMA_signal_1872, new_AGEMA_signal_1871, sbox_inst_38_T2}), .b ({new_AGEMA_signal_3000, new_AGEMA_signal_2999, sbox_inst_38_n20}), .c ({output0_s2[78], output0_s1[78], output0_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U14 ( .a ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, sbox_inst_38_n19}), .b ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, sbox_inst_38_n18}), .c ({new_AGEMA_signal_3000, new_AGEMA_signal_2999, sbox_inst_38_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U13 ( .a ({new_AGEMA_signal_1870, new_AGEMA_signal_1869, sbox_inst_38_T1}), .b ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, sbox_inst_38_T5}), .c ({new_AGEMA_signal_2674, new_AGEMA_signal_2673, sbox_inst_38_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U11 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, input_array[153]}), .b ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, sbox_inst_38_n16}), .c ({output0_s2[118], output0_s1[118], output0_s0[118]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U10 ( .a ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, sbox_inst_38_n15}), .b ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, sbox_inst_38_T5}), .c ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, sbox_inst_38_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U9 ( .a ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, sbox_inst_38_n15}), .b ({new_AGEMA_signal_3004, new_AGEMA_signal_3003, sbox_inst_38_n14}), .c ({output0_s2[158], output0_s1[158], output0_s0[158]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U8 ( .a ({new_AGEMA_signal_2274, new_AGEMA_signal_2273, sbox_inst_38_n13}), .b ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, sbox_inst_38_n12}), .c ({new_AGEMA_signal_3004, new_AGEMA_signal_3003, sbox_inst_38_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_U7 ( .a ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, sbox_inst_38_T6}), .b ({new_AGEMA_signal_1126, new_AGEMA_signal_1125, input_array[155]}), .c ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, sbox_inst_38_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_t5_AND_U1 ( .a ({new_AGEMA_signal_1086, new_AGEMA_signal_1085, input_array[153]}), .b ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, sbox_inst_38_T3}), .clk (clk), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_2280, new_AGEMA_signal_2279, sbox_inst_38_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_38_t6_AND_U1 ( .a ({new_AGEMA_signal_1864, new_AGEMA_signal_1863, sbox_inst_38_L0}), .b ({new_AGEMA_signal_1870, new_AGEMA_signal_1869, sbox_inst_38_T1}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, sbox_inst_38_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U15 ( .a ({new_AGEMA_signal_1146, new_AGEMA_signal_1145, sbox_inst_37_T2}), .b ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, sbox_inst_37_n20}), .c ({output0_s2[77], output0_s1[77], output0_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U14 ( .a ({new_AGEMA_signal_2286, new_AGEMA_signal_2285, sbox_inst_37_n19}), .b ({new_AGEMA_signal_2284, new_AGEMA_signal_2283, sbox_inst_37_n18}), .c ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, sbox_inst_37_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U13 ( .a ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, sbox_inst_37_T1}), .b ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, sbox_inst_37_T5}), .c ({new_AGEMA_signal_2284, new_AGEMA_signal_2283, sbox_inst_37_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U11 ( .a ({input0_s2[149], input0_s1[149], input0_s0[149]}), .b ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, sbox_inst_37_n16}), .c ({output0_s2[117], output0_s1[117], output0_s0[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U10 ( .a ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, sbox_inst_37_n15}), .b ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, sbox_inst_37_T5}), .c ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, sbox_inst_37_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U9 ( .a ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, sbox_inst_37_n15}), .b ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, sbox_inst_37_n14}), .c ({output0_s2[157], output0_s1[157], output0_s0[157]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U8 ( .a ({new_AGEMA_signal_1878, new_AGEMA_signal_1877, sbox_inst_37_n13}), .b ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, sbox_inst_37_n12}), .c ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, sbox_inst_37_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_U7 ( .a ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, sbox_inst_37_T6}), .b ({input0_s2[151], input0_s1[151], input0_s0[151]}), .c ({new_AGEMA_signal_2290, new_AGEMA_signal_2289, sbox_inst_37_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_t5_AND_U1 ( .a ({input0_s2[149], input0_s1[149], input0_s0[149]}), .b ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, sbox_inst_37_T3}), .clk (clk), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1884, new_AGEMA_signal_1883, sbox_inst_37_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_37_t6_AND_U1 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, sbox_inst_37_L0}), .b ({new_AGEMA_signal_1144, new_AGEMA_signal_1143, sbox_inst_37_T1}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, sbox_inst_37_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U15 ( .a ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, sbox_inst_36_T2}), .b ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, sbox_inst_36_n20}), .c ({output0_s2[76], output0_s1[76], output0_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U14 ( .a ({new_AGEMA_signal_2296, new_AGEMA_signal_2295, sbox_inst_36_n19}), .b ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, sbox_inst_36_n18}), .c ({new_AGEMA_signal_2692, new_AGEMA_signal_2691, sbox_inst_36_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U13 ( .a ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, sbox_inst_36_T1}), .b ({new_AGEMA_signal_1894, new_AGEMA_signal_1893, sbox_inst_36_T5}), .c ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, sbox_inst_36_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U11 ( .a ({input0_s2[145], input0_s1[145], input0_s0[145]}), .b ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, sbox_inst_36_n16}), .c ({output0_s2[116], output0_s1[116], output0_s0[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U10 ( .a ({new_AGEMA_signal_1890, new_AGEMA_signal_1889, sbox_inst_36_n15}), .b ({new_AGEMA_signal_1894, new_AGEMA_signal_1893, sbox_inst_36_T5}), .c ({new_AGEMA_signal_2298, new_AGEMA_signal_2297, sbox_inst_36_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U9 ( .a ({new_AGEMA_signal_1890, new_AGEMA_signal_1889, sbox_inst_36_n15}), .b ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, sbox_inst_36_n14}), .c ({output0_s2[156], output0_s1[156], output0_s0[156]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U8 ( .a ({new_AGEMA_signal_1888, new_AGEMA_signal_1887, sbox_inst_36_n13}), .b ({new_AGEMA_signal_2300, new_AGEMA_signal_2299, sbox_inst_36_n12}), .c ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, sbox_inst_36_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_U7 ( .a ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, sbox_inst_36_T6}), .b ({input0_s2[147], input0_s1[147], input0_s0[147]}), .c ({new_AGEMA_signal_2300, new_AGEMA_signal_2299, sbox_inst_36_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_t5_AND_U1 ( .a ({input0_s2[145], input0_s1[145], input0_s0[145]}), .b ({new_AGEMA_signal_1168, new_AGEMA_signal_1167, sbox_inst_36_T3}), .clk (clk), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_1894, new_AGEMA_signal_1893, sbox_inst_36_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_36_t6_AND_U1 ( .a ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, sbox_inst_36_L0}), .b ({new_AGEMA_signal_1164, new_AGEMA_signal_1163, sbox_inst_36_T1}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({new_AGEMA_signal_1896, new_AGEMA_signal_1895, sbox_inst_36_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U15 ( .a ({new_AGEMA_signal_1186, new_AGEMA_signal_1185, sbox_inst_35_T2}), .b ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, sbox_inst_35_n20}), .c ({output0_s2[75], output0_s1[75], output0_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U14 ( .a ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, sbox_inst_35_n19}), .b ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, sbox_inst_35_n18}), .c ({new_AGEMA_signal_2700, new_AGEMA_signal_2699, sbox_inst_35_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U13 ( .a ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, sbox_inst_35_T1}), .b ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, sbox_inst_35_T5}), .c ({new_AGEMA_signal_2304, new_AGEMA_signal_2303, sbox_inst_35_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U11 ( .a ({input0_s2[141], input0_s1[141], input0_s0[141]}), .b ({new_AGEMA_signal_2308, new_AGEMA_signal_2307, sbox_inst_35_n16}), .c ({output0_s2[115], output0_s1[115], output0_s0[115]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U10 ( .a ({new_AGEMA_signal_1900, new_AGEMA_signal_1899, sbox_inst_35_n15}), .b ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, sbox_inst_35_T5}), .c ({new_AGEMA_signal_2308, new_AGEMA_signal_2307, sbox_inst_35_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U9 ( .a ({new_AGEMA_signal_1900, new_AGEMA_signal_1899, sbox_inst_35_n15}), .b ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, sbox_inst_35_n14}), .c ({output0_s2[155], output0_s1[155], output0_s0[155]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U8 ( .a ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, sbox_inst_35_n13}), .b ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, sbox_inst_35_n12}), .c ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, sbox_inst_35_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_U7 ( .a ({new_AGEMA_signal_1906, new_AGEMA_signal_1905, sbox_inst_35_T6}), .b ({input0_s2[143], input0_s1[143], input0_s0[143]}), .c ({new_AGEMA_signal_2310, new_AGEMA_signal_2309, sbox_inst_35_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_t5_AND_U1 ( .a ({input0_s2[141], input0_s1[141], input0_s0[141]}), .b ({new_AGEMA_signal_1188, new_AGEMA_signal_1187, sbox_inst_35_T3}), .clk (clk), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, sbox_inst_35_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_35_t6_AND_U1 ( .a ({new_AGEMA_signal_1176, new_AGEMA_signal_1175, sbox_inst_35_L0}), .b ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, sbox_inst_35_T1}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({new_AGEMA_signal_1906, new_AGEMA_signal_1905, sbox_inst_35_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U15 ( .a ({new_AGEMA_signal_1206, new_AGEMA_signal_1205, sbox_inst_34_T2}), .b ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, sbox_inst_34_n20}), .c ({output0_s2[74], output0_s1[74], output0_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U14 ( .a ({new_AGEMA_signal_2316, new_AGEMA_signal_2315, sbox_inst_34_n19}), .b ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, sbox_inst_34_n18}), .c ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, sbox_inst_34_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U13 ( .a ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, sbox_inst_34_T1}), .b ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, sbox_inst_34_T5}), .c ({new_AGEMA_signal_2314, new_AGEMA_signal_2313, sbox_inst_34_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U11 ( .a ({input0_s2[137], input0_s1[137], input0_s0[137]}), .b ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, sbox_inst_34_n16}), .c ({output0_s2[114], output0_s1[114], output0_s0[114]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U10 ( .a ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, sbox_inst_34_n15}), .b ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, sbox_inst_34_T5}), .c ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, sbox_inst_34_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U9 ( .a ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, sbox_inst_34_n15}), .b ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, sbox_inst_34_n14}), .c ({output0_s2[154], output0_s1[154], output0_s0[154]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U8 ( .a ({new_AGEMA_signal_1908, new_AGEMA_signal_1907, sbox_inst_34_n13}), .b ({new_AGEMA_signal_2320, new_AGEMA_signal_2319, sbox_inst_34_n12}), .c ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, sbox_inst_34_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_U7 ( .a ({new_AGEMA_signal_1916, new_AGEMA_signal_1915, sbox_inst_34_T6}), .b ({input0_s2[139], input0_s1[139], input0_s0[139]}), .c ({new_AGEMA_signal_2320, new_AGEMA_signal_2319, sbox_inst_34_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_t5_AND_U1 ( .a ({input0_s2[137], input0_s1[137], input0_s0[137]}), .b ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, sbox_inst_34_T3}), .clk (clk), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_1914, new_AGEMA_signal_1913, sbox_inst_34_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_34_t6_AND_U1 ( .a ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, sbox_inst_34_L0}), .b ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, sbox_inst_34_T1}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({new_AGEMA_signal_1916, new_AGEMA_signal_1915, sbox_inst_34_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U15 ( .a ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, sbox_inst_33_T2}), .b ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, sbox_inst_33_n20}), .c ({output0_s2[73], output0_s1[73], output0_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U14 ( .a ({new_AGEMA_signal_2326, new_AGEMA_signal_2325, sbox_inst_33_n19}), .b ({new_AGEMA_signal_2324, new_AGEMA_signal_2323, sbox_inst_33_n18}), .c ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, sbox_inst_33_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U13 ( .a ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, sbox_inst_33_T1}), .b ({new_AGEMA_signal_1924, new_AGEMA_signal_1923, sbox_inst_33_T5}), .c ({new_AGEMA_signal_2324, new_AGEMA_signal_2323, sbox_inst_33_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U11 ( .a ({input0_s2[133], input0_s1[133], input0_s0[133]}), .b ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, sbox_inst_33_n16}), .c ({output0_s2[113], output0_s1[113], output0_s0[113]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U10 ( .a ({new_AGEMA_signal_1920, new_AGEMA_signal_1919, sbox_inst_33_n15}), .b ({new_AGEMA_signal_1924, new_AGEMA_signal_1923, sbox_inst_33_T5}), .c ({new_AGEMA_signal_2328, new_AGEMA_signal_2327, sbox_inst_33_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U9 ( .a ({new_AGEMA_signal_1920, new_AGEMA_signal_1919, sbox_inst_33_n15}), .b ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, sbox_inst_33_n14}), .c ({output0_s2[153], output0_s1[153], output0_s0[153]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U8 ( .a ({new_AGEMA_signal_1918, new_AGEMA_signal_1917, sbox_inst_33_n13}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, sbox_inst_33_n12}), .c ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, sbox_inst_33_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_U7 ( .a ({new_AGEMA_signal_1926, new_AGEMA_signal_1925, sbox_inst_33_T6}), .b ({input0_s2[135], input0_s1[135], input0_s0[135]}), .c ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, sbox_inst_33_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_t5_AND_U1 ( .a ({input0_s2[133], input0_s1[133], input0_s0[133]}), .b ({new_AGEMA_signal_1228, new_AGEMA_signal_1227, sbox_inst_33_T3}), .clk (clk), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1924, new_AGEMA_signal_1923, sbox_inst_33_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_33_t6_AND_U1 ( .a ({new_AGEMA_signal_1216, new_AGEMA_signal_1215, sbox_inst_33_L0}), .b ({new_AGEMA_signal_1224, new_AGEMA_signal_1223, sbox_inst_33_T1}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({new_AGEMA_signal_1926, new_AGEMA_signal_1925, sbox_inst_33_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U15 ( .a ({new_AGEMA_signal_1246, new_AGEMA_signal_1245, sbox_inst_32_T2}), .b ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, sbox_inst_32_n20}), .c ({output0_s2[72], output0_s1[72], output0_s0[72]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U14 ( .a ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, sbox_inst_32_n19}), .b ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, sbox_inst_32_n18}), .c ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, sbox_inst_32_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U13 ( .a ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, sbox_inst_32_T1}), .b ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, sbox_inst_32_T5}), .c ({new_AGEMA_signal_2334, new_AGEMA_signal_2333, sbox_inst_32_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U11 ( .a ({input0_s2[129], input0_s1[129], input0_s0[129]}), .b ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, sbox_inst_32_n16}), .c ({output0_s2[112], output0_s1[112], output0_s0[112]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U10 ( .a ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, sbox_inst_32_n15}), .b ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, sbox_inst_32_T5}), .c ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, sbox_inst_32_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U9 ( .a ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, sbox_inst_32_n15}), .b ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, sbox_inst_32_n14}), .c ({output0_s2[152], output0_s1[152], output0_s0[152]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U8 ( .a ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, sbox_inst_32_n13}), .b ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, sbox_inst_32_n12}), .c ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, sbox_inst_32_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_U7 ( .a ({new_AGEMA_signal_1936, new_AGEMA_signal_1935, sbox_inst_32_T6}), .b ({input0_s2[131], input0_s1[131], input0_s0[131]}), .c ({new_AGEMA_signal_2340, new_AGEMA_signal_2339, sbox_inst_32_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_t5_AND_U1 ( .a ({input0_s2[129], input0_s1[129], input0_s0[129]}), .b ({new_AGEMA_signal_1248, new_AGEMA_signal_1247, sbox_inst_32_T3}), .clk (clk), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, sbox_inst_32_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_32_t6_AND_U1 ( .a ({new_AGEMA_signal_1236, new_AGEMA_signal_1235, sbox_inst_32_L0}), .b ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, sbox_inst_32_T1}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({new_AGEMA_signal_1936, new_AGEMA_signal_1935, sbox_inst_32_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U15 ( .a ({new_AGEMA_signal_1266, new_AGEMA_signal_1265, sbox_inst_31_T2}), .b ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, sbox_inst_31_n20}), .c ({output0_s2[71], output0_s1[71], output0_s0[71]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U14 ( .a ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, sbox_inst_31_n19}), .b ({new_AGEMA_signal_2344, new_AGEMA_signal_2343, sbox_inst_31_n18}), .c ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, sbox_inst_31_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U13 ( .a ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, sbox_inst_31_T1}), .b ({new_AGEMA_signal_1944, new_AGEMA_signal_1943, sbox_inst_31_T5}), .c ({new_AGEMA_signal_2344, new_AGEMA_signal_2343, sbox_inst_31_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U11 ( .a ({input0_s2[125], input0_s1[125], input0_s0[125]}), .b ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, sbox_inst_31_n16}), .c ({output0_s2[111], output0_s1[111], output0_s0[111]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U10 ( .a ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, sbox_inst_31_n15}), .b ({new_AGEMA_signal_1944, new_AGEMA_signal_1943, sbox_inst_31_T5}), .c ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, sbox_inst_31_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U9 ( .a ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, sbox_inst_31_n15}), .b ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, sbox_inst_31_n14}), .c ({output0_s2[151], output0_s1[151], output0_s0[151]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U8 ( .a ({new_AGEMA_signal_1938, new_AGEMA_signal_1937, sbox_inst_31_n13}), .b ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, sbox_inst_31_n12}), .c ({new_AGEMA_signal_2736, new_AGEMA_signal_2735, sbox_inst_31_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_U7 ( .a ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, sbox_inst_31_T6}), .b ({input0_s2[127], input0_s1[127], input0_s0[127]}), .c ({new_AGEMA_signal_2350, new_AGEMA_signal_2349, sbox_inst_31_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_t5_AND_U1 ( .a ({input0_s2[125], input0_s1[125], input0_s0[125]}), .b ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, sbox_inst_31_T3}), .clk (clk), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1944, new_AGEMA_signal_1943, sbox_inst_31_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_31_t6_AND_U1 ( .a ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, sbox_inst_31_L0}), .b ({new_AGEMA_signal_1264, new_AGEMA_signal_1263, sbox_inst_31_T1}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, sbox_inst_31_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U15 ( .a ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, sbox_inst_30_T2}), .b ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, sbox_inst_30_n20}), .c ({output0_s2[70], output0_s1[70], output0_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U14 ( .a ({new_AGEMA_signal_2356, new_AGEMA_signal_2355, sbox_inst_30_n19}), .b ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, sbox_inst_30_n18}), .c ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, sbox_inst_30_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U13 ( .a ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, sbox_inst_30_T1}), .b ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, sbox_inst_30_T5}), .c ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, sbox_inst_30_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U11 ( .a ({input0_s2[121], input0_s1[121], input0_s0[121]}), .b ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, sbox_inst_30_n16}), .c ({output0_s2[110], output0_s1[110], output0_s0[110]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U10 ( .a ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, sbox_inst_30_n15}), .b ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, sbox_inst_30_T5}), .c ({new_AGEMA_signal_2358, new_AGEMA_signal_2357, sbox_inst_30_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U9 ( .a ({new_AGEMA_signal_1950, new_AGEMA_signal_1949, sbox_inst_30_n15}), .b ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, sbox_inst_30_n14}), .c ({output0_s2[150], output0_s1[150], output0_s0[150]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U8 ( .a ({new_AGEMA_signal_1948, new_AGEMA_signal_1947, sbox_inst_30_n13}), .b ({new_AGEMA_signal_2360, new_AGEMA_signal_2359, sbox_inst_30_n12}), .c ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, sbox_inst_30_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_U7 ( .a ({new_AGEMA_signal_1956, new_AGEMA_signal_1955, sbox_inst_30_T6}), .b ({input0_s2[123], input0_s1[123], input0_s0[123]}), .c ({new_AGEMA_signal_2360, new_AGEMA_signal_2359, sbox_inst_30_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_t5_AND_U1 ( .a ({input0_s2[121], input0_s1[121], input0_s0[121]}), .b ({new_AGEMA_signal_1288, new_AGEMA_signal_1287, sbox_inst_30_T3}), .clk (clk), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, sbox_inst_30_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_30_t6_AND_U1 ( .a ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, sbox_inst_30_L0}), .b ({new_AGEMA_signal_1284, new_AGEMA_signal_1283, sbox_inst_30_T1}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({new_AGEMA_signal_1956, new_AGEMA_signal_1955, sbox_inst_30_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U15 ( .a ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, sbox_inst_29_T2}), .b ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, sbox_inst_29_n20}), .c ({output0_s2[69], output0_s1[69], output0_s0[69]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U14 ( .a ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, sbox_inst_29_n19}), .b ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, sbox_inst_29_n18}), .c ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, sbox_inst_29_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U13 ( .a ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, sbox_inst_29_T1}), .b ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, sbox_inst_29_T5}), .c ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, sbox_inst_29_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U11 ( .a ({input0_s2[117], input0_s1[117], input0_s0[117]}), .b ({new_AGEMA_signal_2368, new_AGEMA_signal_2367, sbox_inst_29_n16}), .c ({output0_s2[109], output0_s1[109], output0_s0[109]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U10 ( .a ({new_AGEMA_signal_1960, new_AGEMA_signal_1959, sbox_inst_29_n15}), .b ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, sbox_inst_29_T5}), .c ({new_AGEMA_signal_2368, new_AGEMA_signal_2367, sbox_inst_29_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U9 ( .a ({new_AGEMA_signal_1960, new_AGEMA_signal_1959, sbox_inst_29_n15}), .b ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, sbox_inst_29_n14}), .c ({output0_s2[149], output0_s1[149], output0_s0[149]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U8 ( .a ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, sbox_inst_29_n13}), .b ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, sbox_inst_29_n12}), .c ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, sbox_inst_29_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_U7 ( .a ({new_AGEMA_signal_1966, new_AGEMA_signal_1965, sbox_inst_29_T6}), .b ({input0_s2[119], input0_s1[119], input0_s0[119]}), .c ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, sbox_inst_29_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_t5_AND_U1 ( .a ({input0_s2[117], input0_s1[117], input0_s0[117]}), .b ({new_AGEMA_signal_1308, new_AGEMA_signal_1307, sbox_inst_29_T3}), .clk (clk), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, sbox_inst_29_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_29_t6_AND_U1 ( .a ({new_AGEMA_signal_1296, new_AGEMA_signal_1295, sbox_inst_29_L0}), .b ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, sbox_inst_29_T1}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({new_AGEMA_signal_1966, new_AGEMA_signal_1965, sbox_inst_29_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U15 ( .a ({new_AGEMA_signal_1326, new_AGEMA_signal_1325, sbox_inst_28_T2}), .b ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, sbox_inst_28_n20}), .c ({output0_s2[68], output0_s1[68], output0_s0[68]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U14 ( .a ({new_AGEMA_signal_2376, new_AGEMA_signal_2375, sbox_inst_28_n19}), .b ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, sbox_inst_28_n18}), .c ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, sbox_inst_28_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U13 ( .a ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, sbox_inst_28_T1}), .b ({new_AGEMA_signal_1974, new_AGEMA_signal_1973, sbox_inst_28_T5}), .c ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, sbox_inst_28_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U11 ( .a ({input0_s2[113], input0_s1[113], input0_s0[113]}), .b ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, sbox_inst_28_n16}), .c ({output0_s2[108], output0_s1[108], output0_s0[108]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U10 ( .a ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, sbox_inst_28_n15}), .b ({new_AGEMA_signal_1974, new_AGEMA_signal_1973, sbox_inst_28_T5}), .c ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, sbox_inst_28_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U9 ( .a ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, sbox_inst_28_n15}), .b ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, sbox_inst_28_n14}), .c ({output0_s2[148], output0_s1[148], output0_s0[148]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U8 ( .a ({new_AGEMA_signal_1968, new_AGEMA_signal_1967, sbox_inst_28_n13}), .b ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, sbox_inst_28_n12}), .c ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, sbox_inst_28_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_U7 ( .a ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, sbox_inst_28_T6}), .b ({input0_s2[115], input0_s1[115], input0_s0[115]}), .c ({new_AGEMA_signal_2380, new_AGEMA_signal_2379, sbox_inst_28_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_t5_AND_U1 ( .a ({input0_s2[113], input0_s1[113], input0_s0[113]}), .b ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, sbox_inst_28_T3}), .clk (clk), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_1974, new_AGEMA_signal_1973, sbox_inst_28_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_28_t6_AND_U1 ( .a ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, sbox_inst_28_L0}), .b ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, sbox_inst_28_T1}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, sbox_inst_28_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U15 ( .a ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, sbox_inst_27_T2}), .b ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, sbox_inst_27_n20}), .c ({output0_s2[67], output0_s1[67], output0_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U14 ( .a ({new_AGEMA_signal_2386, new_AGEMA_signal_2385, sbox_inst_27_n19}), .b ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, sbox_inst_27_n18}), .c ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, sbox_inst_27_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U13 ( .a ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, sbox_inst_27_T1}), .b ({new_AGEMA_signal_1984, new_AGEMA_signal_1983, sbox_inst_27_T5}), .c ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, sbox_inst_27_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U11 ( .a ({input0_s2[109], input0_s1[109], input0_s0[109]}), .b ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, sbox_inst_27_n16}), .c ({output0_s2[107], output0_s1[107], output0_s0[107]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U10 ( .a ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, sbox_inst_27_n15}), .b ({new_AGEMA_signal_1984, new_AGEMA_signal_1983, sbox_inst_27_T5}), .c ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, sbox_inst_27_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U9 ( .a ({new_AGEMA_signal_1980, new_AGEMA_signal_1979, sbox_inst_27_n15}), .b ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, sbox_inst_27_n14}), .c ({output0_s2[147], output0_s1[147], output0_s0[147]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U8 ( .a ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, sbox_inst_27_n13}), .b ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, sbox_inst_27_n12}), .c ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, sbox_inst_27_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_U7 ( .a ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, sbox_inst_27_T6}), .b ({input0_s2[111], input0_s1[111], input0_s0[111]}), .c ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, sbox_inst_27_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_t5_AND_U1 ( .a ({input0_s2[109], input0_s1[109], input0_s0[109]}), .b ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, sbox_inst_27_T3}), .clk (clk), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1984, new_AGEMA_signal_1983, sbox_inst_27_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_27_t6_AND_U1 ( .a ({new_AGEMA_signal_1336, new_AGEMA_signal_1335, sbox_inst_27_L0}), .b ({new_AGEMA_signal_1344, new_AGEMA_signal_1343, sbox_inst_27_T1}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({new_AGEMA_signal_1986, new_AGEMA_signal_1985, sbox_inst_27_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U15 ( .a ({new_AGEMA_signal_1366, new_AGEMA_signal_1365, sbox_inst_26_T2}), .b ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, sbox_inst_26_n20}), .c ({output0_s2[66], output0_s1[66], output0_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U14 ( .a ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, sbox_inst_26_n19}), .b ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, sbox_inst_26_n18}), .c ({new_AGEMA_signal_2772, new_AGEMA_signal_2771, sbox_inst_26_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U13 ( .a ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, sbox_inst_26_T1}), .b ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, sbox_inst_26_T5}), .c ({new_AGEMA_signal_2394, new_AGEMA_signal_2393, sbox_inst_26_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U11 ( .a ({input0_s2[105], input0_s1[105], input0_s0[105]}), .b ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, sbox_inst_26_n16}), .c ({output0_s2[106], output0_s1[106], output0_s0[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U10 ( .a ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, sbox_inst_26_n15}), .b ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, sbox_inst_26_T5}), .c ({new_AGEMA_signal_2398, new_AGEMA_signal_2397, sbox_inst_26_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U9 ( .a ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, sbox_inst_26_n15}), .b ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, sbox_inst_26_n14}), .c ({output0_s2[146], output0_s1[146], output0_s0[146]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U8 ( .a ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, sbox_inst_26_n13}), .b ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, sbox_inst_26_n12}), .c ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, sbox_inst_26_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_U7 ( .a ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, sbox_inst_26_T6}), .b ({input0_s2[107], input0_s1[107], input0_s0[107]}), .c ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, sbox_inst_26_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_t5_AND_U1 ( .a ({input0_s2[105], input0_s1[105], input0_s0[105]}), .b ({new_AGEMA_signal_1368, new_AGEMA_signal_1367, sbox_inst_26_T3}), .clk (clk), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, sbox_inst_26_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_26_t6_AND_U1 ( .a ({new_AGEMA_signal_1356, new_AGEMA_signal_1355, sbox_inst_26_L0}), .b ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, sbox_inst_26_T1}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, sbox_inst_26_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U15 ( .a ({new_AGEMA_signal_1386, new_AGEMA_signal_1385, sbox_inst_25_T2}), .b ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, sbox_inst_25_n20}), .c ({output0_s2[65], output0_s1[65], output0_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U14 ( .a ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, sbox_inst_25_n19}), .b ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, sbox_inst_25_n18}), .c ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, sbox_inst_25_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U13 ( .a ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, sbox_inst_25_T1}), .b ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, sbox_inst_25_T5}), .c ({new_AGEMA_signal_2404, new_AGEMA_signal_2403, sbox_inst_25_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U11 ( .a ({input0_s2[101], input0_s1[101], input0_s0[101]}), .b ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, sbox_inst_25_n16}), .c ({output0_s2[105], output0_s1[105], output0_s0[105]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U10 ( .a ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, sbox_inst_25_n15}), .b ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, sbox_inst_25_T5}), .c ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, sbox_inst_25_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U9 ( .a ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, sbox_inst_25_n15}), .b ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, sbox_inst_25_n14}), .c ({output0_s2[145], output0_s1[145], output0_s0[145]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U8 ( .a ({new_AGEMA_signal_1998, new_AGEMA_signal_1997, sbox_inst_25_n13}), .b ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, sbox_inst_25_n12}), .c ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, sbox_inst_25_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_U7 ( .a ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, sbox_inst_25_T6}), .b ({input0_s2[103], input0_s1[103], input0_s0[103]}), .c ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, sbox_inst_25_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_t5_AND_U1 ( .a ({input0_s2[101], input0_s1[101], input0_s0[101]}), .b ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, sbox_inst_25_T3}), .clk (clk), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_2004, new_AGEMA_signal_2003, sbox_inst_25_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_25_t6_AND_U1 ( .a ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, sbox_inst_25_L0}), .b ({new_AGEMA_signal_1384, new_AGEMA_signal_1383, sbox_inst_25_T1}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, sbox_inst_25_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U15 ( .a ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, sbox_inst_24_T2}), .b ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, sbox_inst_24_n20}), .c ({output0_s2[64], output0_s1[64], output0_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U14 ( .a ({new_AGEMA_signal_2416, new_AGEMA_signal_2415, sbox_inst_24_n19}), .b ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, sbox_inst_24_n18}), .c ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, sbox_inst_24_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U13 ( .a ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, sbox_inst_24_T1}), .b ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, sbox_inst_24_T5}), .c ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, sbox_inst_24_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U11 ( .a ({input0_s2[97], input0_s1[97], input0_s0[97]}), .b ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, sbox_inst_24_n16}), .c ({output0_s2[104], output0_s1[104], output0_s0[104]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U10 ( .a ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, sbox_inst_24_n15}), .b ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, sbox_inst_24_T5}), .c ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, sbox_inst_24_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U9 ( .a ({new_AGEMA_signal_2010, new_AGEMA_signal_2009, sbox_inst_24_n15}), .b ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, sbox_inst_24_n14}), .c ({output0_s2[144], output0_s1[144], output0_s0[144]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U8 ( .a ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, sbox_inst_24_n13}), .b ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, sbox_inst_24_n12}), .c ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, sbox_inst_24_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_U7 ( .a ({new_AGEMA_signal_2016, new_AGEMA_signal_2015, sbox_inst_24_T6}), .b ({input0_s2[99], input0_s1[99], input0_s0[99]}), .c ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, sbox_inst_24_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_t5_AND_U1 ( .a ({input0_s2[97], input0_s1[97], input0_s0[97]}), .b ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, sbox_inst_24_T3}), .clk (clk), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, sbox_inst_24_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_24_t6_AND_U1 ( .a ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, sbox_inst_24_L0}), .b ({new_AGEMA_signal_1404, new_AGEMA_signal_1403, sbox_inst_24_T1}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({new_AGEMA_signal_2016, new_AGEMA_signal_2015, sbox_inst_24_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U15 ( .a ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, sbox_inst_23_T2}), .b ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, sbox_inst_23_n20}), .c ({output0_s2[63], output0_s1[63], output0_s0[63]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U14 ( .a ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, sbox_inst_23_n19}), .b ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, sbox_inst_23_n18}), .c ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, sbox_inst_23_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U13 ( .a ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, sbox_inst_23_T1}), .b ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, sbox_inst_23_T5}), .c ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, sbox_inst_23_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U11 ( .a ({input0_s2[93], input0_s1[93], input0_s0[93]}), .b ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, sbox_inst_23_n16}), .c ({output0_s2[103], output0_s1[103], output0_s0[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U10 ( .a ({new_AGEMA_signal_2020, new_AGEMA_signal_2019, sbox_inst_23_n15}), .b ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, sbox_inst_23_T5}), .c ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, sbox_inst_23_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U9 ( .a ({new_AGEMA_signal_2020, new_AGEMA_signal_2019, sbox_inst_23_n15}), .b ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, sbox_inst_23_n14}), .c ({output0_s2[143], output0_s1[143], output0_s0[143]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U8 ( .a ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, sbox_inst_23_n13}), .b ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, sbox_inst_23_n12}), .c ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, sbox_inst_23_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_U7 ( .a ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, sbox_inst_23_T6}), .b ({input0_s2[95], input0_s1[95], input0_s0[95]}), .c ({new_AGEMA_signal_2430, new_AGEMA_signal_2429, sbox_inst_23_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_t5_AND_U1 ( .a ({input0_s2[93], input0_s1[93], input0_s0[93]}), .b ({new_AGEMA_signal_1428, new_AGEMA_signal_1427, sbox_inst_23_T3}), .clk (clk), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, sbox_inst_23_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_23_t6_AND_U1 ( .a ({new_AGEMA_signal_1416, new_AGEMA_signal_1415, sbox_inst_23_L0}), .b ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, sbox_inst_23_T1}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, sbox_inst_23_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U15 ( .a ({new_AGEMA_signal_1446, new_AGEMA_signal_1445, sbox_inst_22_T2}), .b ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, sbox_inst_22_n20}), .c ({output0_s2[62], output0_s1[62], output0_s0[62]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U14 ( .a ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, sbox_inst_22_n19}), .b ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, sbox_inst_22_n18}), .c ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, sbox_inst_22_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U13 ( .a ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, sbox_inst_22_T1}), .b ({new_AGEMA_signal_2034, new_AGEMA_signal_2033, sbox_inst_22_T5}), .c ({new_AGEMA_signal_2434, new_AGEMA_signal_2433, sbox_inst_22_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U11 ( .a ({input0_s2[89], input0_s1[89], input0_s0[89]}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, sbox_inst_22_n16}), .c ({output0_s2[102], output0_s1[102], output0_s0[102]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U10 ( .a ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, sbox_inst_22_n15}), .b ({new_AGEMA_signal_2034, new_AGEMA_signal_2033, sbox_inst_22_T5}), .c ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, sbox_inst_22_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U9 ( .a ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, sbox_inst_22_n15}), .b ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, sbox_inst_22_n14}), .c ({output0_s2[142], output0_s1[142], output0_s0[142]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U8 ( .a ({new_AGEMA_signal_2028, new_AGEMA_signal_2027, sbox_inst_22_n13}), .b ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, sbox_inst_22_n12}), .c ({new_AGEMA_signal_2808, new_AGEMA_signal_2807, sbox_inst_22_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_U7 ( .a ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, sbox_inst_22_T6}), .b ({input0_s2[91], input0_s1[91], input0_s0[91]}), .c ({new_AGEMA_signal_2440, new_AGEMA_signal_2439, sbox_inst_22_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_t5_AND_U1 ( .a ({input0_s2[89], input0_s1[89], input0_s0[89]}), .b ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, sbox_inst_22_T3}), .clk (clk), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_2034, new_AGEMA_signal_2033, sbox_inst_22_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_22_t6_AND_U1 ( .a ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, sbox_inst_22_L0}), .b ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, sbox_inst_22_T1}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, sbox_inst_22_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U15 ( .a ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, sbox_inst_21_T2}), .b ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, sbox_inst_21_n20}), .c ({output0_s2[61], output0_s1[61], output0_s0[61]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U14 ( .a ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, sbox_inst_21_n19}), .b ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, sbox_inst_21_n18}), .c ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, sbox_inst_21_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U13 ( .a ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, sbox_inst_21_T1}), .b ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, sbox_inst_21_T5}), .c ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, sbox_inst_21_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U11 ( .a ({input0_s2[85], input0_s1[85], input0_s0[85]}), .b ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, sbox_inst_21_n16}), .c ({output0_s2[101], output0_s1[101], output0_s0[101]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U10 ( .a ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, sbox_inst_21_n15}), .b ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, sbox_inst_21_T5}), .c ({new_AGEMA_signal_2448, new_AGEMA_signal_2447, sbox_inst_21_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U9 ( .a ({new_AGEMA_signal_2040, new_AGEMA_signal_2039, sbox_inst_21_n15}), .b ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, sbox_inst_21_n14}), .c ({output0_s2[141], output0_s1[141], output0_s0[141]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U8 ( .a ({new_AGEMA_signal_2038, new_AGEMA_signal_2037, sbox_inst_21_n13}), .b ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, sbox_inst_21_n12}), .c ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, sbox_inst_21_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_U7 ( .a ({new_AGEMA_signal_2046, new_AGEMA_signal_2045, sbox_inst_21_T6}), .b ({input0_s2[87], input0_s1[87], input0_s0[87]}), .c ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, sbox_inst_21_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_t5_AND_U1 ( .a ({input0_s2[85], input0_s1[85], input0_s0[85]}), .b ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, sbox_inst_21_T3}), .clk (clk), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, sbox_inst_21_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_21_t6_AND_U1 ( .a ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, sbox_inst_21_L0}), .b ({new_AGEMA_signal_1464, new_AGEMA_signal_1463, sbox_inst_21_T1}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({new_AGEMA_signal_2046, new_AGEMA_signal_2045, sbox_inst_21_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U15 ( .a ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, sbox_inst_20_T2}), .b ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, sbox_inst_20_n20}), .c ({output0_s2[60], output0_s1[60], output0_s0[60]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U14 ( .a ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, sbox_inst_20_n19}), .b ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, sbox_inst_20_n18}), .c ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, sbox_inst_20_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U13 ( .a ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, sbox_inst_20_T1}), .b ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, sbox_inst_20_T5}), .c ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, sbox_inst_20_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U11 ( .a ({input0_s2[81], input0_s1[81], input0_s0[81]}), .b ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, sbox_inst_20_n16}), .c ({output0_s2[100], output0_s1[100], output0_s0[100]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U10 ( .a ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, sbox_inst_20_n15}), .b ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, sbox_inst_20_T5}), .c ({new_AGEMA_signal_2458, new_AGEMA_signal_2457, sbox_inst_20_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U9 ( .a ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, sbox_inst_20_n15}), .b ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, sbox_inst_20_n14}), .c ({output0_s2[140], output0_s1[140], output0_s0[140]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U8 ( .a ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, sbox_inst_20_n13}), .b ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, sbox_inst_20_n12}), .c ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, sbox_inst_20_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_U7 ( .a ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, sbox_inst_20_T6}), .b ({input0_s2[83], input0_s1[83], input0_s0[83]}), .c ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, sbox_inst_20_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_t5_AND_U1 ( .a ({input0_s2[81], input0_s1[81], input0_s0[81]}), .b ({new_AGEMA_signal_1488, new_AGEMA_signal_1487, sbox_inst_20_T3}), .clk (clk), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, sbox_inst_20_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_20_t6_AND_U1 ( .a ({new_AGEMA_signal_1476, new_AGEMA_signal_1475, sbox_inst_20_L0}), .b ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, sbox_inst_20_T1}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, sbox_inst_20_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U15 ( .a ({new_AGEMA_signal_1506, new_AGEMA_signal_1505, sbox_inst_19_T2}), .b ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, sbox_inst_19_n20}), .c ({output0_s2[59], output0_s1[59], output0_s0[59]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U14 ( .a ({new_AGEMA_signal_2466, new_AGEMA_signal_2465, sbox_inst_19_n19}), .b ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, sbox_inst_19_n18}), .c ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, sbox_inst_19_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U13 ( .a ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, sbox_inst_19_T1}), .b ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, sbox_inst_19_T5}), .c ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, sbox_inst_19_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U11 ( .a ({input0_s2[77], input0_s1[77], input0_s0[77]}), .b ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, sbox_inst_19_n16}), .c ({output0_s2[99], output0_s1[99], output0_s0[99]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U10 ( .a ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, sbox_inst_19_n15}), .b ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, sbox_inst_19_T5}), .c ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, sbox_inst_19_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U9 ( .a ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, sbox_inst_19_n15}), .b ({new_AGEMA_signal_2832, new_AGEMA_signal_2831, sbox_inst_19_n14}), .c ({output0_s2[139], output0_s1[139], output0_s0[139]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U8 ( .a ({new_AGEMA_signal_2058, new_AGEMA_signal_2057, sbox_inst_19_n13}), .b ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, sbox_inst_19_n12}), .c ({new_AGEMA_signal_2832, new_AGEMA_signal_2831, sbox_inst_19_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_U7 ( .a ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, sbox_inst_19_T6}), .b ({input0_s2[79], input0_s1[79], input0_s0[79]}), .c ({new_AGEMA_signal_2470, new_AGEMA_signal_2469, sbox_inst_19_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_t5_AND_U1 ( .a ({input0_s2[77], input0_s1[77], input0_s0[77]}), .b ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, sbox_inst_19_T3}), .clk (clk), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_2064, new_AGEMA_signal_2063, sbox_inst_19_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_19_t6_AND_U1 ( .a ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, sbox_inst_19_L0}), .b ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, sbox_inst_19_T1}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, sbox_inst_19_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U15 ( .a ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, sbox_inst_18_T2}), .b ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, sbox_inst_18_n20}), .c ({output0_s2[58], output0_s1[58], output0_s0[58]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U14 ( .a ({new_AGEMA_signal_2476, new_AGEMA_signal_2475, sbox_inst_18_n19}), .b ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, sbox_inst_18_n18}), .c ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, sbox_inst_18_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U13 ( .a ({new_AGEMA_signal_1524, new_AGEMA_signal_1523, sbox_inst_18_T1}), .b ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, sbox_inst_18_T5}), .c ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, sbox_inst_18_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U11 ( .a ({input0_s2[73], input0_s1[73], input0_s0[73]}), .b ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, sbox_inst_18_n16}), .c ({output0_s2[98], output0_s1[98], output0_s0[98]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U10 ( .a ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, sbox_inst_18_n15}), .b ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, sbox_inst_18_T5}), .c ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, sbox_inst_18_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U9 ( .a ({new_AGEMA_signal_2070, new_AGEMA_signal_2069, sbox_inst_18_n15}), .b ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, sbox_inst_18_n14}), .c ({output0_s2[138], output0_s1[138], output0_s0[138]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U8 ( .a ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, sbox_inst_18_n13}), .b ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, sbox_inst_18_n12}), .c ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, sbox_inst_18_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_U7 ( .a ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, sbox_inst_18_T6}), .b ({input0_s2[75], input0_s1[75], input0_s0[75]}), .c ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, sbox_inst_18_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_t5_AND_U1 ( .a ({input0_s2[73], input0_s1[73], input0_s0[73]}), .b ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, sbox_inst_18_T3}), .clk (clk), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, sbox_inst_18_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_18_t6_AND_U1 ( .a ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, sbox_inst_18_L0}), .b ({new_AGEMA_signal_1524, new_AGEMA_signal_1523, sbox_inst_18_T1}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({new_AGEMA_signal_2076, new_AGEMA_signal_2075, sbox_inst_18_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U15 ( .a ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, sbox_inst_17_T2}), .b ({new_AGEMA_signal_2844, new_AGEMA_signal_2843, sbox_inst_17_n20}), .c ({output0_s2[57], output0_s1[57], output0_s0[57]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U14 ( .a ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, sbox_inst_17_n19}), .b ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, sbox_inst_17_n18}), .c ({new_AGEMA_signal_2844, new_AGEMA_signal_2843, sbox_inst_17_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U13 ( .a ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, sbox_inst_17_T1}), .b ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, sbox_inst_17_T5}), .c ({new_AGEMA_signal_2484, new_AGEMA_signal_2483, sbox_inst_17_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U11 ( .a ({input0_s2[69], input0_s1[69], input0_s0[69]}), .b ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, sbox_inst_17_n16}), .c ({output0_s2[97], output0_s1[97], output0_s0[97]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U10 ( .a ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, sbox_inst_17_n15}), .b ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, sbox_inst_17_T5}), .c ({new_AGEMA_signal_2488, new_AGEMA_signal_2487, sbox_inst_17_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U9 ( .a ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, sbox_inst_17_n15}), .b ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, sbox_inst_17_n14}), .c ({output0_s2[137], output0_s1[137], output0_s0[137]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U8 ( .a ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, sbox_inst_17_n13}), .b ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, sbox_inst_17_n12}), .c ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, sbox_inst_17_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_U7 ( .a ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, sbox_inst_17_T6}), .b ({input0_s2[71], input0_s1[71], input0_s0[71]}), .c ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, sbox_inst_17_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_t5_AND_U1 ( .a ({input0_s2[69], input0_s1[69], input0_s0[69]}), .b ({new_AGEMA_signal_1548, new_AGEMA_signal_1547, sbox_inst_17_T3}), .clk (clk), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, sbox_inst_17_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_17_t6_AND_U1 ( .a ({new_AGEMA_signal_1536, new_AGEMA_signal_1535, sbox_inst_17_L0}), .b ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, sbox_inst_17_T1}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, sbox_inst_17_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U15 ( .a ({new_AGEMA_signal_1566, new_AGEMA_signal_1565, sbox_inst_16_T2}), .b ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, sbox_inst_16_n20}), .c ({output0_s2[56], output0_s1[56], output0_s0[56]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U14 ( .a ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, sbox_inst_16_n19}), .b ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, sbox_inst_16_n18}), .c ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, sbox_inst_16_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U13 ( .a ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, sbox_inst_16_T1}), .b ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, sbox_inst_16_T5}), .c ({new_AGEMA_signal_2494, new_AGEMA_signal_2493, sbox_inst_16_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U11 ( .a ({input0_s2[65], input0_s1[65], input0_s0[65]}), .b ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, sbox_inst_16_n16}), .c ({output0_s2[96], output0_s1[96], output0_s0[96]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U10 ( .a ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, sbox_inst_16_n15}), .b ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, sbox_inst_16_T5}), .c ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, sbox_inst_16_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U9 ( .a ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, sbox_inst_16_n15}), .b ({new_AGEMA_signal_2856, new_AGEMA_signal_2855, sbox_inst_16_n14}), .c ({output0_s2[136], output0_s1[136], output0_s0[136]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U8 ( .a ({new_AGEMA_signal_2088, new_AGEMA_signal_2087, sbox_inst_16_n13}), .b ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, sbox_inst_16_n12}), .c ({new_AGEMA_signal_2856, new_AGEMA_signal_2855, sbox_inst_16_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_U7 ( .a ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, sbox_inst_16_T6}), .b ({input0_s2[67], input0_s1[67], input0_s0[67]}), .c ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, sbox_inst_16_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_t5_AND_U1 ( .a ({input0_s2[65], input0_s1[65], input0_s0[65]}), .b ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, sbox_inst_16_T3}), .clk (clk), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_2094, new_AGEMA_signal_2093, sbox_inst_16_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_16_t6_AND_U1 ( .a ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, sbox_inst_16_L0}), .b ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, sbox_inst_16_T1}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, sbox_inst_16_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U15 ( .a ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, sbox_inst_15_T2}), .b ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, sbox_inst_15_n20}), .c ({output0_s2[55], output0_s1[55], output0_s0[55]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U14 ( .a ({new_AGEMA_signal_2506, new_AGEMA_signal_2505, sbox_inst_15_n19}), .b ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, sbox_inst_15_n18}), .c ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, sbox_inst_15_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U13 ( .a ({new_AGEMA_signal_1584, new_AGEMA_signal_1583, sbox_inst_15_T1}), .b ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, sbox_inst_15_T5}), .c ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, sbox_inst_15_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U11 ( .a ({input0_s2[61], input0_s1[61], input0_s0[61]}), .b ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, sbox_inst_15_n16}), .c ({output0_s2[95], output0_s1[95], output0_s0[95]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U10 ( .a ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, sbox_inst_15_n15}), .b ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, sbox_inst_15_T5}), .c ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, sbox_inst_15_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U9 ( .a ({new_AGEMA_signal_2100, new_AGEMA_signal_2099, sbox_inst_15_n15}), .b ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, sbox_inst_15_n14}), .c ({output0_s2[135], output0_s1[135], output0_s0[135]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U8 ( .a ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, sbox_inst_15_n13}), .b ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, sbox_inst_15_n12}), .c ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, sbox_inst_15_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_U7 ( .a ({new_AGEMA_signal_2106, new_AGEMA_signal_2105, sbox_inst_15_T6}), .b ({input0_s2[63], input0_s1[63], input0_s0[63]}), .c ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, sbox_inst_15_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_t5_AND_U1 ( .a ({input0_s2[61], input0_s1[61], input0_s0[61]}), .b ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, sbox_inst_15_T3}), .clk (clk), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, sbox_inst_15_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_15_t6_AND_U1 ( .a ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, sbox_inst_15_L0}), .b ({new_AGEMA_signal_1584, new_AGEMA_signal_1583, sbox_inst_15_T1}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({new_AGEMA_signal_2106, new_AGEMA_signal_2105, sbox_inst_15_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U15 ( .a ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, sbox_inst_14_T2}), .b ({new_AGEMA_signal_2868, new_AGEMA_signal_2867, sbox_inst_14_n20}), .c ({output0_s2[54], output0_s1[54], output0_s0[54]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U14 ( .a ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, sbox_inst_14_n19}), .b ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, sbox_inst_14_n18}), .c ({new_AGEMA_signal_2868, new_AGEMA_signal_2867, sbox_inst_14_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U13 ( .a ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, sbox_inst_14_T1}), .b ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, sbox_inst_14_T5}), .c ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, sbox_inst_14_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U11 ( .a ({input0_s2[57], input0_s1[57], input0_s0[57]}), .b ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, sbox_inst_14_n16}), .c ({output0_s2[94], output0_s1[94], output0_s0[94]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U10 ( .a ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, sbox_inst_14_n15}), .b ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, sbox_inst_14_T5}), .c ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, sbox_inst_14_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U9 ( .a ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, sbox_inst_14_n15}), .b ({new_AGEMA_signal_2872, new_AGEMA_signal_2871, sbox_inst_14_n14}), .c ({output0_s2[134], output0_s1[134], output0_s0[134]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U8 ( .a ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, sbox_inst_14_n13}), .b ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, sbox_inst_14_n12}), .c ({new_AGEMA_signal_2872, new_AGEMA_signal_2871, sbox_inst_14_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_U7 ( .a ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, sbox_inst_14_T6}), .b ({input0_s2[59], input0_s1[59], input0_s0[59]}), .c ({new_AGEMA_signal_2520, new_AGEMA_signal_2519, sbox_inst_14_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_t5_AND_U1 ( .a ({input0_s2[57], input0_s1[57], input0_s0[57]}), .b ({new_AGEMA_signal_1608, new_AGEMA_signal_1607, sbox_inst_14_T3}), .clk (clk), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, sbox_inst_14_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_14_t6_AND_U1 ( .a ({new_AGEMA_signal_1596, new_AGEMA_signal_1595, sbox_inst_14_L0}), .b ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, sbox_inst_14_T1}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, sbox_inst_14_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U15 ( .a ({new_AGEMA_signal_1626, new_AGEMA_signal_1625, sbox_inst_13_T2}), .b ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, sbox_inst_13_n20}), .c ({output0_s2[53], output0_s1[53], output0_s0[53]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U14 ( .a ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, sbox_inst_13_n19}), .b ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, sbox_inst_13_n18}), .c ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, sbox_inst_13_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U13 ( .a ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, sbox_inst_13_T1}), .b ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, sbox_inst_13_T5}), .c ({new_AGEMA_signal_2524, new_AGEMA_signal_2523, sbox_inst_13_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U11 ( .a ({input0_s2[53], input0_s1[53], input0_s0[53]}), .b ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, sbox_inst_13_n16}), .c ({output0_s2[93], output0_s1[93], output0_s0[93]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U10 ( .a ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, sbox_inst_13_n15}), .b ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, sbox_inst_13_T5}), .c ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, sbox_inst_13_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U9 ( .a ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, sbox_inst_13_n15}), .b ({new_AGEMA_signal_2880, new_AGEMA_signal_2879, sbox_inst_13_n14}), .c ({output0_s2[133], output0_s1[133], output0_s0[133]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U8 ( .a ({new_AGEMA_signal_2118, new_AGEMA_signal_2117, sbox_inst_13_n13}), .b ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, sbox_inst_13_n12}), .c ({new_AGEMA_signal_2880, new_AGEMA_signal_2879, sbox_inst_13_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_U7 ( .a ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, sbox_inst_13_T6}), .b ({input0_s2[55], input0_s1[55], input0_s0[55]}), .c ({new_AGEMA_signal_2530, new_AGEMA_signal_2529, sbox_inst_13_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_t5_AND_U1 ( .a ({input0_s2[53], input0_s1[53], input0_s0[53]}), .b ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, sbox_inst_13_T3}), .clk (clk), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_2124, new_AGEMA_signal_2123, sbox_inst_13_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_13_t6_AND_U1 ( .a ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, sbox_inst_13_L0}), .b ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, sbox_inst_13_T1}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, sbox_inst_13_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U15 ( .a ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, sbox_inst_12_T2}), .b ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, sbox_inst_12_n20}), .c ({output0_s2[52], output0_s1[52], output0_s0[52]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U14 ( .a ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, sbox_inst_12_n19}), .b ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, sbox_inst_12_n18}), .c ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, sbox_inst_12_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U13 ( .a ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, sbox_inst_12_T1}), .b ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, sbox_inst_12_T5}), .c ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, sbox_inst_12_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U11 ( .a ({input0_s2[49], input0_s1[49], input0_s0[49]}), .b ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, sbox_inst_12_n16}), .c ({output0_s2[92], output0_s1[92], output0_s0[92]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U10 ( .a ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, sbox_inst_12_n15}), .b ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, sbox_inst_12_T5}), .c ({new_AGEMA_signal_2538, new_AGEMA_signal_2537, sbox_inst_12_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U9 ( .a ({new_AGEMA_signal_2130, new_AGEMA_signal_2129, sbox_inst_12_n15}), .b ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, sbox_inst_12_n14}), .c ({output0_s2[132], output0_s1[132], output0_s0[132]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U8 ( .a ({new_AGEMA_signal_2128, new_AGEMA_signal_2127, sbox_inst_12_n13}), .b ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, sbox_inst_12_n12}), .c ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, sbox_inst_12_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_U7 ( .a ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, sbox_inst_12_T6}), .b ({input0_s2[51], input0_s1[51], input0_s0[51]}), .c ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, sbox_inst_12_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_t5_AND_U1 ( .a ({input0_s2[49], input0_s1[49], input0_s0[49]}), .b ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, sbox_inst_12_T3}), .clk (clk), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, sbox_inst_12_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_12_t6_AND_U1 ( .a ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, sbox_inst_12_L0}), .b ({new_AGEMA_signal_1644, new_AGEMA_signal_1643, sbox_inst_12_T1}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({new_AGEMA_signal_2136, new_AGEMA_signal_2135, sbox_inst_12_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U15 ( .a ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, sbox_inst_11_T2}), .b ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, sbox_inst_11_n20}), .c ({output0_s2[51], output0_s1[51], output0_s0[51]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U14 ( .a ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, sbox_inst_11_n19}), .b ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, sbox_inst_11_n18}), .c ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, sbox_inst_11_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U13 ( .a ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, sbox_inst_11_T1}), .b ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, sbox_inst_11_T5}), .c ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, sbox_inst_11_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U11 ( .a ({input0_s2[45], input0_s1[45], input0_s0[45]}), .b ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, sbox_inst_11_n16}), .c ({output0_s2[91], output0_s1[91], output0_s0[91]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U10 ( .a ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, sbox_inst_11_n15}), .b ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, sbox_inst_11_T5}), .c ({new_AGEMA_signal_2548, new_AGEMA_signal_2547, sbox_inst_11_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U9 ( .a ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, sbox_inst_11_n15}), .b ({new_AGEMA_signal_2896, new_AGEMA_signal_2895, sbox_inst_11_n14}), .c ({output0_s2[131], output0_s1[131], output0_s0[131]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U8 ( .a ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, sbox_inst_11_n13}), .b ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, sbox_inst_11_n12}), .c ({new_AGEMA_signal_2896, new_AGEMA_signal_2895, sbox_inst_11_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_U7 ( .a ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, sbox_inst_11_T6}), .b ({input0_s2[47], input0_s1[47], input0_s0[47]}), .c ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, sbox_inst_11_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_t5_AND_U1 ( .a ({input0_s2[45], input0_s1[45], input0_s0[45]}), .b ({new_AGEMA_signal_1668, new_AGEMA_signal_1667, sbox_inst_11_T3}), .clk (clk), .r ({Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, sbox_inst_11_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_11_t6_AND_U1 ( .a ({new_AGEMA_signal_1656, new_AGEMA_signal_1655, sbox_inst_11_L0}), .b ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, sbox_inst_11_T1}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771]}), .c ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, sbox_inst_11_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U15 ( .a ({new_AGEMA_signal_1686, new_AGEMA_signal_1685, sbox_inst_10_T2}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, sbox_inst_10_n20}), .c ({output0_s2[50], output0_s1[50], output0_s0[50]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U14 ( .a ({new_AGEMA_signal_2556, new_AGEMA_signal_2555, sbox_inst_10_n19}), .b ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, sbox_inst_10_n18}), .c ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, sbox_inst_10_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U13 ( .a ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, sbox_inst_10_T1}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, sbox_inst_10_T5}), .c ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, sbox_inst_10_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U11 ( .a ({input0_s2[41], input0_s1[41], input0_s0[41]}), .b ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, sbox_inst_10_n16}), .c ({output0_s2[90], output0_s1[90], output0_s0[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U10 ( .a ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, sbox_inst_10_n15}), .b ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, sbox_inst_10_T5}), .c ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, sbox_inst_10_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U9 ( .a ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, sbox_inst_10_n15}), .b ({new_AGEMA_signal_2904, new_AGEMA_signal_2903, sbox_inst_10_n14}), .c ({output0_s2[130], output0_s1[130], output0_s0[130]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U8 ( .a ({new_AGEMA_signal_2148, new_AGEMA_signal_2147, sbox_inst_10_n13}), .b ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, sbox_inst_10_n12}), .c ({new_AGEMA_signal_2904, new_AGEMA_signal_2903, sbox_inst_10_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_U7 ( .a ({new_AGEMA_signal_2156, new_AGEMA_signal_2155, sbox_inst_10_T6}), .b ({input0_s2[43], input0_s1[43], input0_s0[43]}), .c ({new_AGEMA_signal_2560, new_AGEMA_signal_2559, sbox_inst_10_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_t5_AND_U1 ( .a ({input0_s2[41], input0_s1[41], input0_s0[41]}), .b ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, sbox_inst_10_T3}), .clk (clk), .r ({Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_2154, new_AGEMA_signal_2153, sbox_inst_10_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_10_t6_AND_U1 ( .a ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, sbox_inst_10_L0}), .b ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, sbox_inst_10_T1}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777]}), .c ({new_AGEMA_signal_2156, new_AGEMA_signal_2155, sbox_inst_10_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U15 ( .a ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, sbox_inst_9_T2}), .b ({new_AGEMA_signal_2908, new_AGEMA_signal_2907, sbox_inst_9_n20}), .c ({output0_s2[49], output0_s1[49], output0_s0[49]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U14 ( .a ({new_AGEMA_signal_2566, new_AGEMA_signal_2565, sbox_inst_9_n19}), .b ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, sbox_inst_9_n18}), .c ({new_AGEMA_signal_2908, new_AGEMA_signal_2907, sbox_inst_9_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U13 ( .a ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, sbox_inst_9_T1}), .b ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, sbox_inst_9_T5}), .c ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, sbox_inst_9_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U11 ( .a ({input0_s2[37], input0_s1[37], input0_s0[37]}), .b ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, sbox_inst_9_n16}), .c ({output0_s2[89], output0_s1[89], output0_s0[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U10 ( .a ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, sbox_inst_9_n15}), .b ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, sbox_inst_9_T5}), .c ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, sbox_inst_9_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U9 ( .a ({new_AGEMA_signal_2160, new_AGEMA_signal_2159, sbox_inst_9_n15}), .b ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, sbox_inst_9_n14}), .c ({output0_s2[129], output0_s1[129], output0_s0[129]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U8 ( .a ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, sbox_inst_9_n13}), .b ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, sbox_inst_9_n12}), .c ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, sbox_inst_9_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_U7 ( .a ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, sbox_inst_9_T6}), .b ({input0_s2[39], input0_s1[39], input0_s0[39]}), .c ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, sbox_inst_9_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_t5_AND_U1 ( .a ({input0_s2[37], input0_s1[37], input0_s0[37]}), .b ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, sbox_inst_9_T3}), .clk (clk), .r ({Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, sbox_inst_9_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_9_t6_AND_U1 ( .a ({new_AGEMA_signal_1696, new_AGEMA_signal_1695, sbox_inst_9_L0}), .b ({new_AGEMA_signal_1704, new_AGEMA_signal_1703, sbox_inst_9_T1}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783]}), .c ({new_AGEMA_signal_2166, new_AGEMA_signal_2165, sbox_inst_9_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U15 ( .a ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, sbox_inst_8_T2}), .b ({new_AGEMA_signal_2916, new_AGEMA_signal_2915, sbox_inst_8_n20}), .c ({output0_s2[48], output0_s1[48], output0_s0[48]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U14 ( .a ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, sbox_inst_8_n19}), .b ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, sbox_inst_8_n18}), .c ({new_AGEMA_signal_2916, new_AGEMA_signal_2915, sbox_inst_8_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U13 ( .a ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, sbox_inst_8_T1}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, sbox_inst_8_T5}), .c ({new_AGEMA_signal_2574, new_AGEMA_signal_2573, sbox_inst_8_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U11 ( .a ({input0_s2[33], input0_s1[33], input0_s0[33]}), .b ({new_AGEMA_signal_2578, new_AGEMA_signal_2577, sbox_inst_8_n16}), .c ({output0_s2[88], output0_s1[88], output0_s0[88]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U10 ( .a ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, sbox_inst_8_n15}), .b ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, sbox_inst_8_T5}), .c ({new_AGEMA_signal_2578, new_AGEMA_signal_2577, sbox_inst_8_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U9 ( .a ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, sbox_inst_8_n15}), .b ({new_AGEMA_signal_2920, new_AGEMA_signal_2919, sbox_inst_8_n14}), .c ({output0_s2[128], output0_s1[128], output0_s0[128]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U8 ( .a ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, sbox_inst_8_n13}), .b ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, sbox_inst_8_n12}), .c ({new_AGEMA_signal_2920, new_AGEMA_signal_2919, sbox_inst_8_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_U7 ( .a ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, sbox_inst_8_T6}), .b ({input0_s2[35], input0_s1[35], input0_s0[35]}), .c ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, sbox_inst_8_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_t5_AND_U1 ( .a ({input0_s2[33], input0_s1[33], input0_s0[33]}), .b ({new_AGEMA_signal_1728, new_AGEMA_signal_1727, sbox_inst_8_T3}), .clk (clk), .r ({Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, sbox_inst_8_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_8_t6_AND_U1 ( .a ({new_AGEMA_signal_1716, new_AGEMA_signal_1715, sbox_inst_8_L0}), .b ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, sbox_inst_8_T1}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789]}), .c ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, sbox_inst_8_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U15 ( .a ({new_AGEMA_signal_1746, new_AGEMA_signal_1745, sbox_inst_7_T2}), .b ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, sbox_inst_7_n20}), .c ({output0_s2[47], output0_s1[47], output0_s0[47]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U14 ( .a ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, sbox_inst_7_n19}), .b ({new_AGEMA_signal_2584, new_AGEMA_signal_2583, sbox_inst_7_n18}), .c ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, sbox_inst_7_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U13 ( .a ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, sbox_inst_7_T1}), .b ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, sbox_inst_7_T5}), .c ({new_AGEMA_signal_2584, new_AGEMA_signal_2583, sbox_inst_7_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U11 ( .a ({input0_s2[29], input0_s1[29], input0_s0[29]}), .b ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, sbox_inst_7_n16}), .c ({output0_s2[87], output0_s1[87], output0_s0[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U10 ( .a ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, sbox_inst_7_n15}), .b ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, sbox_inst_7_T5}), .c ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, sbox_inst_7_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U9 ( .a ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, sbox_inst_7_n15}), .b ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, sbox_inst_7_n14}), .c ({output0_s2[127], output0_s1[127], output0_s0[127]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U8 ( .a ({new_AGEMA_signal_2178, new_AGEMA_signal_2177, sbox_inst_7_n13}), .b ({new_AGEMA_signal_2590, new_AGEMA_signal_2589, sbox_inst_7_n12}), .c ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, sbox_inst_7_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_U7 ( .a ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, sbox_inst_7_T6}), .b ({input0_s2[31], input0_s1[31], input0_s0[31]}), .c ({new_AGEMA_signal_2590, new_AGEMA_signal_2589, sbox_inst_7_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_t5_AND_U1 ( .a ({input0_s2[29], input0_s1[29], input0_s0[29]}), .b ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, sbox_inst_7_T3}), .clk (clk), .r ({Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_2184, new_AGEMA_signal_2183, sbox_inst_7_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_7_t6_AND_U1 ( .a ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, sbox_inst_7_L0}), .b ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, sbox_inst_7_T1}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795]}), .c ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, sbox_inst_7_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U15 ( .a ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, sbox_inst_6_T2}), .b ({new_AGEMA_signal_2932, new_AGEMA_signal_2931, sbox_inst_6_n20}), .c ({output0_s2[46], output0_s1[46], output0_s0[46]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U14 ( .a ({new_AGEMA_signal_2596, new_AGEMA_signal_2595, sbox_inst_6_n19}), .b ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, sbox_inst_6_n18}), .c ({new_AGEMA_signal_2932, new_AGEMA_signal_2931, sbox_inst_6_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U13 ( .a ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, sbox_inst_6_T1}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, sbox_inst_6_T5}), .c ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, sbox_inst_6_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U11 ( .a ({input0_s2[25], input0_s1[25], input0_s0[25]}), .b ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, sbox_inst_6_n16}), .c ({output0_s2[86], output0_s1[86], output0_s0[86]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U10 ( .a ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, sbox_inst_6_n15}), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, sbox_inst_6_T5}), .c ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, sbox_inst_6_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U9 ( .a ({new_AGEMA_signal_2190, new_AGEMA_signal_2189, sbox_inst_6_n15}), .b ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, sbox_inst_6_n14}), .c ({output0_s2[126], output0_s1[126], output0_s0[126]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U8 ( .a ({new_AGEMA_signal_2188, new_AGEMA_signal_2187, sbox_inst_6_n13}), .b ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, sbox_inst_6_n12}), .c ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, sbox_inst_6_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_U7 ( .a ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, sbox_inst_6_T6}), .b ({input0_s2[27], input0_s1[27], input0_s0[27]}), .c ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, sbox_inst_6_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_t5_AND_U1 ( .a ({input0_s2[25], input0_s1[25], input0_s0[25]}), .b ({new_AGEMA_signal_1768, new_AGEMA_signal_1767, sbox_inst_6_T3}), .clk (clk), .r ({Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, sbox_inst_6_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_6_t6_AND_U1 ( .a ({new_AGEMA_signal_1756, new_AGEMA_signal_1755, sbox_inst_6_L0}), .b ({new_AGEMA_signal_1764, new_AGEMA_signal_1763, sbox_inst_6_T1}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801]}), .c ({new_AGEMA_signal_2196, new_AGEMA_signal_2195, sbox_inst_6_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U15 ( .a ({new_AGEMA_signal_1786, new_AGEMA_signal_1785, sbox_inst_5_T2}), .b ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, sbox_inst_5_n20}), .c ({output0_s2[45], output0_s1[45], output0_s0[45]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U14 ( .a ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, sbox_inst_5_n19}), .b ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, sbox_inst_5_n18}), .c ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, sbox_inst_5_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U13 ( .a ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, sbox_inst_5_T1}), .b ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, sbox_inst_5_T5}), .c ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, sbox_inst_5_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U11 ( .a ({input0_s2[21], input0_s1[21], input0_s0[21]}), .b ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, sbox_inst_5_n16}), .c ({output0_s2[85], output0_s1[85], output0_s0[85]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U10 ( .a ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, sbox_inst_5_n15}), .b ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, sbox_inst_5_T5}), .c ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, sbox_inst_5_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U9 ( .a ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, sbox_inst_5_n15}), .b ({new_AGEMA_signal_2944, new_AGEMA_signal_2943, sbox_inst_5_n14}), .c ({output0_s2[125], output0_s1[125], output0_s0[125]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U8 ( .a ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, sbox_inst_5_n13}), .b ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, sbox_inst_5_n12}), .c ({new_AGEMA_signal_2944, new_AGEMA_signal_2943, sbox_inst_5_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_U7 ( .a ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, sbox_inst_5_T6}), .b ({input0_s2[23], input0_s1[23], input0_s0[23]}), .c ({new_AGEMA_signal_2610, new_AGEMA_signal_2609, sbox_inst_5_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_t5_AND_U1 ( .a ({input0_s2[21], input0_s1[21], input0_s0[21]}), .b ({new_AGEMA_signal_1788, new_AGEMA_signal_1787, sbox_inst_5_T3}), .clk (clk), .r ({Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, sbox_inst_5_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_5_t6_AND_U1 ( .a ({new_AGEMA_signal_1776, new_AGEMA_signal_1775, sbox_inst_5_L0}), .b ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, sbox_inst_5_T1}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807]}), .c ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, sbox_inst_5_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U15 ( .a ({new_AGEMA_signal_1806, new_AGEMA_signal_1805, sbox_inst_4_T2}), .b ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, sbox_inst_4_n20}), .c ({output0_s2[44], output0_s1[44], output0_s0[44]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U14 ( .a ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, sbox_inst_4_n19}), .b ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, sbox_inst_4_n18}), .c ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, sbox_inst_4_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U13 ( .a ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, sbox_inst_4_T1}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, sbox_inst_4_T5}), .c ({new_AGEMA_signal_2614, new_AGEMA_signal_2613, sbox_inst_4_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U11 ( .a ({input0_s2[17], input0_s1[17], input0_s0[17]}), .b ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, sbox_inst_4_n16}), .c ({output0_s2[84], output0_s1[84], output0_s0[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U10 ( .a ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, sbox_inst_4_n15}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, sbox_inst_4_T5}), .c ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, sbox_inst_4_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U9 ( .a ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, sbox_inst_4_n15}), .b ({new_AGEMA_signal_2952, new_AGEMA_signal_2951, sbox_inst_4_n14}), .c ({output0_s2[124], output0_s1[124], output0_s0[124]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U8 ( .a ({new_AGEMA_signal_2208, new_AGEMA_signal_2207, sbox_inst_4_n13}), .b ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, sbox_inst_4_n12}), .c ({new_AGEMA_signal_2952, new_AGEMA_signal_2951, sbox_inst_4_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_U7 ( .a ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, sbox_inst_4_T6}), .b ({input0_s2[19], input0_s1[19], input0_s0[19]}), .c ({new_AGEMA_signal_2620, new_AGEMA_signal_2619, sbox_inst_4_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_t5_AND_U1 ( .a ({input0_s2[17], input0_s1[17], input0_s0[17]}), .b ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, sbox_inst_4_T3}), .clk (clk), .r ({Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_2214, new_AGEMA_signal_2213, sbox_inst_4_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_4_t6_AND_U1 ( .a ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, sbox_inst_4_L0}), .b ({new_AGEMA_signal_1804, new_AGEMA_signal_1803, sbox_inst_4_T1}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813]}), .c ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, sbox_inst_4_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U15 ( .a ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, sbox_inst_3_T2}), .b ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, sbox_inst_3_n20}), .c ({output0_s2[43], output0_s1[43], output0_s0[43]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U14 ( .a ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, sbox_inst_3_n19}), .b ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, sbox_inst_3_n18}), .c ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, sbox_inst_3_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U13 ( .a ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, sbox_inst_3_T1}), .b ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, sbox_inst_3_T5}), .c ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, sbox_inst_3_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U11 ( .a ({input0_s2[13], input0_s1[13], input0_s0[13]}), .b ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, sbox_inst_3_n16}), .c ({output0_s2[83], output0_s1[83], output0_s0[83]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U10 ( .a ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, sbox_inst_3_n15}), .b ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, sbox_inst_3_T5}), .c ({new_AGEMA_signal_2628, new_AGEMA_signal_2627, sbox_inst_3_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U9 ( .a ({new_AGEMA_signal_2220, new_AGEMA_signal_2219, sbox_inst_3_n15}), .b ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, sbox_inst_3_n14}), .c ({output0_s2[123], output0_s1[123], output0_s0[123]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U8 ( .a ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, sbox_inst_3_n13}), .b ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, sbox_inst_3_n12}), .c ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, sbox_inst_3_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_U7 ( .a ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, sbox_inst_3_T6}), .b ({input0_s2[15], input0_s1[15], input0_s0[15]}), .c ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, sbox_inst_3_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_t5_AND_U1 ( .a ({input0_s2[13], input0_s1[13], input0_s0[13]}), .b ({new_AGEMA_signal_1828, new_AGEMA_signal_1827, sbox_inst_3_T3}), .clk (clk), .r ({Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, sbox_inst_3_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_3_t6_AND_U1 ( .a ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, sbox_inst_3_L0}), .b ({new_AGEMA_signal_1824, new_AGEMA_signal_1823, sbox_inst_3_T1}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819]}), .c ({new_AGEMA_signal_2226, new_AGEMA_signal_2225, sbox_inst_3_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U15 ( .a ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, sbox_inst_2_T2}), .b ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, sbox_inst_2_n20}), .c ({output0_s2[42], output0_s1[42], output0_s0[42]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U14 ( .a ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, sbox_inst_2_n19}), .b ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, sbox_inst_2_n18}), .c ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, sbox_inst_2_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U13 ( .a ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, sbox_inst_2_T1}), .b ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, sbox_inst_2_T5}), .c ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, sbox_inst_2_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U11 ( .a ({input0_s2[9], input0_s1[9], input0_s0[9]}), .b ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, sbox_inst_2_n16}), .c ({output0_s2[82], output0_s1[82], output0_s0[82]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U10 ( .a ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, sbox_inst_2_n15}), .b ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, sbox_inst_2_T5}), .c ({new_AGEMA_signal_2638, new_AGEMA_signal_2637, sbox_inst_2_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U9 ( .a ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, sbox_inst_2_n15}), .b ({new_AGEMA_signal_2968, new_AGEMA_signal_2967, sbox_inst_2_n14}), .c ({output0_s2[122], output0_s1[122], output0_s0[122]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U8 ( .a ({new_AGEMA_signal_2228, new_AGEMA_signal_2227, sbox_inst_2_n13}), .b ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, sbox_inst_2_n12}), .c ({new_AGEMA_signal_2968, new_AGEMA_signal_2967, sbox_inst_2_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_U7 ( .a ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, sbox_inst_2_T6}), .b ({input0_s2[11], input0_s1[11], input0_s0[11]}), .c ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, sbox_inst_2_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_t5_AND_U1 ( .a ({input0_s2[9], input0_s1[9], input0_s0[9]}), .b ({new_AGEMA_signal_1848, new_AGEMA_signal_1847, sbox_inst_2_T3}), .clk (clk), .r ({Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, sbox_inst_2_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_2_t6_AND_U1 ( .a ({new_AGEMA_signal_1836, new_AGEMA_signal_1835, sbox_inst_2_L0}), .b ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, sbox_inst_2_T1}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825]}), .c ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, sbox_inst_2_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U15 ( .a ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, sbox_inst_1_T2}), .b ({new_AGEMA_signal_3152, new_AGEMA_signal_3151, sbox_inst_1_n20}), .c ({output0_s2[41], output0_s1[41], output0_s0[41]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U14 ( .a ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, sbox_inst_1_n19}), .b ({new_AGEMA_signal_2972, new_AGEMA_signal_2971, sbox_inst_1_n18}), .c ({new_AGEMA_signal_3152, new_AGEMA_signal_3151, sbox_inst_1_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U13 ( .a ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, sbox_inst_1_T1}), .b ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, sbox_inst_1_T5}), .c ({new_AGEMA_signal_2972, new_AGEMA_signal_2971, sbox_inst_1_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U11 ( .a ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, input_array_5}), .b ({new_AGEMA_signal_2976, new_AGEMA_signal_2975, sbox_inst_1_n16}), .c ({output0_s2[81], output0_s1[81], output0_s0[81]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U10 ( .a ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, sbox_inst_1_n15}), .b ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, sbox_inst_1_T5}), .c ({new_AGEMA_signal_2976, new_AGEMA_signal_2975, sbox_inst_1_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U9 ( .a ({new_AGEMA_signal_2646, new_AGEMA_signal_2645, sbox_inst_1_n15}), .b ({new_AGEMA_signal_3156, new_AGEMA_signal_3155, sbox_inst_1_n14}), .c ({output0_s2[121], output0_s1[121], output0_s0[121]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U8 ( .a ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, sbox_inst_1_n13}), .b ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, sbox_inst_1_n12}), .c ({new_AGEMA_signal_3156, new_AGEMA_signal_3155, sbox_inst_1_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_U7 ( .a ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, sbox_inst_1_T6}), .b ({input0_s2[7], input0_s1[7], input0_s0[7]}), .c ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, sbox_inst_1_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_t5_AND_U1 ( .a ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, input_array_5}), .b ({new_AGEMA_signal_2248, new_AGEMA_signal_2247, sbox_inst_1_T3}), .clk (clk), .r ({Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_2650, new_AGEMA_signal_2649, sbox_inst_1_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_1_t6_AND_U1 ( .a ({new_AGEMA_signal_2238, new_AGEMA_signal_2237, sbox_inst_1_L0}), .b ({new_AGEMA_signal_2244, new_AGEMA_signal_2243, sbox_inst_1_T1}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831]}), .c ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, sbox_inst_1_T6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U15 ( .a ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, sbox_inst_0_T2}), .b ({new_AGEMA_signal_3160, new_AGEMA_signal_3159, sbox_inst_0_n20}), .c ({output0_s2[40], output0_s1[40], output0_s0[40]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U14 ( .a ({new_AGEMA_signal_2984, new_AGEMA_signal_2983, sbox_inst_0_n19}), .b ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, sbox_inst_0_n18}), .c ({new_AGEMA_signal_3160, new_AGEMA_signal_3159, sbox_inst_0_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U13 ( .a ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, sbox_inst_0_T1}), .b ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, sbox_inst_0_T5}), .c ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, sbox_inst_0_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U11 ( .a ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, input_array_1}), .b ({new_AGEMA_signal_2986, new_AGEMA_signal_2985, sbox_inst_0_n16}), .c ({output0_s2[80], output0_s1[80], output0_s0[80]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U10 ( .a ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, sbox_inst_0_n15}), .b ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, sbox_inst_0_T5}), .c ({new_AGEMA_signal_2986, new_AGEMA_signal_2985, sbox_inst_0_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U9 ( .a ({new_AGEMA_signal_2656, new_AGEMA_signal_2655, sbox_inst_0_n15}), .b ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, sbox_inst_0_n14}), .c ({output0_s2[120], output0_s1[120], output0_s0[120]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U8 ( .a ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, sbox_inst_0_n13}), .b ({new_AGEMA_signal_2988, new_AGEMA_signal_2987, sbox_inst_0_n12}), .c ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, sbox_inst_0_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_U7 ( .a ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, sbox_inst_0_T6}), .b ({new_AGEMA_signal_1102, new_AGEMA_signal_1101, input_array_3}), .c ({new_AGEMA_signal_2988, new_AGEMA_signal_2987, sbox_inst_0_n12}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_t5_AND_U1 ( .a ({new_AGEMA_signal_1078, new_AGEMA_signal_1077, input_array_1}), .b ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, sbox_inst_0_T3}), .clk (clk), .r ({Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, sbox_inst_0_T5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) sbox_inst_0_t6_AND_U1 ( .a ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, sbox_inst_0_L0}), .b ({new_AGEMA_signal_2256, new_AGEMA_signal_2255, sbox_inst_0_T1}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837]}), .c ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, sbox_inst_0_T6}) ) ;

endmodule
