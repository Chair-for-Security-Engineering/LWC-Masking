/* modified netlist. Source: module Photon_256 in file ./test/Photon_256.v */
/* clock gating is added to the circuit, the latency increased 6 time(s)  */

module Photon_256_HPC2_ClockGating_d3 (w0_s0, w1_s0, temp_s0, k, p256_sel, clk, w0_s1, w0_s2, w0_s3, w1_s1, w1_s2, w1_s3, temp_s1, temp_s2, temp_s3, Fresh, /*rst,*/ y0_s0, y1_s0, temp_next_s0, temp_next_s1, temp_next_s2, temp_next_s3, y0_s1, y0_s2, y0_s3, y1_s1, y1_s2, y1_s3/*, Synch*/);
    input [127:0] w0_s0 ;
    input [127:0] w1_s0 ;
    input [127:0] temp_s0 ;
    input [3:0] k ;
    input p256_sel ;
    input clk ;
    input [127:0] w0_s1 ;
    input [127:0] w0_s2 ;
    input [127:0] w0_s3 ;
    input [127:0] w1_s1 ;
    input [127:0] w1_s2 ;
    input [127:0] w1_s3 ;
    input [127:0] temp_s1 ;
    input [127:0] temp_s2 ;
    input [127:0] temp_s3 ;
    //input rst ;
    input [6719:0] Fresh ;
    output [127:0] y0_s0 ;
    output [127:0] y1_s0 ;
    output [127:0] temp_next_s0 ;
    output [127:0] temp_next_s1 ;
    output [127:0] temp_next_s2 ;
    output [127:0] temp_next_s3 ;
    output [127:0] y0_s1 ;
    output [127:0] y0_s2 ;
    output [127:0] y0_s3 ;
    output [127:0] y1_s1 ;
    output [127:0] y1_s2 ;
    output [127:0] y1_s3 ;
    //output Synch ;
    wire add_sub1_0_n8 ;
    wire add_sub1_0_n7 ;
    wire add_sub1_0_n6 ;
    wire add_sub1_0_n5 ;
    wire add_sub1_0_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_0_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_0_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_0_subc_rom_sbox_0_ANF_2_t0 ;
    wire add_sub1_1_n8 ;
    wire add_sub1_1_n7 ;
    wire add_sub1_1_n6 ;
    wire add_sub1_1_n5 ;
    wire add_sub1_1_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_1_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_1_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_1_subc_rom_sbox_0_ANF_2_t0 ;
    wire add_sub1_2_n8 ;
    wire add_sub1_2_n7 ;
    wire add_sub1_2_n6 ;
    wire add_sub1_2_n5 ;
    wire add_sub1_2_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_2_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_2_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_2_subc_rom_sbox_0_ANF_2_t0 ;
    wire add_sub1_3_n8 ;
    wire add_sub1_3_n7 ;
    wire add_sub1_3_n6 ;
    wire add_sub1_3_n5 ;
    wire add_sub1_3_addc_rom_ic_out_0_ ;
    wire add_sub1_3_addc_rom_ic_out_1_ ;
    wire add_sub1_3_addc_rom_ic_out_2_ ;
    wire add_sub1_3_addc_rom_ic1_ANF_0_n2 ;
    wire add_sub1_3_addc_rom_ic1_ANF_0_t0 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n21 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n20 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n19 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n18 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n17 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n16 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n15 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n14 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n13 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_n12 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t7 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t6 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t5 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t4 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t3 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t2 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t1 ;
    wire add_sub1_3_addc_rom_rc1_ANF_1_t0 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_7_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_6_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_5_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_4_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_3_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_2_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_1_ANF_2_t0 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n20 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n19 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n18 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n17 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n16 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n15 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n14 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n13 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_n12 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t7 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t6 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t5 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t4 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t3 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t2 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t1 ;
    wire add_sub1_3_subc_rom_sbox_0_ANF_2_t0 ;
    wire mcs1_mcs_mat1_0_n128 ;
    wire mcs1_mcs_mat1_0_n127 ;
    wire mcs1_mcs_mat1_0_n126 ;
    wire mcs1_mcs_mat1_0_n125 ;
    wire mcs1_mcs_mat1_0_n124 ;
    wire mcs1_mcs_mat1_0_n123 ;
    wire mcs1_mcs_mat1_0_n122 ;
    wire mcs1_mcs_mat1_0_n121 ;
    wire mcs1_mcs_mat1_0_n120 ;
    wire mcs1_mcs_mat1_0_n119 ;
    wire mcs1_mcs_mat1_0_n118 ;
    wire mcs1_mcs_mat1_0_n117 ;
    wire mcs1_mcs_mat1_0_n116 ;
    wire mcs1_mcs_mat1_0_n115 ;
    wire mcs1_mcs_mat1_0_n114 ;
    wire mcs1_mcs_mat1_0_n113 ;
    wire mcs1_mcs_mat1_0_n112 ;
    wire mcs1_mcs_mat1_0_n111 ;
    wire mcs1_mcs_mat1_0_n110 ;
    wire mcs1_mcs_mat1_0_n109 ;
    wire mcs1_mcs_mat1_0_n108 ;
    wire mcs1_mcs_mat1_0_n107 ;
    wire mcs1_mcs_mat1_0_n106 ;
    wire mcs1_mcs_mat1_0_n105 ;
    wire mcs1_mcs_mat1_0_n104 ;
    wire mcs1_mcs_mat1_0_n103 ;
    wire mcs1_mcs_mat1_0_n102 ;
    wire mcs1_mcs_mat1_0_n101 ;
    wire mcs1_mcs_mat1_0_n100 ;
    wire mcs1_mcs_mat1_0_n99 ;
    wire mcs1_mcs_mat1_0_n98 ;
    wire mcs1_mcs_mat1_0_n97 ;
    wire mcs1_mcs_mat1_0_n96 ;
    wire mcs1_mcs_mat1_0_n95 ;
    wire mcs1_mcs_mat1_0_n94 ;
    wire mcs1_mcs_mat1_0_n93 ;
    wire mcs1_mcs_mat1_0_n92 ;
    wire mcs1_mcs_mat1_0_n91 ;
    wire mcs1_mcs_mat1_0_n90 ;
    wire mcs1_mcs_mat1_0_n89 ;
    wire mcs1_mcs_mat1_0_n88 ;
    wire mcs1_mcs_mat1_0_n87 ;
    wire mcs1_mcs_mat1_0_n86 ;
    wire mcs1_mcs_mat1_0_n85 ;
    wire mcs1_mcs_mat1_0_n84 ;
    wire mcs1_mcs_mat1_0_n83 ;
    wire mcs1_mcs_mat1_0_n82 ;
    wire mcs1_mcs_mat1_0_n81 ;
    wire mcs1_mcs_mat1_0_n80 ;
    wire mcs1_mcs_mat1_0_n79 ;
    wire mcs1_mcs_mat1_0_n78 ;
    wire mcs1_mcs_mat1_0_n77 ;
    wire mcs1_mcs_mat1_0_n76 ;
    wire mcs1_mcs_mat1_0_n75 ;
    wire mcs1_mcs_mat1_0_n74 ;
    wire mcs1_mcs_mat1_0_n73 ;
    wire mcs1_mcs_mat1_0_n72 ;
    wire mcs1_mcs_mat1_0_n71 ;
    wire mcs1_mcs_mat1_0_n70 ;
    wire mcs1_mcs_mat1_0_n69 ;
    wire mcs1_mcs_mat1_0_n68 ;
    wire mcs1_mcs_mat1_0_n67 ;
    wire mcs1_mcs_mat1_0_n66 ;
    wire mcs1_mcs_mat1_0_n65 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_0_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_1_n128 ;
    wire mcs1_mcs_mat1_1_n127 ;
    wire mcs1_mcs_mat1_1_n126 ;
    wire mcs1_mcs_mat1_1_n125 ;
    wire mcs1_mcs_mat1_1_n124 ;
    wire mcs1_mcs_mat1_1_n123 ;
    wire mcs1_mcs_mat1_1_n122 ;
    wire mcs1_mcs_mat1_1_n121 ;
    wire mcs1_mcs_mat1_1_n120 ;
    wire mcs1_mcs_mat1_1_n119 ;
    wire mcs1_mcs_mat1_1_n118 ;
    wire mcs1_mcs_mat1_1_n117 ;
    wire mcs1_mcs_mat1_1_n116 ;
    wire mcs1_mcs_mat1_1_n115 ;
    wire mcs1_mcs_mat1_1_n114 ;
    wire mcs1_mcs_mat1_1_n113 ;
    wire mcs1_mcs_mat1_1_n112 ;
    wire mcs1_mcs_mat1_1_n111 ;
    wire mcs1_mcs_mat1_1_n110 ;
    wire mcs1_mcs_mat1_1_n109 ;
    wire mcs1_mcs_mat1_1_n108 ;
    wire mcs1_mcs_mat1_1_n107 ;
    wire mcs1_mcs_mat1_1_n106 ;
    wire mcs1_mcs_mat1_1_n105 ;
    wire mcs1_mcs_mat1_1_n104 ;
    wire mcs1_mcs_mat1_1_n103 ;
    wire mcs1_mcs_mat1_1_n102 ;
    wire mcs1_mcs_mat1_1_n101 ;
    wire mcs1_mcs_mat1_1_n100 ;
    wire mcs1_mcs_mat1_1_n99 ;
    wire mcs1_mcs_mat1_1_n98 ;
    wire mcs1_mcs_mat1_1_n97 ;
    wire mcs1_mcs_mat1_1_n96 ;
    wire mcs1_mcs_mat1_1_n95 ;
    wire mcs1_mcs_mat1_1_n94 ;
    wire mcs1_mcs_mat1_1_n93 ;
    wire mcs1_mcs_mat1_1_n92 ;
    wire mcs1_mcs_mat1_1_n91 ;
    wire mcs1_mcs_mat1_1_n90 ;
    wire mcs1_mcs_mat1_1_n89 ;
    wire mcs1_mcs_mat1_1_n88 ;
    wire mcs1_mcs_mat1_1_n87 ;
    wire mcs1_mcs_mat1_1_n86 ;
    wire mcs1_mcs_mat1_1_n85 ;
    wire mcs1_mcs_mat1_1_n84 ;
    wire mcs1_mcs_mat1_1_n83 ;
    wire mcs1_mcs_mat1_1_n82 ;
    wire mcs1_mcs_mat1_1_n81 ;
    wire mcs1_mcs_mat1_1_n80 ;
    wire mcs1_mcs_mat1_1_n79 ;
    wire mcs1_mcs_mat1_1_n78 ;
    wire mcs1_mcs_mat1_1_n77 ;
    wire mcs1_mcs_mat1_1_n76 ;
    wire mcs1_mcs_mat1_1_n75 ;
    wire mcs1_mcs_mat1_1_n74 ;
    wire mcs1_mcs_mat1_1_n73 ;
    wire mcs1_mcs_mat1_1_n72 ;
    wire mcs1_mcs_mat1_1_n71 ;
    wire mcs1_mcs_mat1_1_n70 ;
    wire mcs1_mcs_mat1_1_n69 ;
    wire mcs1_mcs_mat1_1_n68 ;
    wire mcs1_mcs_mat1_1_n67 ;
    wire mcs1_mcs_mat1_1_n66 ;
    wire mcs1_mcs_mat1_1_n65 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_1_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_2_n128 ;
    wire mcs1_mcs_mat1_2_n127 ;
    wire mcs1_mcs_mat1_2_n126 ;
    wire mcs1_mcs_mat1_2_n125 ;
    wire mcs1_mcs_mat1_2_n124 ;
    wire mcs1_mcs_mat1_2_n123 ;
    wire mcs1_mcs_mat1_2_n122 ;
    wire mcs1_mcs_mat1_2_n121 ;
    wire mcs1_mcs_mat1_2_n120 ;
    wire mcs1_mcs_mat1_2_n119 ;
    wire mcs1_mcs_mat1_2_n118 ;
    wire mcs1_mcs_mat1_2_n117 ;
    wire mcs1_mcs_mat1_2_n116 ;
    wire mcs1_mcs_mat1_2_n115 ;
    wire mcs1_mcs_mat1_2_n114 ;
    wire mcs1_mcs_mat1_2_n113 ;
    wire mcs1_mcs_mat1_2_n112 ;
    wire mcs1_mcs_mat1_2_n111 ;
    wire mcs1_mcs_mat1_2_n110 ;
    wire mcs1_mcs_mat1_2_n109 ;
    wire mcs1_mcs_mat1_2_n108 ;
    wire mcs1_mcs_mat1_2_n107 ;
    wire mcs1_mcs_mat1_2_n106 ;
    wire mcs1_mcs_mat1_2_n105 ;
    wire mcs1_mcs_mat1_2_n104 ;
    wire mcs1_mcs_mat1_2_n103 ;
    wire mcs1_mcs_mat1_2_n102 ;
    wire mcs1_mcs_mat1_2_n101 ;
    wire mcs1_mcs_mat1_2_n100 ;
    wire mcs1_mcs_mat1_2_n99 ;
    wire mcs1_mcs_mat1_2_n98 ;
    wire mcs1_mcs_mat1_2_n97 ;
    wire mcs1_mcs_mat1_2_n96 ;
    wire mcs1_mcs_mat1_2_n95 ;
    wire mcs1_mcs_mat1_2_n94 ;
    wire mcs1_mcs_mat1_2_n93 ;
    wire mcs1_mcs_mat1_2_n92 ;
    wire mcs1_mcs_mat1_2_n91 ;
    wire mcs1_mcs_mat1_2_n90 ;
    wire mcs1_mcs_mat1_2_n89 ;
    wire mcs1_mcs_mat1_2_n88 ;
    wire mcs1_mcs_mat1_2_n87 ;
    wire mcs1_mcs_mat1_2_n86 ;
    wire mcs1_mcs_mat1_2_n85 ;
    wire mcs1_mcs_mat1_2_n84 ;
    wire mcs1_mcs_mat1_2_n83 ;
    wire mcs1_mcs_mat1_2_n82 ;
    wire mcs1_mcs_mat1_2_n81 ;
    wire mcs1_mcs_mat1_2_n80 ;
    wire mcs1_mcs_mat1_2_n79 ;
    wire mcs1_mcs_mat1_2_n78 ;
    wire mcs1_mcs_mat1_2_n77 ;
    wire mcs1_mcs_mat1_2_n76 ;
    wire mcs1_mcs_mat1_2_n75 ;
    wire mcs1_mcs_mat1_2_n74 ;
    wire mcs1_mcs_mat1_2_n73 ;
    wire mcs1_mcs_mat1_2_n72 ;
    wire mcs1_mcs_mat1_2_n71 ;
    wire mcs1_mcs_mat1_2_n70 ;
    wire mcs1_mcs_mat1_2_n69 ;
    wire mcs1_mcs_mat1_2_n68 ;
    wire mcs1_mcs_mat1_2_n67 ;
    wire mcs1_mcs_mat1_2_n66 ;
    wire mcs1_mcs_mat1_2_n65 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_2_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_3_n128 ;
    wire mcs1_mcs_mat1_3_n127 ;
    wire mcs1_mcs_mat1_3_n126 ;
    wire mcs1_mcs_mat1_3_n125 ;
    wire mcs1_mcs_mat1_3_n124 ;
    wire mcs1_mcs_mat1_3_n123 ;
    wire mcs1_mcs_mat1_3_n122 ;
    wire mcs1_mcs_mat1_3_n121 ;
    wire mcs1_mcs_mat1_3_n120 ;
    wire mcs1_mcs_mat1_3_n119 ;
    wire mcs1_mcs_mat1_3_n118 ;
    wire mcs1_mcs_mat1_3_n117 ;
    wire mcs1_mcs_mat1_3_n116 ;
    wire mcs1_mcs_mat1_3_n115 ;
    wire mcs1_mcs_mat1_3_n114 ;
    wire mcs1_mcs_mat1_3_n113 ;
    wire mcs1_mcs_mat1_3_n112 ;
    wire mcs1_mcs_mat1_3_n111 ;
    wire mcs1_mcs_mat1_3_n110 ;
    wire mcs1_mcs_mat1_3_n109 ;
    wire mcs1_mcs_mat1_3_n108 ;
    wire mcs1_mcs_mat1_3_n107 ;
    wire mcs1_mcs_mat1_3_n106 ;
    wire mcs1_mcs_mat1_3_n105 ;
    wire mcs1_mcs_mat1_3_n104 ;
    wire mcs1_mcs_mat1_3_n103 ;
    wire mcs1_mcs_mat1_3_n102 ;
    wire mcs1_mcs_mat1_3_n101 ;
    wire mcs1_mcs_mat1_3_n100 ;
    wire mcs1_mcs_mat1_3_n99 ;
    wire mcs1_mcs_mat1_3_n98 ;
    wire mcs1_mcs_mat1_3_n97 ;
    wire mcs1_mcs_mat1_3_n96 ;
    wire mcs1_mcs_mat1_3_n95 ;
    wire mcs1_mcs_mat1_3_n94 ;
    wire mcs1_mcs_mat1_3_n93 ;
    wire mcs1_mcs_mat1_3_n92 ;
    wire mcs1_mcs_mat1_3_n91 ;
    wire mcs1_mcs_mat1_3_n90 ;
    wire mcs1_mcs_mat1_3_n89 ;
    wire mcs1_mcs_mat1_3_n88 ;
    wire mcs1_mcs_mat1_3_n87 ;
    wire mcs1_mcs_mat1_3_n86 ;
    wire mcs1_mcs_mat1_3_n85 ;
    wire mcs1_mcs_mat1_3_n84 ;
    wire mcs1_mcs_mat1_3_n83 ;
    wire mcs1_mcs_mat1_3_n82 ;
    wire mcs1_mcs_mat1_3_n81 ;
    wire mcs1_mcs_mat1_3_n80 ;
    wire mcs1_mcs_mat1_3_n79 ;
    wire mcs1_mcs_mat1_3_n78 ;
    wire mcs1_mcs_mat1_3_n77 ;
    wire mcs1_mcs_mat1_3_n76 ;
    wire mcs1_mcs_mat1_3_n75 ;
    wire mcs1_mcs_mat1_3_n74 ;
    wire mcs1_mcs_mat1_3_n73 ;
    wire mcs1_mcs_mat1_3_n72 ;
    wire mcs1_mcs_mat1_3_n71 ;
    wire mcs1_mcs_mat1_3_n70 ;
    wire mcs1_mcs_mat1_3_n69 ;
    wire mcs1_mcs_mat1_3_n68 ;
    wire mcs1_mcs_mat1_3_n67 ;
    wire mcs1_mcs_mat1_3_n66 ;
    wire mcs1_mcs_mat1_3_n65 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_3_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_4_n128 ;
    wire mcs1_mcs_mat1_4_n127 ;
    wire mcs1_mcs_mat1_4_n126 ;
    wire mcs1_mcs_mat1_4_n125 ;
    wire mcs1_mcs_mat1_4_n124 ;
    wire mcs1_mcs_mat1_4_n123 ;
    wire mcs1_mcs_mat1_4_n122 ;
    wire mcs1_mcs_mat1_4_n121 ;
    wire mcs1_mcs_mat1_4_n120 ;
    wire mcs1_mcs_mat1_4_n119 ;
    wire mcs1_mcs_mat1_4_n118 ;
    wire mcs1_mcs_mat1_4_n117 ;
    wire mcs1_mcs_mat1_4_n116 ;
    wire mcs1_mcs_mat1_4_n115 ;
    wire mcs1_mcs_mat1_4_n114 ;
    wire mcs1_mcs_mat1_4_n113 ;
    wire mcs1_mcs_mat1_4_n112 ;
    wire mcs1_mcs_mat1_4_n111 ;
    wire mcs1_mcs_mat1_4_n110 ;
    wire mcs1_mcs_mat1_4_n109 ;
    wire mcs1_mcs_mat1_4_n108 ;
    wire mcs1_mcs_mat1_4_n107 ;
    wire mcs1_mcs_mat1_4_n106 ;
    wire mcs1_mcs_mat1_4_n105 ;
    wire mcs1_mcs_mat1_4_n104 ;
    wire mcs1_mcs_mat1_4_n103 ;
    wire mcs1_mcs_mat1_4_n102 ;
    wire mcs1_mcs_mat1_4_n101 ;
    wire mcs1_mcs_mat1_4_n100 ;
    wire mcs1_mcs_mat1_4_n99 ;
    wire mcs1_mcs_mat1_4_n98 ;
    wire mcs1_mcs_mat1_4_n97 ;
    wire mcs1_mcs_mat1_4_n96 ;
    wire mcs1_mcs_mat1_4_n95 ;
    wire mcs1_mcs_mat1_4_n94 ;
    wire mcs1_mcs_mat1_4_n93 ;
    wire mcs1_mcs_mat1_4_n92 ;
    wire mcs1_mcs_mat1_4_n91 ;
    wire mcs1_mcs_mat1_4_n90 ;
    wire mcs1_mcs_mat1_4_n89 ;
    wire mcs1_mcs_mat1_4_n88 ;
    wire mcs1_mcs_mat1_4_n87 ;
    wire mcs1_mcs_mat1_4_n86 ;
    wire mcs1_mcs_mat1_4_n85 ;
    wire mcs1_mcs_mat1_4_n84 ;
    wire mcs1_mcs_mat1_4_n83 ;
    wire mcs1_mcs_mat1_4_n82 ;
    wire mcs1_mcs_mat1_4_n81 ;
    wire mcs1_mcs_mat1_4_n80 ;
    wire mcs1_mcs_mat1_4_n79 ;
    wire mcs1_mcs_mat1_4_n78 ;
    wire mcs1_mcs_mat1_4_n77 ;
    wire mcs1_mcs_mat1_4_n76 ;
    wire mcs1_mcs_mat1_4_n75 ;
    wire mcs1_mcs_mat1_4_n74 ;
    wire mcs1_mcs_mat1_4_n73 ;
    wire mcs1_mcs_mat1_4_n72 ;
    wire mcs1_mcs_mat1_4_n71 ;
    wire mcs1_mcs_mat1_4_n70 ;
    wire mcs1_mcs_mat1_4_n69 ;
    wire mcs1_mcs_mat1_4_n68 ;
    wire mcs1_mcs_mat1_4_n67 ;
    wire mcs1_mcs_mat1_4_n66 ;
    wire mcs1_mcs_mat1_4_n65 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_4_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_5_n128 ;
    wire mcs1_mcs_mat1_5_n127 ;
    wire mcs1_mcs_mat1_5_n126 ;
    wire mcs1_mcs_mat1_5_n125 ;
    wire mcs1_mcs_mat1_5_n124 ;
    wire mcs1_mcs_mat1_5_n123 ;
    wire mcs1_mcs_mat1_5_n122 ;
    wire mcs1_mcs_mat1_5_n121 ;
    wire mcs1_mcs_mat1_5_n120 ;
    wire mcs1_mcs_mat1_5_n119 ;
    wire mcs1_mcs_mat1_5_n118 ;
    wire mcs1_mcs_mat1_5_n117 ;
    wire mcs1_mcs_mat1_5_n116 ;
    wire mcs1_mcs_mat1_5_n115 ;
    wire mcs1_mcs_mat1_5_n114 ;
    wire mcs1_mcs_mat1_5_n113 ;
    wire mcs1_mcs_mat1_5_n112 ;
    wire mcs1_mcs_mat1_5_n111 ;
    wire mcs1_mcs_mat1_5_n110 ;
    wire mcs1_mcs_mat1_5_n109 ;
    wire mcs1_mcs_mat1_5_n108 ;
    wire mcs1_mcs_mat1_5_n107 ;
    wire mcs1_mcs_mat1_5_n106 ;
    wire mcs1_mcs_mat1_5_n105 ;
    wire mcs1_mcs_mat1_5_n104 ;
    wire mcs1_mcs_mat1_5_n103 ;
    wire mcs1_mcs_mat1_5_n102 ;
    wire mcs1_mcs_mat1_5_n101 ;
    wire mcs1_mcs_mat1_5_n100 ;
    wire mcs1_mcs_mat1_5_n99 ;
    wire mcs1_mcs_mat1_5_n98 ;
    wire mcs1_mcs_mat1_5_n97 ;
    wire mcs1_mcs_mat1_5_n96 ;
    wire mcs1_mcs_mat1_5_n95 ;
    wire mcs1_mcs_mat1_5_n94 ;
    wire mcs1_mcs_mat1_5_n93 ;
    wire mcs1_mcs_mat1_5_n92 ;
    wire mcs1_mcs_mat1_5_n91 ;
    wire mcs1_mcs_mat1_5_n90 ;
    wire mcs1_mcs_mat1_5_n89 ;
    wire mcs1_mcs_mat1_5_n88 ;
    wire mcs1_mcs_mat1_5_n87 ;
    wire mcs1_mcs_mat1_5_n86 ;
    wire mcs1_mcs_mat1_5_n85 ;
    wire mcs1_mcs_mat1_5_n84 ;
    wire mcs1_mcs_mat1_5_n83 ;
    wire mcs1_mcs_mat1_5_n82 ;
    wire mcs1_mcs_mat1_5_n81 ;
    wire mcs1_mcs_mat1_5_n80 ;
    wire mcs1_mcs_mat1_5_n79 ;
    wire mcs1_mcs_mat1_5_n78 ;
    wire mcs1_mcs_mat1_5_n77 ;
    wire mcs1_mcs_mat1_5_n76 ;
    wire mcs1_mcs_mat1_5_n75 ;
    wire mcs1_mcs_mat1_5_n74 ;
    wire mcs1_mcs_mat1_5_n73 ;
    wire mcs1_mcs_mat1_5_n72 ;
    wire mcs1_mcs_mat1_5_n71 ;
    wire mcs1_mcs_mat1_5_n70 ;
    wire mcs1_mcs_mat1_5_n69 ;
    wire mcs1_mcs_mat1_5_n68 ;
    wire mcs1_mcs_mat1_5_n67 ;
    wire mcs1_mcs_mat1_5_n66 ;
    wire mcs1_mcs_mat1_5_n65 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_5_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_6_n128 ;
    wire mcs1_mcs_mat1_6_n127 ;
    wire mcs1_mcs_mat1_6_n126 ;
    wire mcs1_mcs_mat1_6_n125 ;
    wire mcs1_mcs_mat1_6_n124 ;
    wire mcs1_mcs_mat1_6_n123 ;
    wire mcs1_mcs_mat1_6_n122 ;
    wire mcs1_mcs_mat1_6_n121 ;
    wire mcs1_mcs_mat1_6_n120 ;
    wire mcs1_mcs_mat1_6_n119 ;
    wire mcs1_mcs_mat1_6_n118 ;
    wire mcs1_mcs_mat1_6_n117 ;
    wire mcs1_mcs_mat1_6_n116 ;
    wire mcs1_mcs_mat1_6_n115 ;
    wire mcs1_mcs_mat1_6_n114 ;
    wire mcs1_mcs_mat1_6_n113 ;
    wire mcs1_mcs_mat1_6_n112 ;
    wire mcs1_mcs_mat1_6_n111 ;
    wire mcs1_mcs_mat1_6_n110 ;
    wire mcs1_mcs_mat1_6_n109 ;
    wire mcs1_mcs_mat1_6_n108 ;
    wire mcs1_mcs_mat1_6_n107 ;
    wire mcs1_mcs_mat1_6_n106 ;
    wire mcs1_mcs_mat1_6_n105 ;
    wire mcs1_mcs_mat1_6_n104 ;
    wire mcs1_mcs_mat1_6_n103 ;
    wire mcs1_mcs_mat1_6_n102 ;
    wire mcs1_mcs_mat1_6_n101 ;
    wire mcs1_mcs_mat1_6_n100 ;
    wire mcs1_mcs_mat1_6_n99 ;
    wire mcs1_mcs_mat1_6_n98 ;
    wire mcs1_mcs_mat1_6_n97 ;
    wire mcs1_mcs_mat1_6_n96 ;
    wire mcs1_mcs_mat1_6_n95 ;
    wire mcs1_mcs_mat1_6_n94 ;
    wire mcs1_mcs_mat1_6_n93 ;
    wire mcs1_mcs_mat1_6_n92 ;
    wire mcs1_mcs_mat1_6_n91 ;
    wire mcs1_mcs_mat1_6_n90 ;
    wire mcs1_mcs_mat1_6_n89 ;
    wire mcs1_mcs_mat1_6_n88 ;
    wire mcs1_mcs_mat1_6_n87 ;
    wire mcs1_mcs_mat1_6_n86 ;
    wire mcs1_mcs_mat1_6_n85 ;
    wire mcs1_mcs_mat1_6_n84 ;
    wire mcs1_mcs_mat1_6_n83 ;
    wire mcs1_mcs_mat1_6_n82 ;
    wire mcs1_mcs_mat1_6_n81 ;
    wire mcs1_mcs_mat1_6_n80 ;
    wire mcs1_mcs_mat1_6_n79 ;
    wire mcs1_mcs_mat1_6_n78 ;
    wire mcs1_mcs_mat1_6_n77 ;
    wire mcs1_mcs_mat1_6_n76 ;
    wire mcs1_mcs_mat1_6_n75 ;
    wire mcs1_mcs_mat1_6_n74 ;
    wire mcs1_mcs_mat1_6_n73 ;
    wire mcs1_mcs_mat1_6_n72 ;
    wire mcs1_mcs_mat1_6_n71 ;
    wire mcs1_mcs_mat1_6_n70 ;
    wire mcs1_mcs_mat1_6_n69 ;
    wire mcs1_mcs_mat1_6_n68 ;
    wire mcs1_mcs_mat1_6_n67 ;
    wire mcs1_mcs_mat1_6_n66 ;
    wire mcs1_mcs_mat1_6_n65 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_6_mcs_rom0_31_x0x4 ;
    wire mcs1_mcs_mat1_7_n128 ;
    wire mcs1_mcs_mat1_7_n127 ;
    wire mcs1_mcs_mat1_7_n126 ;
    wire mcs1_mcs_mat1_7_n125 ;
    wire mcs1_mcs_mat1_7_n124 ;
    wire mcs1_mcs_mat1_7_n123 ;
    wire mcs1_mcs_mat1_7_n122 ;
    wire mcs1_mcs_mat1_7_n121 ;
    wire mcs1_mcs_mat1_7_n120 ;
    wire mcs1_mcs_mat1_7_n119 ;
    wire mcs1_mcs_mat1_7_n118 ;
    wire mcs1_mcs_mat1_7_n117 ;
    wire mcs1_mcs_mat1_7_n116 ;
    wire mcs1_mcs_mat1_7_n115 ;
    wire mcs1_mcs_mat1_7_n114 ;
    wire mcs1_mcs_mat1_7_n113 ;
    wire mcs1_mcs_mat1_7_n112 ;
    wire mcs1_mcs_mat1_7_n111 ;
    wire mcs1_mcs_mat1_7_n110 ;
    wire mcs1_mcs_mat1_7_n109 ;
    wire mcs1_mcs_mat1_7_n108 ;
    wire mcs1_mcs_mat1_7_n107 ;
    wire mcs1_mcs_mat1_7_n106 ;
    wire mcs1_mcs_mat1_7_n105 ;
    wire mcs1_mcs_mat1_7_n104 ;
    wire mcs1_mcs_mat1_7_n103 ;
    wire mcs1_mcs_mat1_7_n102 ;
    wire mcs1_mcs_mat1_7_n101 ;
    wire mcs1_mcs_mat1_7_n100 ;
    wire mcs1_mcs_mat1_7_n99 ;
    wire mcs1_mcs_mat1_7_n98 ;
    wire mcs1_mcs_mat1_7_n97 ;
    wire mcs1_mcs_mat1_7_n96 ;
    wire mcs1_mcs_mat1_7_n95 ;
    wire mcs1_mcs_mat1_7_n94 ;
    wire mcs1_mcs_mat1_7_n93 ;
    wire mcs1_mcs_mat1_7_n92 ;
    wire mcs1_mcs_mat1_7_n91 ;
    wire mcs1_mcs_mat1_7_n90 ;
    wire mcs1_mcs_mat1_7_n89 ;
    wire mcs1_mcs_mat1_7_n88 ;
    wire mcs1_mcs_mat1_7_n87 ;
    wire mcs1_mcs_mat1_7_n86 ;
    wire mcs1_mcs_mat1_7_n85 ;
    wire mcs1_mcs_mat1_7_n84 ;
    wire mcs1_mcs_mat1_7_n83 ;
    wire mcs1_mcs_mat1_7_n82 ;
    wire mcs1_mcs_mat1_7_n81 ;
    wire mcs1_mcs_mat1_7_n80 ;
    wire mcs1_mcs_mat1_7_n79 ;
    wire mcs1_mcs_mat1_7_n78 ;
    wire mcs1_mcs_mat1_7_n77 ;
    wire mcs1_mcs_mat1_7_n76 ;
    wire mcs1_mcs_mat1_7_n75 ;
    wire mcs1_mcs_mat1_7_n74 ;
    wire mcs1_mcs_mat1_7_n73 ;
    wire mcs1_mcs_mat1_7_n72 ;
    wire mcs1_mcs_mat1_7_n71 ;
    wire mcs1_mcs_mat1_7_n70 ;
    wire mcs1_mcs_mat1_7_n69 ;
    wire mcs1_mcs_mat1_7_n68 ;
    wire mcs1_mcs_mat1_7_n67 ;
    wire mcs1_mcs_mat1_7_n66 ;
    wire mcs1_mcs_mat1_7_n65 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_1_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_2_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_3_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_4_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_5_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_6_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_7_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_8_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_11_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_n3 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_12_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_13_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_14_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_15_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_16_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_17_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_18_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_20_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_21_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_22_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_n4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_23_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n15 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_24_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_25_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_26_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_27_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n15 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n14 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n13 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_28_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_29_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_n6 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_n5 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_30_x0x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n12 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n11 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n10 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n9 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n8 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_n7 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x3x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x2x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x1x4 ;
    wire mcs1_mcs_mat1_7_mcs_rom0_31_x0x4 ;
    wire [127:0] addc_in ;
    wire [127:0] subc_out ;
    wire [124:1] shiftr_out ;
    wire [255:128] mcs_out ;
    wire [127:0] y0_1 ;
    wire [3:0] add_sub1_0_addc_out ;
    wire [2:0] add_sub1_0_addc_rom_ic_out ;
    wire [3:0] add_sub1_0_addc_rom_rc_out ;
    wire [3:0] add_sub1_1_addc_out ;
    wire [2:0] add_sub1_1_addc_rom_ic_out ;
    wire [3:0] add_sub1_1_addc_rom_rc_out ;
    wire [3:0] add_sub1_2_addc_out ;
    wire [2:0] add_sub1_2_addc_rom_ic_out ;
    wire [3:0] add_sub1_2_addc_rom_rc_out ;
    wire [3:0] add_sub1_3_addc_out ;
    wire [3:0] add_sub1_3_addc_rom_rc_out ;
    wire [127:0] mcs1_mcs_mat1_0_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_1_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_2_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_3_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_4_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_5_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_6_mcs_out ;
    wire [127:0] mcs1_mcs_mat1_7_mcs_out ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10778 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10793 ;
    wire new_AGEMA_signal_10794 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10797 ;
    wire new_AGEMA_signal_10798 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10801 ;
    wire new_AGEMA_signal_10802 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10805 ;
    wire new_AGEMA_signal_10806 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10809 ;
    wire new_AGEMA_signal_10810 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10813 ;
    wire new_AGEMA_signal_10814 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10817 ;
    wire new_AGEMA_signal_10818 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10821 ;
    wire new_AGEMA_signal_10822 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10825 ;
    wire new_AGEMA_signal_10826 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10829 ;
    wire new_AGEMA_signal_10830 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10833 ;
    wire new_AGEMA_signal_10834 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10837 ;
    wire new_AGEMA_signal_10838 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10841 ;
    wire new_AGEMA_signal_10842 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10845 ;
    wire new_AGEMA_signal_10846 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10849 ;
    wire new_AGEMA_signal_10850 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10853 ;
    wire new_AGEMA_signal_10854 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10857 ;
    wire new_AGEMA_signal_10858 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10861 ;
    wire new_AGEMA_signal_10862 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10865 ;
    wire new_AGEMA_signal_10866 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10874 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11197 ;
    wire new_AGEMA_signal_11198 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11201 ;
    wire new_AGEMA_signal_11202 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11205 ;
    wire new_AGEMA_signal_11206 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11209 ;
    wire new_AGEMA_signal_11210 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11213 ;
    wire new_AGEMA_signal_11214 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11217 ;
    wire new_AGEMA_signal_11218 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11221 ;
    wire new_AGEMA_signal_11222 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11225 ;
    wire new_AGEMA_signal_11226 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11229 ;
    wire new_AGEMA_signal_11230 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11233 ;
    wire new_AGEMA_signal_11234 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11237 ;
    wire new_AGEMA_signal_11238 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11241 ;
    wire new_AGEMA_signal_11242 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11245 ;
    wire new_AGEMA_signal_11246 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11249 ;
    wire new_AGEMA_signal_11250 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11253 ;
    wire new_AGEMA_signal_11254 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11257 ;
    wire new_AGEMA_signal_11258 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11261 ;
    wire new_AGEMA_signal_11262 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11265 ;
    wire new_AGEMA_signal_11266 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11269 ;
    wire new_AGEMA_signal_11270 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11273 ;
    wire new_AGEMA_signal_11274 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11277 ;
    wire new_AGEMA_signal_11278 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11281 ;
    wire new_AGEMA_signal_11282 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11285 ;
    wire new_AGEMA_signal_11286 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11289 ;
    wire new_AGEMA_signal_11290 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11293 ;
    wire new_AGEMA_signal_11294 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11297 ;
    wire new_AGEMA_signal_11298 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11301 ;
    wire new_AGEMA_signal_11302 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11305 ;
    wire new_AGEMA_signal_11306 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11309 ;
    wire new_AGEMA_signal_11310 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11313 ;
    wire new_AGEMA_signal_11314 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11317 ;
    wire new_AGEMA_signal_11318 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11321 ;
    wire new_AGEMA_signal_11322 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11645 ;
    wire new_AGEMA_signal_11646 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11649 ;
    wire new_AGEMA_signal_11650 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11653 ;
    wire new_AGEMA_signal_11654 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11657 ;
    wire new_AGEMA_signal_11658 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11661 ;
    wire new_AGEMA_signal_11662 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11665 ;
    wire new_AGEMA_signal_11666 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11669 ;
    wire new_AGEMA_signal_11670 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11673 ;
    wire new_AGEMA_signal_11674 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11677 ;
    wire new_AGEMA_signal_11678 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11681 ;
    wire new_AGEMA_signal_11682 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11685 ;
    wire new_AGEMA_signal_11686 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11689 ;
    wire new_AGEMA_signal_11690 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11693 ;
    wire new_AGEMA_signal_11694 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11697 ;
    wire new_AGEMA_signal_11698 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11701 ;
    wire new_AGEMA_signal_11702 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11705 ;
    wire new_AGEMA_signal_11706 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11709 ;
    wire new_AGEMA_signal_11710 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11713 ;
    wire new_AGEMA_signal_11714 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11717 ;
    wire new_AGEMA_signal_11718 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11721 ;
    wire new_AGEMA_signal_11722 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11725 ;
    wire new_AGEMA_signal_11726 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11729 ;
    wire new_AGEMA_signal_11730 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11733 ;
    wire new_AGEMA_signal_11734 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11737 ;
    wire new_AGEMA_signal_11738 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11741 ;
    wire new_AGEMA_signal_11742 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11745 ;
    wire new_AGEMA_signal_11746 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11749 ;
    wire new_AGEMA_signal_11750 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11753 ;
    wire new_AGEMA_signal_11754 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11757 ;
    wire new_AGEMA_signal_11758 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11761 ;
    wire new_AGEMA_signal_11762 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11765 ;
    wire new_AGEMA_signal_11766 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11769 ;
    wire new_AGEMA_signal_11770 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12087 ;
    wire new_AGEMA_signal_12088 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12091 ;
    wire new_AGEMA_signal_12092 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12095 ;
    wire new_AGEMA_signal_12096 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12099 ;
    wire new_AGEMA_signal_12100 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12103 ;
    wire new_AGEMA_signal_12104 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12107 ;
    wire new_AGEMA_signal_12108 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12111 ;
    wire new_AGEMA_signal_12112 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12115 ;
    wire new_AGEMA_signal_12116 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12119 ;
    wire new_AGEMA_signal_12120 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12123 ;
    wire new_AGEMA_signal_12124 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12127 ;
    wire new_AGEMA_signal_12128 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12131 ;
    wire new_AGEMA_signal_12132 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12135 ;
    wire new_AGEMA_signal_12136 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12139 ;
    wire new_AGEMA_signal_12140 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12143 ;
    wire new_AGEMA_signal_12144 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12147 ;
    wire new_AGEMA_signal_12148 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12151 ;
    wire new_AGEMA_signal_12152 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12155 ;
    wire new_AGEMA_signal_12156 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12159 ;
    wire new_AGEMA_signal_12160 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12163 ;
    wire new_AGEMA_signal_12164 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12167 ;
    wire new_AGEMA_signal_12168 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12171 ;
    wire new_AGEMA_signal_12172 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12175 ;
    wire new_AGEMA_signal_12176 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12179 ;
    wire new_AGEMA_signal_12180 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12183 ;
    wire new_AGEMA_signal_12184 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12187 ;
    wire new_AGEMA_signal_12188 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12191 ;
    wire new_AGEMA_signal_12192 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12195 ;
    wire new_AGEMA_signal_12196 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12199 ;
    wire new_AGEMA_signal_12200 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12313 ;
    wire new_AGEMA_signal_12314 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12317 ;
    wire new_AGEMA_signal_12318 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12321 ;
    wire new_AGEMA_signal_12322 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12325 ;
    wire new_AGEMA_signal_12326 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12329 ;
    wire new_AGEMA_signal_12330 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12333 ;
    wire new_AGEMA_signal_12334 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12337 ;
    wire new_AGEMA_signal_12338 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12341 ;
    wire new_AGEMA_signal_12342 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12345 ;
    wire new_AGEMA_signal_12346 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12349 ;
    wire new_AGEMA_signal_12350 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12353 ;
    wire new_AGEMA_signal_12354 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12357 ;
    wire new_AGEMA_signal_12358 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12361 ;
    wire new_AGEMA_signal_12362 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12365 ;
    wire new_AGEMA_signal_12366 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12369 ;
    wire new_AGEMA_signal_12370 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12373 ;
    wire new_AGEMA_signal_12374 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12377 ;
    wire new_AGEMA_signal_12378 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12381 ;
    wire new_AGEMA_signal_12382 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12385 ;
    wire new_AGEMA_signal_12386 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12389 ;
    wire new_AGEMA_signal_12390 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12393 ;
    wire new_AGEMA_signal_12394 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12397 ;
    wire new_AGEMA_signal_12398 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12401 ;
    wire new_AGEMA_signal_12402 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12405 ;
    wire new_AGEMA_signal_12406 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12409 ;
    wire new_AGEMA_signal_12410 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12413 ;
    wire new_AGEMA_signal_12414 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12417 ;
    wire new_AGEMA_signal_12418 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12421 ;
    wire new_AGEMA_signal_12422 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12425 ;
    wire new_AGEMA_signal_12426 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12429 ;
    wire new_AGEMA_signal_12430 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12433 ;
    wire new_AGEMA_signal_12434 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12437 ;
    wire new_AGEMA_signal_12438 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12441 ;
    wire new_AGEMA_signal_12442 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12445 ;
    wire new_AGEMA_signal_12446 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12449 ;
    wire new_AGEMA_signal_12450 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12453 ;
    wire new_AGEMA_signal_12454 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12457 ;
    wire new_AGEMA_signal_12458 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12461 ;
    wire new_AGEMA_signal_12462 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12465 ;
    wire new_AGEMA_signal_12466 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12469 ;
    wire new_AGEMA_signal_12470 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12473 ;
    wire new_AGEMA_signal_12474 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12477 ;
    wire new_AGEMA_signal_12478 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12481 ;
    wire new_AGEMA_signal_12482 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12485 ;
    wire new_AGEMA_signal_12486 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12489 ;
    wire new_AGEMA_signal_12490 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12493 ;
    wire new_AGEMA_signal_12494 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12497 ;
    wire new_AGEMA_signal_12498 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12501 ;
    wire new_AGEMA_signal_12502 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12505 ;
    wire new_AGEMA_signal_12506 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12509 ;
    wire new_AGEMA_signal_12510 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12513 ;
    wire new_AGEMA_signal_12514 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12517 ;
    wire new_AGEMA_signal_12518 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12521 ;
    wire new_AGEMA_signal_12522 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12525 ;
    wire new_AGEMA_signal_12526 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12529 ;
    wire new_AGEMA_signal_12530 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12533 ;
    wire new_AGEMA_signal_12534 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12537 ;
    wire new_AGEMA_signal_12538 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12541 ;
    wire new_AGEMA_signal_12542 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12545 ;
    wire new_AGEMA_signal_12546 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12549 ;
    wire new_AGEMA_signal_12550 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12553 ;
    wire new_AGEMA_signal_12554 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12557 ;
    wire new_AGEMA_signal_12558 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12561 ;
    wire new_AGEMA_signal_12562 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12565 ;
    wire new_AGEMA_signal_12566 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12569 ;
    wire new_AGEMA_signal_12570 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12573 ;
    wire new_AGEMA_signal_12574 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12577 ;
    wire new_AGEMA_signal_12578 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12581 ;
    wire new_AGEMA_signal_12582 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12585 ;
    wire new_AGEMA_signal_12586 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12589 ;
    wire new_AGEMA_signal_12590 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12593 ;
    wire new_AGEMA_signal_12594 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12597 ;
    wire new_AGEMA_signal_12598 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12601 ;
    wire new_AGEMA_signal_12602 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12605 ;
    wire new_AGEMA_signal_12606 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12609 ;
    wire new_AGEMA_signal_12610 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12613 ;
    wire new_AGEMA_signal_12614 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12617 ;
    wire new_AGEMA_signal_12618 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12621 ;
    wire new_AGEMA_signal_12622 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12625 ;
    wire new_AGEMA_signal_12626 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12629 ;
    wire new_AGEMA_signal_12630 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12633 ;
    wire new_AGEMA_signal_12634 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12637 ;
    wire new_AGEMA_signal_12638 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12641 ;
    wire new_AGEMA_signal_12642 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12645 ;
    wire new_AGEMA_signal_12646 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12649 ;
    wire new_AGEMA_signal_12650 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12653 ;
    wire new_AGEMA_signal_12654 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12657 ;
    wire new_AGEMA_signal_12658 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12661 ;
    wire new_AGEMA_signal_12662 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12665 ;
    wire new_AGEMA_signal_12666 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12669 ;
    wire new_AGEMA_signal_12670 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12673 ;
    wire new_AGEMA_signal_12674 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12677 ;
    wire new_AGEMA_signal_12678 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12681 ;
    wire new_AGEMA_signal_12682 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12685 ;
    wire new_AGEMA_signal_12686 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12689 ;
    wire new_AGEMA_signal_12690 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12693 ;
    wire new_AGEMA_signal_12694 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12697 ;
    wire new_AGEMA_signal_12698 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12701 ;
    wire new_AGEMA_signal_12702 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12705 ;
    wire new_AGEMA_signal_12706 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12709 ;
    wire new_AGEMA_signal_12710 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12713 ;
    wire new_AGEMA_signal_12714 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12717 ;
    wire new_AGEMA_signal_12718 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12721 ;
    wire new_AGEMA_signal_12722 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12725 ;
    wire new_AGEMA_signal_12726 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12729 ;
    wire new_AGEMA_signal_12730 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12733 ;
    wire new_AGEMA_signal_12734 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12737 ;
    wire new_AGEMA_signal_12738 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12741 ;
    wire new_AGEMA_signal_12742 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12745 ;
    wire new_AGEMA_signal_12746 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12749 ;
    wire new_AGEMA_signal_12750 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12753 ;
    wire new_AGEMA_signal_12754 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12757 ;
    wire new_AGEMA_signal_12758 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12761 ;
    wire new_AGEMA_signal_12762 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12765 ;
    wire new_AGEMA_signal_12766 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12769 ;
    wire new_AGEMA_signal_12770 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12773 ;
    wire new_AGEMA_signal_12774 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12777 ;
    wire new_AGEMA_signal_12778 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12781 ;
    wire new_AGEMA_signal_12782 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12785 ;
    wire new_AGEMA_signal_12786 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12789 ;
    wire new_AGEMA_signal_12790 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12793 ;
    wire new_AGEMA_signal_12794 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12797 ;
    wire new_AGEMA_signal_12798 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12801 ;
    wire new_AGEMA_signal_12802 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12805 ;
    wire new_AGEMA_signal_12806 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12809 ;
    wire new_AGEMA_signal_12810 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12813 ;
    wire new_AGEMA_signal_12814 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12817 ;
    wire new_AGEMA_signal_12818 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12821 ;
    wire new_AGEMA_signal_12822 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12825 ;
    wire new_AGEMA_signal_12826 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12829 ;
    wire new_AGEMA_signal_12830 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12833 ;
    wire new_AGEMA_signal_12834 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12837 ;
    wire new_AGEMA_signal_12838 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12841 ;
    wire new_AGEMA_signal_12842 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12845 ;
    wire new_AGEMA_signal_12846 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12849 ;
    wire new_AGEMA_signal_12850 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_12853 ;
    wire new_AGEMA_signal_12854 ;
    wire new_AGEMA_signal_12855 ;
    wire new_AGEMA_signal_12856 ;
    wire new_AGEMA_signal_12857 ;
    wire new_AGEMA_signal_12858 ;
    wire new_AGEMA_signal_12859 ;
    wire new_AGEMA_signal_12860 ;
    wire new_AGEMA_signal_12861 ;
    wire new_AGEMA_signal_12862 ;
    wire new_AGEMA_signal_12863 ;
    wire new_AGEMA_signal_12864 ;
    wire new_AGEMA_signal_12865 ;
    wire new_AGEMA_signal_12866 ;
    wire new_AGEMA_signal_12867 ;
    wire new_AGEMA_signal_12868 ;
    wire new_AGEMA_signal_12869 ;
    wire new_AGEMA_signal_12870 ;
    wire new_AGEMA_signal_12871 ;
    wire new_AGEMA_signal_12872 ;
    wire new_AGEMA_signal_12873 ;
    wire new_AGEMA_signal_12874 ;
    wire new_AGEMA_signal_12875 ;
    wire new_AGEMA_signal_12876 ;
    wire new_AGEMA_signal_12877 ;
    wire new_AGEMA_signal_12878 ;
    wire new_AGEMA_signal_12879 ;
    wire new_AGEMA_signal_12880 ;
    wire new_AGEMA_signal_12881 ;
    wire new_AGEMA_signal_12882 ;
    wire new_AGEMA_signal_12883 ;
    wire new_AGEMA_signal_12884 ;
    wire new_AGEMA_signal_12885 ;
    wire new_AGEMA_signal_12886 ;
    wire new_AGEMA_signal_12887 ;
    wire new_AGEMA_signal_12888 ;
    wire new_AGEMA_signal_12889 ;
    wire new_AGEMA_signal_12890 ;
    wire new_AGEMA_signal_12891 ;
    wire new_AGEMA_signal_12892 ;
    wire new_AGEMA_signal_12893 ;
    wire new_AGEMA_signal_12894 ;
    wire new_AGEMA_signal_12895 ;
    wire new_AGEMA_signal_12896 ;
    wire new_AGEMA_signal_12897 ;
    wire new_AGEMA_signal_12898 ;
    wire new_AGEMA_signal_12899 ;
    wire new_AGEMA_signal_12900 ;
    wire new_AGEMA_signal_12901 ;
    wire new_AGEMA_signal_12902 ;
    wire new_AGEMA_signal_12903 ;
    wire new_AGEMA_signal_12904 ;
    wire new_AGEMA_signal_12905 ;
    wire new_AGEMA_signal_12906 ;
    wire new_AGEMA_signal_12907 ;
    wire new_AGEMA_signal_12908 ;
    wire new_AGEMA_signal_12909 ;
    wire new_AGEMA_signal_12910 ;
    wire new_AGEMA_signal_12911 ;
    wire new_AGEMA_signal_12912 ;
    wire new_AGEMA_signal_12913 ;
    wire new_AGEMA_signal_12914 ;
    wire new_AGEMA_signal_12915 ;
    wire new_AGEMA_signal_12916 ;
    wire new_AGEMA_signal_12917 ;
    wire new_AGEMA_signal_12918 ;
    wire new_AGEMA_signal_12919 ;
    wire new_AGEMA_signal_12920 ;
    wire new_AGEMA_signal_12921 ;
    wire new_AGEMA_signal_12922 ;
    wire new_AGEMA_signal_12923 ;
    wire new_AGEMA_signal_12924 ;
    wire new_AGEMA_signal_12925 ;
    wire new_AGEMA_signal_12926 ;
    wire new_AGEMA_signal_12927 ;
    wire new_AGEMA_signal_12928 ;
    wire new_AGEMA_signal_12929 ;
    wire new_AGEMA_signal_12930 ;
    wire new_AGEMA_signal_12931 ;
    wire new_AGEMA_signal_12932 ;
    wire new_AGEMA_signal_12933 ;
    wire new_AGEMA_signal_12934 ;
    wire new_AGEMA_signal_12935 ;
    wire new_AGEMA_signal_12936 ;
    wire new_AGEMA_signal_12937 ;
    wire new_AGEMA_signal_12938 ;
    wire new_AGEMA_signal_12939 ;
    wire new_AGEMA_signal_12940 ;
    wire new_AGEMA_signal_12941 ;
    wire new_AGEMA_signal_12942 ;
    wire new_AGEMA_signal_12943 ;
    wire new_AGEMA_signal_12944 ;
    wire new_AGEMA_signal_12945 ;
    wire new_AGEMA_signal_12946 ;
    wire new_AGEMA_signal_12947 ;
    wire new_AGEMA_signal_12948 ;
    wire new_AGEMA_signal_12949 ;
    wire new_AGEMA_signal_12950 ;
    wire new_AGEMA_signal_12951 ;
    wire new_AGEMA_signal_12952 ;
    wire new_AGEMA_signal_12953 ;
    wire new_AGEMA_signal_12954 ;
    wire new_AGEMA_signal_12955 ;
    wire new_AGEMA_signal_12956 ;
    wire new_AGEMA_signal_12957 ;
    wire new_AGEMA_signal_12958 ;
    wire new_AGEMA_signal_12959 ;
    wire new_AGEMA_signal_12960 ;
    wire new_AGEMA_signal_12961 ;
    wire new_AGEMA_signal_12962 ;
    wire new_AGEMA_signal_12963 ;
    wire new_AGEMA_signal_12964 ;
    wire new_AGEMA_signal_12965 ;
    wire new_AGEMA_signal_12966 ;
    wire new_AGEMA_signal_12967 ;
    wire new_AGEMA_signal_12968 ;
    wire new_AGEMA_signal_12969 ;
    wire new_AGEMA_signal_12970 ;
    wire new_AGEMA_signal_12971 ;
    wire new_AGEMA_signal_12972 ;
    wire new_AGEMA_signal_12973 ;
    wire new_AGEMA_signal_12974 ;
    wire new_AGEMA_signal_12975 ;
    wire new_AGEMA_signal_12976 ;
    wire new_AGEMA_signal_12977 ;
    wire new_AGEMA_signal_12978 ;
    wire new_AGEMA_signal_12979 ;
    wire new_AGEMA_signal_12980 ;
    wire new_AGEMA_signal_12981 ;
    wire new_AGEMA_signal_12982 ;
    wire new_AGEMA_signal_12983 ;
    wire new_AGEMA_signal_12984 ;
    wire new_AGEMA_signal_12985 ;
    wire new_AGEMA_signal_12986 ;
    wire new_AGEMA_signal_12987 ;
    wire new_AGEMA_signal_12988 ;
    wire new_AGEMA_signal_12989 ;
    wire new_AGEMA_signal_12990 ;
    wire new_AGEMA_signal_12991 ;
    wire new_AGEMA_signal_12992 ;
    wire new_AGEMA_signal_12993 ;
    wire new_AGEMA_signal_12994 ;
    wire new_AGEMA_signal_12995 ;
    wire new_AGEMA_signal_12996 ;
    wire new_AGEMA_signal_12997 ;
    wire new_AGEMA_signal_12998 ;
    wire new_AGEMA_signal_12999 ;
    wire new_AGEMA_signal_13000 ;
    wire new_AGEMA_signal_13001 ;
    wire new_AGEMA_signal_13002 ;
    wire new_AGEMA_signal_13003 ;
    wire new_AGEMA_signal_13004 ;
    wire new_AGEMA_signal_13005 ;
    wire new_AGEMA_signal_13006 ;
    wire new_AGEMA_signal_13007 ;
    wire new_AGEMA_signal_13008 ;
    wire new_AGEMA_signal_13009 ;
    wire new_AGEMA_signal_13010 ;
    wire new_AGEMA_signal_13011 ;
    wire new_AGEMA_signal_13012 ;
    wire new_AGEMA_signal_13013 ;
    wire new_AGEMA_signal_13014 ;
    wire new_AGEMA_signal_13015 ;
    wire new_AGEMA_signal_13016 ;
    wire new_AGEMA_signal_13017 ;
    wire new_AGEMA_signal_13018 ;
    wire new_AGEMA_signal_13019 ;
    wire new_AGEMA_signal_13020 ;
    wire new_AGEMA_signal_13021 ;
    wire new_AGEMA_signal_13022 ;
    wire new_AGEMA_signal_13023 ;
    wire new_AGEMA_signal_13024 ;
    wire new_AGEMA_signal_13025 ;
    wire new_AGEMA_signal_13026 ;
    wire new_AGEMA_signal_13027 ;
    wire new_AGEMA_signal_13028 ;
    wire new_AGEMA_signal_13029 ;
    wire new_AGEMA_signal_13030 ;
    wire new_AGEMA_signal_13031 ;
    wire new_AGEMA_signal_13032 ;
    wire new_AGEMA_signal_13033 ;
    wire new_AGEMA_signal_13034 ;
    wire new_AGEMA_signal_13035 ;
    wire new_AGEMA_signal_13036 ;
    wire new_AGEMA_signal_13037 ;
    wire new_AGEMA_signal_13038 ;
    wire new_AGEMA_signal_13039 ;
    wire new_AGEMA_signal_13040 ;
    wire new_AGEMA_signal_13041 ;
    wire new_AGEMA_signal_13042 ;
    wire new_AGEMA_signal_13043 ;
    wire new_AGEMA_signal_13044 ;
    wire new_AGEMA_signal_13045 ;
    wire new_AGEMA_signal_13046 ;
    wire new_AGEMA_signal_13047 ;
    wire new_AGEMA_signal_13048 ;
    wire new_AGEMA_signal_13049 ;
    wire new_AGEMA_signal_13050 ;
    wire new_AGEMA_signal_13051 ;
    wire new_AGEMA_signal_13052 ;
    wire new_AGEMA_signal_13053 ;
    wire new_AGEMA_signal_13054 ;
    wire new_AGEMA_signal_13055 ;
    wire new_AGEMA_signal_13056 ;
    wire new_AGEMA_signal_13057 ;
    wire new_AGEMA_signal_13058 ;
    wire new_AGEMA_signal_13059 ;
    wire new_AGEMA_signal_13060 ;
    wire new_AGEMA_signal_13061 ;
    wire new_AGEMA_signal_13062 ;
    wire new_AGEMA_signal_13063 ;
    wire new_AGEMA_signal_13064 ;
    wire new_AGEMA_signal_13065 ;
    wire new_AGEMA_signal_13066 ;
    wire new_AGEMA_signal_13067 ;
    wire new_AGEMA_signal_13068 ;
    wire new_AGEMA_signal_13069 ;
    wire new_AGEMA_signal_13070 ;
    wire new_AGEMA_signal_13071 ;
    wire new_AGEMA_signal_13072 ;
    wire new_AGEMA_signal_13073 ;
    wire new_AGEMA_signal_13074 ;
    wire new_AGEMA_signal_13075 ;
    wire new_AGEMA_signal_13076 ;
    wire new_AGEMA_signal_13077 ;
    wire new_AGEMA_signal_13078 ;
    wire new_AGEMA_signal_13079 ;
    wire new_AGEMA_signal_13080 ;
    wire new_AGEMA_signal_13081 ;
    wire new_AGEMA_signal_13082 ;
    wire new_AGEMA_signal_13083 ;
    wire new_AGEMA_signal_13084 ;
    wire new_AGEMA_signal_13085 ;
    wire new_AGEMA_signal_13086 ;
    wire new_AGEMA_signal_13087 ;
    wire new_AGEMA_signal_13088 ;
    wire new_AGEMA_signal_13089 ;
    wire new_AGEMA_signal_13090 ;
    wire new_AGEMA_signal_13091 ;
    wire new_AGEMA_signal_13092 ;
    wire new_AGEMA_signal_13093 ;
    wire new_AGEMA_signal_13094 ;
    wire new_AGEMA_signal_13095 ;
    wire new_AGEMA_signal_13096 ;
    wire new_AGEMA_signal_13097 ;
    wire new_AGEMA_signal_13098 ;
    wire new_AGEMA_signal_13099 ;
    wire new_AGEMA_signal_13100 ;
    wire new_AGEMA_signal_13101 ;
    wire new_AGEMA_signal_13102 ;
    wire new_AGEMA_signal_13103 ;
    wire new_AGEMA_signal_13104 ;
    wire new_AGEMA_signal_13105 ;
    wire new_AGEMA_signal_13106 ;
    wire new_AGEMA_signal_13107 ;
    wire new_AGEMA_signal_13108 ;
    wire new_AGEMA_signal_13109 ;
    wire new_AGEMA_signal_13110 ;
    wire new_AGEMA_signal_13111 ;
    wire new_AGEMA_signal_13112 ;
    wire new_AGEMA_signal_13113 ;
    wire new_AGEMA_signal_13114 ;
    wire new_AGEMA_signal_13115 ;
    wire new_AGEMA_signal_13116 ;
    wire new_AGEMA_signal_13117 ;
    wire new_AGEMA_signal_13118 ;
    wire new_AGEMA_signal_13119 ;
    wire new_AGEMA_signal_13120 ;
    wire new_AGEMA_signal_13121 ;
    wire new_AGEMA_signal_13122 ;
    wire new_AGEMA_signal_13123 ;
    wire new_AGEMA_signal_13124 ;
    wire new_AGEMA_signal_13125 ;
    wire new_AGEMA_signal_13126 ;
    wire new_AGEMA_signal_13127 ;
    wire new_AGEMA_signal_13128 ;
    wire new_AGEMA_signal_13129 ;
    wire new_AGEMA_signal_13130 ;
    wire new_AGEMA_signal_13131 ;
    wire new_AGEMA_signal_13132 ;
    wire new_AGEMA_signal_13133 ;
    wire new_AGEMA_signal_13134 ;
    wire new_AGEMA_signal_13135 ;
    wire new_AGEMA_signal_13136 ;
    wire new_AGEMA_signal_13137 ;
    wire new_AGEMA_signal_13138 ;
    wire new_AGEMA_signal_13139 ;
    wire new_AGEMA_signal_13140 ;
    wire new_AGEMA_signal_13141 ;
    wire new_AGEMA_signal_13142 ;
    wire new_AGEMA_signal_13143 ;
    wire new_AGEMA_signal_13144 ;
    wire new_AGEMA_signal_13145 ;
    wire new_AGEMA_signal_13146 ;
    wire new_AGEMA_signal_13147 ;
    wire new_AGEMA_signal_13148 ;
    wire new_AGEMA_signal_13149 ;
    wire new_AGEMA_signal_13150 ;
    wire new_AGEMA_signal_13151 ;
    wire new_AGEMA_signal_13152 ;
    wire new_AGEMA_signal_13153 ;
    wire new_AGEMA_signal_13154 ;
    wire new_AGEMA_signal_13155 ;
    wire new_AGEMA_signal_13156 ;
    wire new_AGEMA_signal_13157 ;
    wire new_AGEMA_signal_13158 ;
    wire new_AGEMA_signal_13159 ;
    wire new_AGEMA_signal_13160 ;
    wire new_AGEMA_signal_13161 ;
    wire new_AGEMA_signal_13162 ;
    wire new_AGEMA_signal_13163 ;
    wire new_AGEMA_signal_13164 ;
    wire new_AGEMA_signal_13165 ;
    wire new_AGEMA_signal_13166 ;
    wire new_AGEMA_signal_13167 ;
    wire new_AGEMA_signal_13168 ;
    wire new_AGEMA_signal_13169 ;
    wire new_AGEMA_signal_13170 ;
    wire new_AGEMA_signal_13171 ;
    wire new_AGEMA_signal_13172 ;
    wire new_AGEMA_signal_13173 ;
    wire new_AGEMA_signal_13174 ;
    wire new_AGEMA_signal_13175 ;
    wire new_AGEMA_signal_13176 ;
    wire new_AGEMA_signal_13177 ;
    wire new_AGEMA_signal_13178 ;
    wire new_AGEMA_signal_13179 ;
    wire new_AGEMA_signal_13180 ;
    wire new_AGEMA_signal_13181 ;
    wire new_AGEMA_signal_13182 ;
    wire new_AGEMA_signal_13183 ;
    wire new_AGEMA_signal_13184 ;
    wire new_AGEMA_signal_13185 ;
    wire new_AGEMA_signal_13186 ;
    wire new_AGEMA_signal_13187 ;
    wire new_AGEMA_signal_13188 ;
    wire new_AGEMA_signal_13189 ;
    wire new_AGEMA_signal_13190 ;
    wire new_AGEMA_signal_13191 ;
    wire new_AGEMA_signal_13192 ;
    wire new_AGEMA_signal_13193 ;
    wire new_AGEMA_signal_13194 ;
    wire new_AGEMA_signal_13195 ;
    wire new_AGEMA_signal_13196 ;
    wire new_AGEMA_signal_13197 ;
    wire new_AGEMA_signal_13198 ;
    wire new_AGEMA_signal_13199 ;
    wire new_AGEMA_signal_13200 ;
    wire new_AGEMA_signal_13201 ;
    wire new_AGEMA_signal_13202 ;
    wire new_AGEMA_signal_13203 ;
    wire new_AGEMA_signal_13204 ;
    wire new_AGEMA_signal_13205 ;
    wire new_AGEMA_signal_13206 ;
    wire new_AGEMA_signal_13207 ;
    wire new_AGEMA_signal_13208 ;
    wire new_AGEMA_signal_13209 ;
    wire new_AGEMA_signal_13210 ;
    wire new_AGEMA_signal_13211 ;
    wire new_AGEMA_signal_13212 ;
    wire new_AGEMA_signal_13213 ;
    wire new_AGEMA_signal_13214 ;
    wire new_AGEMA_signal_13215 ;
    wire new_AGEMA_signal_13216 ;
    wire new_AGEMA_signal_13217 ;
    wire new_AGEMA_signal_13218 ;
    wire new_AGEMA_signal_13219 ;
    wire new_AGEMA_signal_13220 ;
    wire new_AGEMA_signal_13221 ;
    wire new_AGEMA_signal_13222 ;
    wire new_AGEMA_signal_13223 ;
    wire new_AGEMA_signal_13224 ;
    wire new_AGEMA_signal_13225 ;
    wire new_AGEMA_signal_13226 ;
    wire new_AGEMA_signal_13227 ;
    wire new_AGEMA_signal_13228 ;
    wire new_AGEMA_signal_13229 ;
    wire new_AGEMA_signal_13230 ;
    wire new_AGEMA_signal_13231 ;
    wire new_AGEMA_signal_13232 ;
    wire new_AGEMA_signal_13233 ;
    wire new_AGEMA_signal_13234 ;
    wire new_AGEMA_signal_13235 ;
    wire new_AGEMA_signal_13236 ;
    wire new_AGEMA_signal_13237 ;
    wire new_AGEMA_signal_13238 ;
    wire new_AGEMA_signal_13239 ;
    wire new_AGEMA_signal_13240 ;
    wire new_AGEMA_signal_13241 ;
    wire new_AGEMA_signal_13242 ;
    wire new_AGEMA_signal_13243 ;
    wire new_AGEMA_signal_13244 ;
    wire new_AGEMA_signal_13245 ;
    wire new_AGEMA_signal_13246 ;
    wire new_AGEMA_signal_13247 ;
    wire new_AGEMA_signal_13248 ;
    wire new_AGEMA_signal_13249 ;
    wire new_AGEMA_signal_13250 ;
    wire new_AGEMA_signal_13251 ;
    wire new_AGEMA_signal_13252 ;
    wire new_AGEMA_signal_13253 ;
    wire new_AGEMA_signal_13254 ;
    wire new_AGEMA_signal_13255 ;
    wire new_AGEMA_signal_13256 ;
    wire new_AGEMA_signal_13257 ;
    wire new_AGEMA_signal_13258 ;
    wire new_AGEMA_signal_13259 ;
    wire new_AGEMA_signal_13260 ;
    wire new_AGEMA_signal_13261 ;
    wire new_AGEMA_signal_13262 ;
    wire new_AGEMA_signal_13263 ;
    wire new_AGEMA_signal_13264 ;
    wire new_AGEMA_signal_13265 ;
    wire new_AGEMA_signal_13266 ;
    wire new_AGEMA_signal_13267 ;
    wire new_AGEMA_signal_13268 ;
    wire new_AGEMA_signal_13269 ;
    wire new_AGEMA_signal_13270 ;
    wire new_AGEMA_signal_13271 ;
    wire new_AGEMA_signal_13272 ;
    wire new_AGEMA_signal_13273 ;
    wire new_AGEMA_signal_13274 ;
    wire new_AGEMA_signal_13275 ;
    wire new_AGEMA_signal_13276 ;
    wire new_AGEMA_signal_13277 ;
    wire new_AGEMA_signal_13278 ;
    wire new_AGEMA_signal_13279 ;
    wire new_AGEMA_signal_13280 ;
    wire new_AGEMA_signal_13281 ;
    wire new_AGEMA_signal_13282 ;
    wire new_AGEMA_signal_13283 ;
    wire new_AGEMA_signal_13284 ;
    wire new_AGEMA_signal_13285 ;
    wire new_AGEMA_signal_13286 ;
    wire new_AGEMA_signal_13287 ;
    wire new_AGEMA_signal_13288 ;
    wire new_AGEMA_signal_13289 ;
    wire new_AGEMA_signal_13290 ;
    wire new_AGEMA_signal_13291 ;
    wire new_AGEMA_signal_13292 ;
    wire new_AGEMA_signal_13293 ;
    wire new_AGEMA_signal_13294 ;
    wire new_AGEMA_signal_13295 ;
    wire new_AGEMA_signal_13296 ;
    wire new_AGEMA_signal_13297 ;
    wire new_AGEMA_signal_13298 ;
    wire new_AGEMA_signal_13299 ;
    wire new_AGEMA_signal_13300 ;
    wire new_AGEMA_signal_13301 ;
    wire new_AGEMA_signal_13302 ;
    wire new_AGEMA_signal_13303 ;
    wire new_AGEMA_signal_13304 ;
    wire new_AGEMA_signal_13305 ;
    wire new_AGEMA_signal_13306 ;
    wire new_AGEMA_signal_13307 ;
    wire new_AGEMA_signal_13308 ;
    wire new_AGEMA_signal_13309 ;
    wire new_AGEMA_signal_13310 ;
    wire new_AGEMA_signal_13311 ;
    wire new_AGEMA_signal_13312 ;
    wire new_AGEMA_signal_13313 ;
    wire new_AGEMA_signal_13314 ;
    wire new_AGEMA_signal_13315 ;
    wire new_AGEMA_signal_13316 ;
    wire new_AGEMA_signal_13317 ;
    wire new_AGEMA_signal_13318 ;
    wire new_AGEMA_signal_13319 ;
    wire new_AGEMA_signal_13320 ;
    wire new_AGEMA_signal_13321 ;
    wire new_AGEMA_signal_13322 ;
    wire new_AGEMA_signal_13323 ;
    wire new_AGEMA_signal_13324 ;
    wire new_AGEMA_signal_13325 ;
    wire new_AGEMA_signal_13326 ;
    wire new_AGEMA_signal_13327 ;
    wire new_AGEMA_signal_13328 ;
    wire new_AGEMA_signal_13329 ;
    wire new_AGEMA_signal_13330 ;
    wire new_AGEMA_signal_13331 ;
    wire new_AGEMA_signal_13332 ;
    wire new_AGEMA_signal_13333 ;
    wire new_AGEMA_signal_13334 ;
    wire new_AGEMA_signal_13335 ;
    wire new_AGEMA_signal_13336 ;
    wire new_AGEMA_signal_13337 ;
    wire new_AGEMA_signal_13338 ;
    wire new_AGEMA_signal_13339 ;
    wire new_AGEMA_signal_13340 ;
    wire new_AGEMA_signal_13341 ;
    wire new_AGEMA_signal_13342 ;
    wire new_AGEMA_signal_13343 ;
    wire new_AGEMA_signal_13344 ;
    wire new_AGEMA_signal_13345 ;
    wire new_AGEMA_signal_13346 ;
    wire new_AGEMA_signal_13347 ;
    wire new_AGEMA_signal_13348 ;
    wire new_AGEMA_signal_13349 ;
    wire new_AGEMA_signal_13350 ;
    wire new_AGEMA_signal_13351 ;
    wire new_AGEMA_signal_13352 ;
    wire new_AGEMA_signal_13353 ;
    wire new_AGEMA_signal_13354 ;
    wire new_AGEMA_signal_13355 ;
    wire new_AGEMA_signal_13356 ;
    wire new_AGEMA_signal_13357 ;
    wire new_AGEMA_signal_13358 ;
    wire new_AGEMA_signal_13359 ;
    wire new_AGEMA_signal_13360 ;
    wire new_AGEMA_signal_13361 ;
    wire new_AGEMA_signal_13362 ;
    wire new_AGEMA_signal_13363 ;
    wire new_AGEMA_signal_13364 ;
    wire new_AGEMA_signal_13365 ;
    wire new_AGEMA_signal_13366 ;
    wire new_AGEMA_signal_13367 ;
    wire new_AGEMA_signal_13368 ;
    wire new_AGEMA_signal_13369 ;
    wire new_AGEMA_signal_13370 ;
    wire new_AGEMA_signal_13371 ;
    wire new_AGEMA_signal_13372 ;
    wire new_AGEMA_signal_13373 ;
    wire new_AGEMA_signal_13374 ;
    wire new_AGEMA_signal_13375 ;
    wire new_AGEMA_signal_13376 ;
    wire new_AGEMA_signal_13377 ;
    wire new_AGEMA_signal_13378 ;
    wire new_AGEMA_signal_13379 ;
    wire new_AGEMA_signal_13380 ;
    wire new_AGEMA_signal_13381 ;
    wire new_AGEMA_signal_13382 ;
    wire new_AGEMA_signal_13383 ;
    wire new_AGEMA_signal_13384 ;
    wire new_AGEMA_signal_13385 ;
    wire new_AGEMA_signal_13386 ;
    wire new_AGEMA_signal_13387 ;
    wire new_AGEMA_signal_13388 ;
    wire new_AGEMA_signal_13389 ;
    wire new_AGEMA_signal_13390 ;
    wire new_AGEMA_signal_13391 ;
    wire new_AGEMA_signal_13392 ;
    wire new_AGEMA_signal_13393 ;
    wire new_AGEMA_signal_13394 ;
    wire new_AGEMA_signal_13395 ;
    wire new_AGEMA_signal_13396 ;
    wire new_AGEMA_signal_13397 ;
    wire new_AGEMA_signal_13398 ;
    wire new_AGEMA_signal_13399 ;
    wire new_AGEMA_signal_13400 ;
    wire new_AGEMA_signal_13401 ;
    wire new_AGEMA_signal_13402 ;
    wire new_AGEMA_signal_13403 ;
    wire new_AGEMA_signal_13404 ;
    wire new_AGEMA_signal_13405 ;
    wire new_AGEMA_signal_13406 ;
    wire new_AGEMA_signal_13407 ;
    wire new_AGEMA_signal_13408 ;
    wire new_AGEMA_signal_13409 ;
    wire new_AGEMA_signal_13410 ;
    wire new_AGEMA_signal_13411 ;
    wire new_AGEMA_signal_13412 ;
    wire new_AGEMA_signal_13413 ;
    wire new_AGEMA_signal_13414 ;
    wire new_AGEMA_signal_13415 ;
    wire new_AGEMA_signal_13416 ;
    wire new_AGEMA_signal_13417 ;
    wire new_AGEMA_signal_13418 ;
    wire new_AGEMA_signal_13419 ;
    wire new_AGEMA_signal_13420 ;
    wire new_AGEMA_signal_13421 ;
    wire new_AGEMA_signal_13422 ;
    wire new_AGEMA_signal_13423 ;
    wire new_AGEMA_signal_13424 ;
    wire new_AGEMA_signal_13425 ;
    wire new_AGEMA_signal_13426 ;
    wire new_AGEMA_signal_13427 ;
    wire new_AGEMA_signal_13428 ;
    wire new_AGEMA_signal_13429 ;
    wire new_AGEMA_signal_13430 ;
    wire new_AGEMA_signal_13431 ;
    wire new_AGEMA_signal_13432 ;
    wire new_AGEMA_signal_13433 ;
    wire new_AGEMA_signal_13434 ;
    wire new_AGEMA_signal_13435 ;
    wire new_AGEMA_signal_13436 ;
    wire new_AGEMA_signal_13437 ;
    wire new_AGEMA_signal_13438 ;
    wire new_AGEMA_signal_13439 ;
    wire new_AGEMA_signal_13440 ;
    wire new_AGEMA_signal_13441 ;
    wire new_AGEMA_signal_13442 ;
    wire new_AGEMA_signal_13443 ;
    wire new_AGEMA_signal_13444 ;
    wire new_AGEMA_signal_13445 ;
    wire new_AGEMA_signal_13446 ;
    wire new_AGEMA_signal_13447 ;
    wire new_AGEMA_signal_13448 ;
    wire new_AGEMA_signal_13449 ;
    wire new_AGEMA_signal_13450 ;
    wire new_AGEMA_signal_13451 ;
    wire new_AGEMA_signal_13452 ;
    wire new_AGEMA_signal_13453 ;
    wire new_AGEMA_signal_13454 ;
    wire new_AGEMA_signal_13455 ;
    wire new_AGEMA_signal_13456 ;
    wire new_AGEMA_signal_13457 ;
    wire new_AGEMA_signal_13458 ;
    wire new_AGEMA_signal_13459 ;
    wire new_AGEMA_signal_13460 ;
    wire new_AGEMA_signal_13461 ;
    wire new_AGEMA_signal_13462 ;
    wire new_AGEMA_signal_13463 ;
    wire new_AGEMA_signal_13464 ;
    wire new_AGEMA_signal_13465 ;
    wire new_AGEMA_signal_13466 ;
    wire new_AGEMA_signal_13467 ;
    wire new_AGEMA_signal_13468 ;
    wire new_AGEMA_signal_13469 ;
    wire new_AGEMA_signal_13470 ;
    wire new_AGEMA_signal_13471 ;
    wire new_AGEMA_signal_13472 ;
    wire new_AGEMA_signal_13473 ;
    wire new_AGEMA_signal_13474 ;
    wire new_AGEMA_signal_13475 ;
    wire new_AGEMA_signal_13476 ;
    wire new_AGEMA_signal_13477 ;
    wire new_AGEMA_signal_13478 ;
    wire new_AGEMA_signal_13479 ;
    wire new_AGEMA_signal_13480 ;
    wire new_AGEMA_signal_13481 ;
    wire new_AGEMA_signal_13482 ;
    wire new_AGEMA_signal_13483 ;
    wire new_AGEMA_signal_13484 ;
    wire new_AGEMA_signal_13485 ;
    wire new_AGEMA_signal_13486 ;
    wire new_AGEMA_signal_13487 ;
    wire new_AGEMA_signal_13488 ;
    wire new_AGEMA_signal_13489 ;
    wire new_AGEMA_signal_13490 ;
    wire new_AGEMA_signal_13491 ;
    wire new_AGEMA_signal_13492 ;
    wire new_AGEMA_signal_13493 ;
    wire new_AGEMA_signal_13494 ;
    wire new_AGEMA_signal_13495 ;
    wire new_AGEMA_signal_13496 ;
    wire new_AGEMA_signal_13497 ;
    wire new_AGEMA_signal_13498 ;
    wire new_AGEMA_signal_13499 ;
    wire new_AGEMA_signal_13500 ;
    wire new_AGEMA_signal_13501 ;
    wire new_AGEMA_signal_13502 ;
    wire new_AGEMA_signal_13503 ;
    wire new_AGEMA_signal_13504 ;
    wire new_AGEMA_signal_13505 ;
    wire new_AGEMA_signal_13506 ;
    wire new_AGEMA_signal_13507 ;
    wire new_AGEMA_signal_13508 ;
    wire new_AGEMA_signal_13509 ;
    wire new_AGEMA_signal_13510 ;
    wire new_AGEMA_signal_13511 ;
    wire new_AGEMA_signal_13512 ;
    wire new_AGEMA_signal_13513 ;
    wire new_AGEMA_signal_13514 ;
    wire new_AGEMA_signal_13515 ;
    wire new_AGEMA_signal_13516 ;
    wire new_AGEMA_signal_13517 ;
    wire new_AGEMA_signal_13518 ;
    wire new_AGEMA_signal_13519 ;
    wire new_AGEMA_signal_13520 ;
    wire new_AGEMA_signal_13521 ;
    wire new_AGEMA_signal_13522 ;
    wire new_AGEMA_signal_13523 ;
    wire new_AGEMA_signal_13524 ;
    wire new_AGEMA_signal_13525 ;
    wire new_AGEMA_signal_13526 ;
    wire new_AGEMA_signal_13527 ;
    wire new_AGEMA_signal_13528 ;
    wire new_AGEMA_signal_13529 ;
    wire new_AGEMA_signal_13530 ;
    wire new_AGEMA_signal_13531 ;
    wire new_AGEMA_signal_13532 ;
    wire new_AGEMA_signal_13533 ;
    wire new_AGEMA_signal_13534 ;
    wire new_AGEMA_signal_13535 ;
    wire new_AGEMA_signal_13536 ;
    wire new_AGEMA_signal_13537 ;
    wire new_AGEMA_signal_13538 ;
    wire new_AGEMA_signal_13539 ;
    wire new_AGEMA_signal_13540 ;
    wire new_AGEMA_signal_13541 ;
    wire new_AGEMA_signal_13542 ;
    wire new_AGEMA_signal_13543 ;
    wire new_AGEMA_signal_13544 ;
    wire new_AGEMA_signal_13545 ;
    wire new_AGEMA_signal_13546 ;
    wire new_AGEMA_signal_13547 ;
    wire new_AGEMA_signal_13548 ;
    wire new_AGEMA_signal_13549 ;
    wire new_AGEMA_signal_13550 ;
    wire new_AGEMA_signal_13551 ;
    wire new_AGEMA_signal_13552 ;
    wire new_AGEMA_signal_13553 ;
    wire new_AGEMA_signal_13554 ;
    wire new_AGEMA_signal_13555 ;
    wire new_AGEMA_signal_13556 ;
    wire new_AGEMA_signal_13557 ;
    wire new_AGEMA_signal_13558 ;
    wire new_AGEMA_signal_13559 ;
    wire new_AGEMA_signal_13560 ;
    wire new_AGEMA_signal_13561 ;
    wire new_AGEMA_signal_13562 ;
    wire new_AGEMA_signal_13563 ;
    wire new_AGEMA_signal_13564 ;
    wire new_AGEMA_signal_13565 ;
    wire new_AGEMA_signal_13566 ;
    wire new_AGEMA_signal_13567 ;
    wire new_AGEMA_signal_13568 ;
    wire new_AGEMA_signal_13569 ;
    wire new_AGEMA_signal_13570 ;
    wire new_AGEMA_signal_13571 ;
    wire new_AGEMA_signal_13572 ;
    wire new_AGEMA_signal_13573 ;
    wire new_AGEMA_signal_13574 ;
    wire new_AGEMA_signal_13575 ;
    wire new_AGEMA_signal_13576 ;
    wire new_AGEMA_signal_13577 ;
    wire new_AGEMA_signal_13578 ;
    wire new_AGEMA_signal_13579 ;
    wire new_AGEMA_signal_13580 ;
    wire new_AGEMA_signal_13581 ;
    wire new_AGEMA_signal_13582 ;
    wire new_AGEMA_signal_13583 ;
    wire new_AGEMA_signal_13584 ;
    wire new_AGEMA_signal_13585 ;
    wire new_AGEMA_signal_13586 ;
    wire new_AGEMA_signal_13587 ;
    wire new_AGEMA_signal_13588 ;
    wire new_AGEMA_signal_13589 ;
    wire new_AGEMA_signal_13590 ;
    wire new_AGEMA_signal_13591 ;
    wire new_AGEMA_signal_13592 ;
    wire new_AGEMA_signal_13593 ;
    wire new_AGEMA_signal_13594 ;
    wire new_AGEMA_signal_13595 ;
    wire new_AGEMA_signal_13596 ;
    wire new_AGEMA_signal_13597 ;
    wire new_AGEMA_signal_13598 ;
    wire new_AGEMA_signal_13599 ;
    wire new_AGEMA_signal_13600 ;
    wire new_AGEMA_signal_13601 ;
    wire new_AGEMA_signal_13602 ;
    wire new_AGEMA_signal_13603 ;
    wire new_AGEMA_signal_13604 ;
    wire new_AGEMA_signal_13605 ;
    wire new_AGEMA_signal_13606 ;
    wire new_AGEMA_signal_13607 ;
    wire new_AGEMA_signal_13608 ;
    wire new_AGEMA_signal_13609 ;
    wire new_AGEMA_signal_13610 ;
    wire new_AGEMA_signal_13611 ;
    wire new_AGEMA_signal_13612 ;
    wire new_AGEMA_signal_13613 ;
    wire new_AGEMA_signal_13614 ;
    wire new_AGEMA_signal_13615 ;
    wire new_AGEMA_signal_13616 ;
    wire new_AGEMA_signal_13617 ;
    wire new_AGEMA_signal_13618 ;
    wire new_AGEMA_signal_13619 ;
    wire new_AGEMA_signal_13620 ;
    wire new_AGEMA_signal_13621 ;
    wire new_AGEMA_signal_13622 ;
    wire new_AGEMA_signal_13623 ;
    wire new_AGEMA_signal_13624 ;
    wire new_AGEMA_signal_13625 ;
    wire new_AGEMA_signal_13626 ;
    wire new_AGEMA_signal_13627 ;
    wire new_AGEMA_signal_13628 ;
    wire new_AGEMA_signal_13629 ;
    wire new_AGEMA_signal_13630 ;
    wire new_AGEMA_signal_13631 ;
    wire new_AGEMA_signal_13632 ;
    wire new_AGEMA_signal_13633 ;
    wire new_AGEMA_signal_13634 ;
    wire new_AGEMA_signal_13635 ;
    wire new_AGEMA_signal_13636 ;
    wire new_AGEMA_signal_13637 ;
    wire new_AGEMA_signal_13638 ;
    wire new_AGEMA_signal_13639 ;
    wire new_AGEMA_signal_13640 ;
    wire new_AGEMA_signal_13641 ;
    wire new_AGEMA_signal_13642 ;
    wire new_AGEMA_signal_13643 ;
    wire new_AGEMA_signal_13644 ;
    wire new_AGEMA_signal_13645 ;
    wire new_AGEMA_signal_13646 ;
    wire new_AGEMA_signal_13647 ;
    wire new_AGEMA_signal_13648 ;
    wire new_AGEMA_signal_13649 ;
    wire new_AGEMA_signal_13650 ;
    wire new_AGEMA_signal_13651 ;
    wire new_AGEMA_signal_13652 ;
    wire new_AGEMA_signal_13653 ;
    wire new_AGEMA_signal_13654 ;
    wire new_AGEMA_signal_13655 ;
    wire new_AGEMA_signal_13656 ;
    wire new_AGEMA_signal_13657 ;
    wire new_AGEMA_signal_13658 ;
    wire new_AGEMA_signal_13659 ;
    wire new_AGEMA_signal_13660 ;
    wire new_AGEMA_signal_13661 ;
    wire new_AGEMA_signal_13662 ;
    wire new_AGEMA_signal_13663 ;
    wire new_AGEMA_signal_13664 ;
    wire new_AGEMA_signal_13665 ;
    wire new_AGEMA_signal_13666 ;
    wire new_AGEMA_signal_13667 ;
    wire new_AGEMA_signal_13668 ;
    wire new_AGEMA_signal_13669 ;
    wire new_AGEMA_signal_13670 ;
    wire new_AGEMA_signal_13671 ;
    wire new_AGEMA_signal_13672 ;
    wire new_AGEMA_signal_13673 ;
    wire new_AGEMA_signal_13674 ;
    wire new_AGEMA_signal_13675 ;
    wire new_AGEMA_signal_13676 ;
    wire new_AGEMA_signal_13677 ;
    wire new_AGEMA_signal_13678 ;
    wire new_AGEMA_signal_13679 ;
    wire new_AGEMA_signal_13680 ;
    wire new_AGEMA_signal_13681 ;
    wire new_AGEMA_signal_13682 ;
    wire new_AGEMA_signal_13683 ;
    wire new_AGEMA_signal_13684 ;
    wire new_AGEMA_signal_13685 ;
    wire new_AGEMA_signal_13686 ;
    wire new_AGEMA_signal_13687 ;
    wire new_AGEMA_signal_13688 ;
    wire new_AGEMA_signal_13689 ;
    wire new_AGEMA_signal_13690 ;
    wire new_AGEMA_signal_13691 ;
    wire new_AGEMA_signal_13692 ;
    wire new_AGEMA_signal_13693 ;
    wire new_AGEMA_signal_13694 ;
    wire new_AGEMA_signal_13695 ;
    wire new_AGEMA_signal_13696 ;
    wire new_AGEMA_signal_13697 ;
    wire new_AGEMA_signal_13698 ;
    wire new_AGEMA_signal_13699 ;
    wire new_AGEMA_signal_13700 ;
    wire new_AGEMA_signal_13701 ;
    wire new_AGEMA_signal_13702 ;
    wire new_AGEMA_signal_13703 ;
    wire new_AGEMA_signal_13704 ;
    wire new_AGEMA_signal_13705 ;
    wire new_AGEMA_signal_13706 ;
    wire new_AGEMA_signal_13707 ;
    wire new_AGEMA_signal_13708 ;
    wire new_AGEMA_signal_13709 ;
    wire new_AGEMA_signal_13710 ;
    wire new_AGEMA_signal_13711 ;
    wire new_AGEMA_signal_13712 ;
    wire new_AGEMA_signal_13713 ;
    wire new_AGEMA_signal_13714 ;
    wire new_AGEMA_signal_13715 ;
    wire new_AGEMA_signal_13716 ;
    wire new_AGEMA_signal_13717 ;
    wire new_AGEMA_signal_13718 ;
    wire new_AGEMA_signal_13719 ;
    wire new_AGEMA_signal_13720 ;
    wire new_AGEMA_signal_13721 ;
    wire new_AGEMA_signal_13722 ;
    wire new_AGEMA_signal_13723 ;
    wire new_AGEMA_signal_13724 ;
    wire new_AGEMA_signal_13725 ;
    wire new_AGEMA_signal_13726 ;
    wire new_AGEMA_signal_13727 ;
    wire new_AGEMA_signal_13728 ;
    wire new_AGEMA_signal_13729 ;
    wire new_AGEMA_signal_13730 ;
    wire new_AGEMA_signal_13731 ;
    wire new_AGEMA_signal_13732 ;
    wire new_AGEMA_signal_13733 ;
    wire new_AGEMA_signal_13734 ;
    wire new_AGEMA_signal_13735 ;
    wire new_AGEMA_signal_13736 ;
    wire new_AGEMA_signal_13737 ;
    wire new_AGEMA_signal_13738 ;
    wire new_AGEMA_signal_13739 ;
    wire new_AGEMA_signal_13740 ;
    wire new_AGEMA_signal_13741 ;
    wire new_AGEMA_signal_13742 ;
    wire new_AGEMA_signal_13743 ;
    wire new_AGEMA_signal_13744 ;
    wire new_AGEMA_signal_13745 ;
    wire new_AGEMA_signal_13746 ;
    wire new_AGEMA_signal_13747 ;
    wire new_AGEMA_signal_13748 ;
    wire new_AGEMA_signal_13749 ;
    wire new_AGEMA_signal_13750 ;
    wire new_AGEMA_signal_13751 ;
    wire new_AGEMA_signal_13752 ;
    wire new_AGEMA_signal_13753 ;
    wire new_AGEMA_signal_13754 ;
    wire new_AGEMA_signal_13755 ;
    wire new_AGEMA_signal_13756 ;
    wire new_AGEMA_signal_13757 ;
    wire new_AGEMA_signal_13758 ;
    wire new_AGEMA_signal_13759 ;
    wire new_AGEMA_signal_13760 ;
    wire new_AGEMA_signal_13761 ;
    wire new_AGEMA_signal_13762 ;
    wire new_AGEMA_signal_13763 ;
    wire new_AGEMA_signal_13764 ;
    wire new_AGEMA_signal_13765 ;
    wire new_AGEMA_signal_13766 ;
    wire new_AGEMA_signal_13767 ;
    wire new_AGEMA_signal_13768 ;
    wire new_AGEMA_signal_13769 ;
    wire new_AGEMA_signal_13770 ;
    wire new_AGEMA_signal_13771 ;
    wire new_AGEMA_signal_13772 ;
    wire new_AGEMA_signal_13773 ;
    wire new_AGEMA_signal_13774 ;
    wire new_AGEMA_signal_13775 ;
    wire new_AGEMA_signal_13776 ;
    wire new_AGEMA_signal_13777 ;
    wire new_AGEMA_signal_13778 ;
    wire new_AGEMA_signal_13779 ;
    wire new_AGEMA_signal_13780 ;
    wire new_AGEMA_signal_13781 ;
    wire new_AGEMA_signal_13782 ;
    wire new_AGEMA_signal_13783 ;
    wire new_AGEMA_signal_13784 ;
    wire new_AGEMA_signal_13785 ;
    wire new_AGEMA_signal_13786 ;
    wire new_AGEMA_signal_13787 ;
    wire new_AGEMA_signal_13788 ;
    wire new_AGEMA_signal_13789 ;
    wire new_AGEMA_signal_13790 ;
    wire new_AGEMA_signal_13791 ;
    wire new_AGEMA_signal_13792 ;
    wire new_AGEMA_signal_13793 ;
    wire new_AGEMA_signal_13794 ;
    wire new_AGEMA_signal_13795 ;
    wire new_AGEMA_signal_13796 ;
    wire new_AGEMA_signal_13797 ;
    wire new_AGEMA_signal_13798 ;
    wire new_AGEMA_signal_13799 ;
    wire new_AGEMA_signal_13800 ;
    wire new_AGEMA_signal_13801 ;
    wire new_AGEMA_signal_13802 ;
    wire new_AGEMA_signal_13803 ;
    wire new_AGEMA_signal_13804 ;
    wire new_AGEMA_signal_13805 ;
    wire new_AGEMA_signal_13806 ;
    wire new_AGEMA_signal_13807 ;
    wire new_AGEMA_signal_13808 ;
    wire new_AGEMA_signal_13809 ;
    wire new_AGEMA_signal_13810 ;
    wire new_AGEMA_signal_13811 ;
    wire new_AGEMA_signal_13812 ;
    wire new_AGEMA_signal_13813 ;
    wire new_AGEMA_signal_13814 ;
    wire new_AGEMA_signal_13815 ;
    wire new_AGEMA_signal_13816 ;
    wire new_AGEMA_signal_13817 ;
    wire new_AGEMA_signal_13818 ;
    wire new_AGEMA_signal_13819 ;
    wire new_AGEMA_signal_13820 ;
    wire new_AGEMA_signal_13821 ;
    wire new_AGEMA_signal_13822 ;
    wire new_AGEMA_signal_13823 ;
    wire new_AGEMA_signal_13824 ;
    wire new_AGEMA_signal_13825 ;
    wire new_AGEMA_signal_13826 ;
    wire new_AGEMA_signal_13827 ;
    wire new_AGEMA_signal_13828 ;
    wire new_AGEMA_signal_13829 ;
    wire new_AGEMA_signal_13830 ;
    wire new_AGEMA_signal_13831 ;
    wire new_AGEMA_signal_13832 ;
    wire new_AGEMA_signal_13833 ;
    wire new_AGEMA_signal_13834 ;
    wire new_AGEMA_signal_13835 ;
    wire new_AGEMA_signal_13836 ;
    wire new_AGEMA_signal_13837 ;
    wire new_AGEMA_signal_13838 ;
    wire new_AGEMA_signal_13839 ;
    wire new_AGEMA_signal_13840 ;
    wire new_AGEMA_signal_13841 ;
    wire new_AGEMA_signal_13842 ;
    wire new_AGEMA_signal_13843 ;
    wire new_AGEMA_signal_13844 ;
    wire new_AGEMA_signal_13845 ;
    wire new_AGEMA_signal_13846 ;
    wire new_AGEMA_signal_13847 ;
    wire new_AGEMA_signal_13848 ;
    wire new_AGEMA_signal_13849 ;
    wire new_AGEMA_signal_13850 ;
    wire new_AGEMA_signal_13851 ;
    wire new_AGEMA_signal_13852 ;
    wire new_AGEMA_signal_13853 ;
    wire new_AGEMA_signal_13854 ;
    wire new_AGEMA_signal_13855 ;
    wire new_AGEMA_signal_13856 ;
    wire new_AGEMA_signal_13857 ;
    wire new_AGEMA_signal_13858 ;
    wire new_AGEMA_signal_13859 ;
    wire new_AGEMA_signal_13860 ;
    wire new_AGEMA_signal_13861 ;
    wire new_AGEMA_signal_13862 ;
    wire new_AGEMA_signal_13863 ;
    wire new_AGEMA_signal_13864 ;
    wire new_AGEMA_signal_13865 ;
    wire new_AGEMA_signal_13866 ;
    wire new_AGEMA_signal_13867 ;
    wire new_AGEMA_signal_13868 ;
    wire new_AGEMA_signal_13869 ;
    wire new_AGEMA_signal_13870 ;
    wire new_AGEMA_signal_13871 ;
    wire new_AGEMA_signal_13872 ;
    wire new_AGEMA_signal_13873 ;
    wire new_AGEMA_signal_13874 ;
    wire new_AGEMA_signal_13875 ;
    wire new_AGEMA_signal_13876 ;
    wire new_AGEMA_signal_13877 ;
    wire new_AGEMA_signal_13878 ;
    wire new_AGEMA_signal_13879 ;
    wire new_AGEMA_signal_13880 ;
    wire new_AGEMA_signal_13881 ;
    wire new_AGEMA_signal_13882 ;
    wire new_AGEMA_signal_13883 ;
    wire new_AGEMA_signal_13884 ;
    wire new_AGEMA_signal_13885 ;
    wire new_AGEMA_signal_13886 ;
    wire new_AGEMA_signal_13887 ;
    wire new_AGEMA_signal_13888 ;
    wire new_AGEMA_signal_13889 ;
    wire new_AGEMA_signal_13890 ;
    wire new_AGEMA_signal_13891 ;
    wire new_AGEMA_signal_13892 ;
    wire new_AGEMA_signal_13893 ;
    wire new_AGEMA_signal_13894 ;
    wire new_AGEMA_signal_13895 ;
    wire new_AGEMA_signal_13896 ;
    wire new_AGEMA_signal_13897 ;
    wire new_AGEMA_signal_13898 ;
    wire new_AGEMA_signal_13899 ;
    wire new_AGEMA_signal_13900 ;
    wire new_AGEMA_signal_13901 ;
    wire new_AGEMA_signal_13902 ;
    wire new_AGEMA_signal_13903 ;
    wire new_AGEMA_signal_13904 ;
    wire new_AGEMA_signal_13905 ;
    wire new_AGEMA_signal_13906 ;
    wire new_AGEMA_signal_13907 ;
    wire new_AGEMA_signal_13908 ;
    wire new_AGEMA_signal_13909 ;
    wire new_AGEMA_signal_13910 ;
    wire new_AGEMA_signal_13911 ;
    wire new_AGEMA_signal_13912 ;
    wire new_AGEMA_signal_13913 ;
    wire new_AGEMA_signal_13914 ;
    wire new_AGEMA_signal_13915 ;
    wire new_AGEMA_signal_13916 ;
    wire new_AGEMA_signal_13917 ;
    wire new_AGEMA_signal_13918 ;
    wire new_AGEMA_signal_13919 ;
    wire new_AGEMA_signal_13920 ;
    wire new_AGEMA_signal_13921 ;
    wire new_AGEMA_signal_13922 ;
    wire new_AGEMA_signal_13923 ;
    wire new_AGEMA_signal_13924 ;
    wire new_AGEMA_signal_13925 ;
    wire new_AGEMA_signal_13926 ;
    wire new_AGEMA_signal_13927 ;
    wire new_AGEMA_signal_13928 ;
    wire new_AGEMA_signal_13929 ;
    wire new_AGEMA_signal_13930 ;
    wire new_AGEMA_signal_13931 ;
    wire new_AGEMA_signal_13932 ;
    wire new_AGEMA_signal_13933 ;
    wire new_AGEMA_signal_13934 ;
    wire new_AGEMA_signal_13935 ;
    wire new_AGEMA_signal_13936 ;
    wire new_AGEMA_signal_13937 ;
    wire new_AGEMA_signal_13938 ;
    wire new_AGEMA_signal_13939 ;
    wire new_AGEMA_signal_13940 ;
    wire new_AGEMA_signal_13941 ;
    wire new_AGEMA_signal_13942 ;
    wire new_AGEMA_signal_13943 ;
    wire new_AGEMA_signal_13944 ;
    wire new_AGEMA_signal_13945 ;
    wire new_AGEMA_signal_13946 ;
    wire new_AGEMA_signal_13947 ;
    wire new_AGEMA_signal_13948 ;
    wire new_AGEMA_signal_13949 ;
    wire new_AGEMA_signal_13950 ;
    wire new_AGEMA_signal_13951 ;
    wire new_AGEMA_signal_13952 ;
    wire new_AGEMA_signal_13953 ;
    wire new_AGEMA_signal_13954 ;
    wire new_AGEMA_signal_13955 ;
    wire new_AGEMA_signal_13956 ;
    wire new_AGEMA_signal_13957 ;
    wire new_AGEMA_signal_13958 ;
    wire new_AGEMA_signal_13959 ;
    wire new_AGEMA_signal_13960 ;
    wire new_AGEMA_signal_13961 ;
    wire new_AGEMA_signal_13962 ;
    wire new_AGEMA_signal_13963 ;
    wire new_AGEMA_signal_13964 ;
    wire new_AGEMA_signal_13965 ;
    wire new_AGEMA_signal_13966 ;
    wire new_AGEMA_signal_13967 ;
    wire new_AGEMA_signal_13968 ;
    wire new_AGEMA_signal_13969 ;
    wire new_AGEMA_signal_13970 ;
    wire new_AGEMA_signal_13971 ;
    wire new_AGEMA_signal_13972 ;
    wire new_AGEMA_signal_13973 ;
    wire new_AGEMA_signal_13974 ;
    wire new_AGEMA_signal_13975 ;
    wire new_AGEMA_signal_13976 ;
    wire new_AGEMA_signal_13977 ;
    wire new_AGEMA_signal_13978 ;
    wire new_AGEMA_signal_13979 ;
    wire new_AGEMA_signal_13980 ;
    wire new_AGEMA_signal_13981 ;
    wire new_AGEMA_signal_13982 ;
    wire new_AGEMA_signal_13983 ;
    wire new_AGEMA_signal_13984 ;
    wire new_AGEMA_signal_13985 ;
    wire new_AGEMA_signal_13986 ;
    wire new_AGEMA_signal_13987 ;
    wire new_AGEMA_signal_13988 ;
    wire new_AGEMA_signal_13989 ;
    wire new_AGEMA_signal_13990 ;
    wire new_AGEMA_signal_13991 ;
    wire new_AGEMA_signal_13992 ;
    wire new_AGEMA_signal_13993 ;
    wire new_AGEMA_signal_13994 ;
    wire new_AGEMA_signal_13995 ;
    wire new_AGEMA_signal_13996 ;
    wire new_AGEMA_signal_13997 ;
    wire new_AGEMA_signal_13998 ;
    wire new_AGEMA_signal_13999 ;
    wire new_AGEMA_signal_14000 ;
    wire new_AGEMA_signal_14001 ;
    wire new_AGEMA_signal_14002 ;
    wire new_AGEMA_signal_14003 ;
    wire new_AGEMA_signal_14004 ;
    wire new_AGEMA_signal_14005 ;
    wire new_AGEMA_signal_14006 ;
    wire new_AGEMA_signal_14007 ;
    wire new_AGEMA_signal_14008 ;
    wire new_AGEMA_signal_14009 ;
    wire new_AGEMA_signal_14010 ;
    wire new_AGEMA_signal_14011 ;
    wire new_AGEMA_signal_14012 ;
    wire new_AGEMA_signal_14013 ;
    wire new_AGEMA_signal_14014 ;
    wire new_AGEMA_signal_14015 ;
    wire new_AGEMA_signal_14016 ;
    wire new_AGEMA_signal_14017 ;
    wire new_AGEMA_signal_14018 ;
    wire new_AGEMA_signal_14019 ;
    wire new_AGEMA_signal_14020 ;
    wire new_AGEMA_signal_14021 ;
    wire new_AGEMA_signal_14022 ;
    wire new_AGEMA_signal_14023 ;
    wire new_AGEMA_signal_14024 ;
    wire new_AGEMA_signal_14025 ;
    wire new_AGEMA_signal_14026 ;
    wire new_AGEMA_signal_14027 ;
    wire new_AGEMA_signal_14028 ;
    wire new_AGEMA_signal_14029 ;
    wire new_AGEMA_signal_14030 ;
    wire new_AGEMA_signal_14031 ;
    wire new_AGEMA_signal_14032 ;
    wire new_AGEMA_signal_14033 ;
    wire new_AGEMA_signal_14034 ;
    wire new_AGEMA_signal_14035 ;
    wire new_AGEMA_signal_14036 ;
    wire new_AGEMA_signal_14037 ;
    wire new_AGEMA_signal_14038 ;
    wire new_AGEMA_signal_14039 ;
    wire new_AGEMA_signal_14040 ;
    wire new_AGEMA_signal_14041 ;
    wire new_AGEMA_signal_14042 ;
    wire new_AGEMA_signal_14043 ;
    wire new_AGEMA_signal_14044 ;
    wire new_AGEMA_signal_14045 ;
    wire new_AGEMA_signal_14046 ;
    wire new_AGEMA_signal_14047 ;
    wire new_AGEMA_signal_14048 ;
    wire new_AGEMA_signal_14049 ;
    wire new_AGEMA_signal_14050 ;
    wire new_AGEMA_signal_14051 ;
    wire new_AGEMA_signal_14052 ;
    wire new_AGEMA_signal_14053 ;
    wire new_AGEMA_signal_14054 ;
    wire new_AGEMA_signal_14055 ;
    wire new_AGEMA_signal_14056 ;
    wire new_AGEMA_signal_14057 ;
    wire new_AGEMA_signal_14058 ;
    wire new_AGEMA_signal_14059 ;
    wire new_AGEMA_signal_14060 ;
    wire new_AGEMA_signal_14061 ;
    wire new_AGEMA_signal_14062 ;
    wire new_AGEMA_signal_14063 ;
    wire new_AGEMA_signal_14064 ;
    wire new_AGEMA_signal_14065 ;
    wire new_AGEMA_signal_14066 ;
    wire new_AGEMA_signal_14067 ;
    wire new_AGEMA_signal_14068 ;
    wire new_AGEMA_signal_14069 ;
    wire new_AGEMA_signal_14070 ;
    wire new_AGEMA_signal_14071 ;
    wire new_AGEMA_signal_14072 ;
    wire new_AGEMA_signal_14073 ;
    wire new_AGEMA_signal_14074 ;
    wire new_AGEMA_signal_14075 ;
    wire new_AGEMA_signal_14076 ;
    wire new_AGEMA_signal_14077 ;
    wire new_AGEMA_signal_14078 ;
    wire new_AGEMA_signal_14079 ;
    wire new_AGEMA_signal_14080 ;
    wire new_AGEMA_signal_14081 ;
    wire new_AGEMA_signal_14082 ;
    wire new_AGEMA_signal_14083 ;
    wire new_AGEMA_signal_14084 ;
    wire new_AGEMA_signal_14085 ;
    wire new_AGEMA_signal_14086 ;
    wire new_AGEMA_signal_14087 ;
    wire new_AGEMA_signal_14088 ;
    wire new_AGEMA_signal_14089 ;
    wire new_AGEMA_signal_14090 ;
    wire new_AGEMA_signal_14091 ;
    wire new_AGEMA_signal_14092 ;
    wire new_AGEMA_signal_14093 ;
    wire new_AGEMA_signal_14094 ;
    wire new_AGEMA_signal_14095 ;
    wire new_AGEMA_signal_14096 ;
    wire new_AGEMA_signal_14097 ;
    wire new_AGEMA_signal_14098 ;
    wire new_AGEMA_signal_14099 ;
    wire new_AGEMA_signal_14100 ;
    wire new_AGEMA_signal_14101 ;
    wire new_AGEMA_signal_14102 ;
    wire new_AGEMA_signal_14103 ;
    wire new_AGEMA_signal_14104 ;
    wire new_AGEMA_signal_14105 ;
    wire new_AGEMA_signal_14106 ;
    wire new_AGEMA_signal_14107 ;
    wire new_AGEMA_signal_14108 ;
    wire new_AGEMA_signal_14109 ;
    wire new_AGEMA_signal_14110 ;
    wire new_AGEMA_signal_14111 ;
    wire new_AGEMA_signal_14112 ;
    wire new_AGEMA_signal_14113 ;
    wire new_AGEMA_signal_14114 ;
    wire new_AGEMA_signal_14115 ;
    wire new_AGEMA_signal_14116 ;
    wire new_AGEMA_signal_14117 ;
    wire new_AGEMA_signal_14118 ;
    wire new_AGEMA_signal_14119 ;
    wire new_AGEMA_signal_14120 ;
    wire new_AGEMA_signal_14121 ;
    wire new_AGEMA_signal_14122 ;
    wire new_AGEMA_signal_14123 ;
    wire new_AGEMA_signal_14124 ;
    wire new_AGEMA_signal_14125 ;
    wire new_AGEMA_signal_14126 ;
    wire new_AGEMA_signal_14127 ;
    wire new_AGEMA_signal_14128 ;
    wire new_AGEMA_signal_14129 ;
    wire new_AGEMA_signal_14130 ;
    wire new_AGEMA_signal_14131 ;
    wire new_AGEMA_signal_14132 ;
    wire new_AGEMA_signal_14133 ;
    wire new_AGEMA_signal_14134 ;
    wire new_AGEMA_signal_14135 ;
    wire new_AGEMA_signal_14136 ;
    wire new_AGEMA_signal_14137 ;
    wire new_AGEMA_signal_14138 ;
    wire new_AGEMA_signal_14139 ;
    wire new_AGEMA_signal_14140 ;
    wire new_AGEMA_signal_14141 ;
    wire new_AGEMA_signal_14142 ;
    wire new_AGEMA_signal_14143 ;
    wire new_AGEMA_signal_14144 ;
    wire new_AGEMA_signal_14145 ;
    wire new_AGEMA_signal_14146 ;
    wire new_AGEMA_signal_14147 ;
    wire new_AGEMA_signal_14148 ;
    wire new_AGEMA_signal_14149 ;
    wire new_AGEMA_signal_14150 ;
    wire new_AGEMA_signal_14151 ;
    wire new_AGEMA_signal_14152 ;
    wire new_AGEMA_signal_14153 ;
    wire new_AGEMA_signal_14154 ;
    wire new_AGEMA_signal_14155 ;
    wire new_AGEMA_signal_14156 ;
    wire new_AGEMA_signal_14157 ;
    wire new_AGEMA_signal_14158 ;
    wire new_AGEMA_signal_14159 ;
    wire new_AGEMA_signal_14160 ;
    wire new_AGEMA_signal_14161 ;
    wire new_AGEMA_signal_14162 ;
    wire new_AGEMA_signal_14163 ;
    wire new_AGEMA_signal_14164 ;
    wire new_AGEMA_signal_14165 ;
    wire new_AGEMA_signal_14166 ;
    wire new_AGEMA_signal_14167 ;
    wire new_AGEMA_signal_14168 ;
    wire new_AGEMA_signal_14169 ;
    wire new_AGEMA_signal_14170 ;
    wire new_AGEMA_signal_14171 ;
    wire new_AGEMA_signal_14172 ;
    wire new_AGEMA_signal_14173 ;
    wire new_AGEMA_signal_14174 ;
    wire new_AGEMA_signal_14175 ;
    wire new_AGEMA_signal_14176 ;
    wire new_AGEMA_signal_14177 ;
    wire new_AGEMA_signal_14178 ;
    wire new_AGEMA_signal_14179 ;
    wire new_AGEMA_signal_14180 ;
    wire new_AGEMA_signal_14181 ;
    wire new_AGEMA_signal_14182 ;
    wire new_AGEMA_signal_14183 ;
    wire new_AGEMA_signal_14184 ;
    wire new_AGEMA_signal_14185 ;
    wire new_AGEMA_signal_14186 ;
    wire new_AGEMA_signal_14187 ;
    wire new_AGEMA_signal_14188 ;
    wire new_AGEMA_signal_14189 ;
    wire new_AGEMA_signal_14190 ;
    wire new_AGEMA_signal_14191 ;
    wire new_AGEMA_signal_14192 ;
    wire new_AGEMA_signal_14193 ;
    wire new_AGEMA_signal_14194 ;
    wire new_AGEMA_signal_14195 ;
    wire new_AGEMA_signal_14196 ;
    wire new_AGEMA_signal_14197 ;
    wire new_AGEMA_signal_14198 ;
    wire new_AGEMA_signal_14199 ;
    wire new_AGEMA_signal_14200 ;
    wire new_AGEMA_signal_14201 ;
    wire new_AGEMA_signal_14202 ;
    wire new_AGEMA_signal_14203 ;
    wire new_AGEMA_signal_14204 ;
    wire new_AGEMA_signal_14205 ;
    wire new_AGEMA_signal_14206 ;
    wire new_AGEMA_signal_14207 ;
    wire new_AGEMA_signal_14208 ;
    wire new_AGEMA_signal_14209 ;
    wire new_AGEMA_signal_14210 ;
    wire new_AGEMA_signal_14211 ;
    wire new_AGEMA_signal_14212 ;
    wire new_AGEMA_signal_14213 ;
    wire new_AGEMA_signal_14214 ;
    wire new_AGEMA_signal_14215 ;
    wire new_AGEMA_signal_14216 ;
    wire new_AGEMA_signal_14217 ;
    wire new_AGEMA_signal_14218 ;
    wire new_AGEMA_signal_14219 ;
    wire new_AGEMA_signal_14220 ;
    wire new_AGEMA_signal_14221 ;
    wire new_AGEMA_signal_14222 ;
    wire new_AGEMA_signal_14223 ;
    wire new_AGEMA_signal_14224 ;
    wire new_AGEMA_signal_14225 ;
    wire new_AGEMA_signal_14226 ;
    wire new_AGEMA_signal_14227 ;
    wire new_AGEMA_signal_14228 ;
    wire new_AGEMA_signal_14229 ;
    wire new_AGEMA_signal_14230 ;
    wire new_AGEMA_signal_14231 ;
    wire new_AGEMA_signal_14232 ;
    wire new_AGEMA_signal_14233 ;
    wire new_AGEMA_signal_14234 ;
    wire new_AGEMA_signal_14235 ;
    wire new_AGEMA_signal_14236 ;
    wire new_AGEMA_signal_14237 ;
    wire new_AGEMA_signal_14238 ;
    wire new_AGEMA_signal_14239 ;
    wire new_AGEMA_signal_14240 ;
    wire new_AGEMA_signal_14241 ;
    wire new_AGEMA_signal_14242 ;
    wire new_AGEMA_signal_14243 ;
    wire new_AGEMA_signal_14244 ;
    wire new_AGEMA_signal_14245 ;
    wire new_AGEMA_signal_14246 ;
    wire new_AGEMA_signal_14247 ;
    wire new_AGEMA_signal_14248 ;
    wire new_AGEMA_signal_14249 ;
    wire new_AGEMA_signal_14250 ;
    wire new_AGEMA_signal_14251 ;
    wire new_AGEMA_signal_14252 ;
    wire new_AGEMA_signal_14253 ;
    wire new_AGEMA_signal_14254 ;
    wire new_AGEMA_signal_14255 ;
    wire new_AGEMA_signal_14256 ;
    wire new_AGEMA_signal_14257 ;
    wire new_AGEMA_signal_14258 ;
    wire new_AGEMA_signal_14259 ;
    wire new_AGEMA_signal_14260 ;
    wire new_AGEMA_signal_14261 ;
    wire new_AGEMA_signal_14262 ;
    wire new_AGEMA_signal_14263 ;
    wire new_AGEMA_signal_14264 ;
    wire new_AGEMA_signal_14265 ;
    wire new_AGEMA_signal_14266 ;
    wire new_AGEMA_signal_14267 ;
    wire new_AGEMA_signal_14268 ;
    wire new_AGEMA_signal_14269 ;
    wire new_AGEMA_signal_14270 ;
    wire new_AGEMA_signal_14271 ;
    wire new_AGEMA_signal_14272 ;
    wire new_AGEMA_signal_14273 ;
    wire new_AGEMA_signal_14274 ;
    wire new_AGEMA_signal_14275 ;
    wire new_AGEMA_signal_14276 ;
    wire new_AGEMA_signal_14277 ;
    wire new_AGEMA_signal_14278 ;
    wire new_AGEMA_signal_14279 ;
    wire new_AGEMA_signal_14280 ;
    wire new_AGEMA_signal_14281 ;
    wire new_AGEMA_signal_14282 ;
    wire new_AGEMA_signal_14283 ;
    wire new_AGEMA_signal_14284 ;
    wire new_AGEMA_signal_14285 ;
    wire new_AGEMA_signal_14286 ;
    wire new_AGEMA_signal_14287 ;
    wire new_AGEMA_signal_14288 ;
    wire new_AGEMA_signal_14289 ;
    wire new_AGEMA_signal_14290 ;
    wire new_AGEMA_signal_14291 ;
    wire new_AGEMA_signal_14292 ;
    wire new_AGEMA_signal_14293 ;
    wire new_AGEMA_signal_14294 ;
    wire new_AGEMA_signal_14295 ;
    wire new_AGEMA_signal_14296 ;
    wire new_AGEMA_signal_14297 ;
    wire new_AGEMA_signal_14298 ;
    wire new_AGEMA_signal_14299 ;
    wire new_AGEMA_signal_14300 ;
    wire new_AGEMA_signal_14301 ;
    wire new_AGEMA_signal_14302 ;
    wire new_AGEMA_signal_14303 ;
    wire new_AGEMA_signal_14304 ;
    wire new_AGEMA_signal_14305 ;
    wire new_AGEMA_signal_14306 ;
    wire new_AGEMA_signal_14307 ;
    wire new_AGEMA_signal_14308 ;
    wire new_AGEMA_signal_14309 ;
    wire new_AGEMA_signal_14310 ;
    wire new_AGEMA_signal_14311 ;
    wire new_AGEMA_signal_14312 ;
    wire new_AGEMA_signal_14313 ;
    wire new_AGEMA_signal_14314 ;
    wire new_AGEMA_signal_14315 ;
    wire new_AGEMA_signal_14316 ;
    wire new_AGEMA_signal_14317 ;
    wire new_AGEMA_signal_14318 ;
    wire new_AGEMA_signal_14319 ;
    wire new_AGEMA_signal_14320 ;
    wire new_AGEMA_signal_14321 ;
    wire new_AGEMA_signal_14322 ;
    wire new_AGEMA_signal_14323 ;
    wire new_AGEMA_signal_14324 ;
    wire new_AGEMA_signal_14325 ;
    wire new_AGEMA_signal_14326 ;
    wire new_AGEMA_signal_14327 ;
    wire new_AGEMA_signal_14328 ;
    wire new_AGEMA_signal_14329 ;
    wire new_AGEMA_signal_14330 ;
    wire new_AGEMA_signal_14331 ;
    wire new_AGEMA_signal_14332 ;
    wire new_AGEMA_signal_14333 ;
    wire new_AGEMA_signal_14334 ;
    wire new_AGEMA_signal_14335 ;
    wire new_AGEMA_signal_14336 ;
    wire new_AGEMA_signal_14337 ;
    wire new_AGEMA_signal_14338 ;
    wire new_AGEMA_signal_14339 ;
    wire new_AGEMA_signal_14340 ;
    wire new_AGEMA_signal_14341 ;
    wire new_AGEMA_signal_14342 ;
    wire new_AGEMA_signal_14343 ;
    wire new_AGEMA_signal_14344 ;
    wire new_AGEMA_signal_14345 ;
    wire new_AGEMA_signal_14346 ;
    wire new_AGEMA_signal_14347 ;
    wire new_AGEMA_signal_14348 ;
    wire new_AGEMA_signal_14349 ;
    wire new_AGEMA_signal_14350 ;
    wire new_AGEMA_signal_14351 ;
    wire new_AGEMA_signal_14352 ;
    wire new_AGEMA_signal_14353 ;
    wire new_AGEMA_signal_14354 ;
    wire new_AGEMA_signal_14355 ;
    wire new_AGEMA_signal_14356 ;
    wire new_AGEMA_signal_14357 ;
    wire new_AGEMA_signal_14358 ;
    wire new_AGEMA_signal_14359 ;
    wire new_AGEMA_signal_14360 ;
    wire new_AGEMA_signal_14361 ;
    wire new_AGEMA_signal_14362 ;
    wire new_AGEMA_signal_14363 ;
    wire new_AGEMA_signal_14364 ;
    wire new_AGEMA_signal_14365 ;
    wire new_AGEMA_signal_14366 ;
    wire new_AGEMA_signal_14367 ;
    wire new_AGEMA_signal_14368 ;
    wire new_AGEMA_signal_14369 ;
    wire new_AGEMA_signal_14370 ;
    wire new_AGEMA_signal_14371 ;
    wire new_AGEMA_signal_14372 ;
    wire new_AGEMA_signal_14373 ;
    wire new_AGEMA_signal_14374 ;
    wire new_AGEMA_signal_14375 ;
    wire new_AGEMA_signal_14376 ;
    wire new_AGEMA_signal_14377 ;
    wire new_AGEMA_signal_14378 ;
    wire new_AGEMA_signal_14379 ;
    wire new_AGEMA_signal_14380 ;
    wire new_AGEMA_signal_14381 ;
    wire new_AGEMA_signal_14382 ;
    wire new_AGEMA_signal_14383 ;
    wire new_AGEMA_signal_14384 ;
    wire new_AGEMA_signal_14385 ;
    wire new_AGEMA_signal_14386 ;
    wire new_AGEMA_signal_14387 ;
    wire new_AGEMA_signal_14388 ;
    wire new_AGEMA_signal_14389 ;
    wire new_AGEMA_signal_14390 ;
    wire new_AGEMA_signal_14391 ;
    wire new_AGEMA_signal_14392 ;
    wire new_AGEMA_signal_14393 ;
    wire new_AGEMA_signal_14394 ;
    wire new_AGEMA_signal_14395 ;
    wire new_AGEMA_signal_14396 ;
    wire new_AGEMA_signal_14397 ;
    wire new_AGEMA_signal_14398 ;
    wire new_AGEMA_signal_14399 ;
    wire new_AGEMA_signal_14400 ;
    wire new_AGEMA_signal_14401 ;
    wire new_AGEMA_signal_14402 ;
    wire new_AGEMA_signal_14403 ;
    wire new_AGEMA_signal_14404 ;
    wire new_AGEMA_signal_14405 ;
    wire new_AGEMA_signal_14406 ;
    wire new_AGEMA_signal_14407 ;
    wire new_AGEMA_signal_14408 ;
    wire new_AGEMA_signal_14409 ;
    wire new_AGEMA_signal_14410 ;
    wire new_AGEMA_signal_14411 ;
    wire new_AGEMA_signal_14412 ;
    wire new_AGEMA_signal_14413 ;
    wire new_AGEMA_signal_14414 ;
    wire new_AGEMA_signal_14415 ;
    wire new_AGEMA_signal_14416 ;
    wire new_AGEMA_signal_14417 ;
    wire new_AGEMA_signal_14418 ;
    wire new_AGEMA_signal_14419 ;
    wire new_AGEMA_signal_14420 ;
    wire new_AGEMA_signal_14421 ;
    wire new_AGEMA_signal_14422 ;
    wire new_AGEMA_signal_14423 ;
    wire new_AGEMA_signal_14424 ;
    wire new_AGEMA_signal_14425 ;
    wire new_AGEMA_signal_14426 ;
    wire new_AGEMA_signal_14427 ;
    wire new_AGEMA_signal_14428 ;
    wire new_AGEMA_signal_14429 ;
    wire new_AGEMA_signal_14430 ;
    wire new_AGEMA_signal_14431 ;
    wire new_AGEMA_signal_14432 ;
    wire new_AGEMA_signal_14433 ;
    wire new_AGEMA_signal_14434 ;
    wire new_AGEMA_signal_14435 ;
    wire new_AGEMA_signal_14436 ;
    wire new_AGEMA_signal_14437 ;
    wire new_AGEMA_signal_14438 ;
    wire new_AGEMA_signal_14439 ;
    wire new_AGEMA_signal_14440 ;
    wire new_AGEMA_signal_14441 ;
    wire new_AGEMA_signal_14442 ;
    wire new_AGEMA_signal_14443 ;
    wire new_AGEMA_signal_14444 ;
    wire new_AGEMA_signal_14445 ;
    wire new_AGEMA_signal_14446 ;
    wire new_AGEMA_signal_14447 ;
    wire new_AGEMA_signal_14448 ;
    wire new_AGEMA_signal_14449 ;
    wire new_AGEMA_signal_14450 ;
    wire new_AGEMA_signal_14451 ;
    wire new_AGEMA_signal_14452 ;
    wire new_AGEMA_signal_14453 ;
    wire new_AGEMA_signal_14454 ;
    wire new_AGEMA_signal_14455 ;
    wire new_AGEMA_signal_14456 ;
    wire new_AGEMA_signal_14457 ;
    wire new_AGEMA_signal_14458 ;
    wire new_AGEMA_signal_14459 ;
    wire new_AGEMA_signal_14460 ;
    wire new_AGEMA_signal_14461 ;
    wire new_AGEMA_signal_14462 ;
    wire new_AGEMA_signal_14463 ;
    wire new_AGEMA_signal_14464 ;
    wire new_AGEMA_signal_14465 ;
    wire new_AGEMA_signal_14466 ;
    wire new_AGEMA_signal_14467 ;
    wire new_AGEMA_signal_14468 ;
    wire new_AGEMA_signal_14469 ;
    wire new_AGEMA_signal_14470 ;
    wire new_AGEMA_signal_14471 ;
    wire new_AGEMA_signal_14472 ;
    wire new_AGEMA_signal_14473 ;
    wire new_AGEMA_signal_14474 ;
    wire new_AGEMA_signal_14475 ;
    wire new_AGEMA_signal_14476 ;
    wire new_AGEMA_signal_14477 ;
    wire new_AGEMA_signal_14478 ;
    wire new_AGEMA_signal_14479 ;
    wire new_AGEMA_signal_14480 ;
    wire new_AGEMA_signal_14481 ;
    wire new_AGEMA_signal_14482 ;
    wire new_AGEMA_signal_14483 ;
    wire new_AGEMA_signal_14484 ;
    wire new_AGEMA_signal_14485 ;
    wire new_AGEMA_signal_14486 ;
    wire new_AGEMA_signal_14487 ;
    wire new_AGEMA_signal_14488 ;
    wire new_AGEMA_signal_14489 ;
    wire new_AGEMA_signal_14490 ;
    wire new_AGEMA_signal_14491 ;
    wire new_AGEMA_signal_14492 ;
    wire new_AGEMA_signal_14493 ;
    wire new_AGEMA_signal_14494 ;
    wire new_AGEMA_signal_14495 ;
    wire new_AGEMA_signal_14496 ;
    wire new_AGEMA_signal_14497 ;
    wire new_AGEMA_signal_14498 ;
    wire new_AGEMA_signal_14499 ;
    wire new_AGEMA_signal_14500 ;
    wire new_AGEMA_signal_14501 ;
    wire new_AGEMA_signal_14502 ;
    wire new_AGEMA_signal_14503 ;
    wire new_AGEMA_signal_14504 ;
    wire new_AGEMA_signal_14505 ;
    wire new_AGEMA_signal_14506 ;
    wire new_AGEMA_signal_14507 ;
    wire new_AGEMA_signal_14508 ;
    wire new_AGEMA_signal_14509 ;
    wire new_AGEMA_signal_14510 ;
    wire new_AGEMA_signal_14511 ;
    wire new_AGEMA_signal_14512 ;
    wire new_AGEMA_signal_14513 ;
    wire new_AGEMA_signal_14514 ;
    wire new_AGEMA_signal_14515 ;
    wire new_AGEMA_signal_14516 ;
    wire new_AGEMA_signal_14517 ;
    wire new_AGEMA_signal_14518 ;
    wire new_AGEMA_signal_14519 ;
    wire new_AGEMA_signal_14520 ;
    wire new_AGEMA_signal_14521 ;
    wire new_AGEMA_signal_14522 ;
    wire new_AGEMA_signal_14523 ;
    wire new_AGEMA_signal_14524 ;
    wire new_AGEMA_signal_14525 ;
    wire new_AGEMA_signal_14526 ;
    wire new_AGEMA_signal_14527 ;
    wire new_AGEMA_signal_14528 ;
    wire new_AGEMA_signal_14529 ;
    wire new_AGEMA_signal_14530 ;
    wire new_AGEMA_signal_14531 ;
    wire new_AGEMA_signal_14532 ;
    wire new_AGEMA_signal_14533 ;
    wire new_AGEMA_signal_14534 ;
    wire new_AGEMA_signal_14535 ;
    wire new_AGEMA_signal_14536 ;
    wire new_AGEMA_signal_14537 ;
    wire new_AGEMA_signal_14538 ;
    wire new_AGEMA_signal_14539 ;
    wire new_AGEMA_signal_14540 ;
    wire new_AGEMA_signal_14541 ;
    wire new_AGEMA_signal_14542 ;
    wire new_AGEMA_signal_14543 ;
    wire new_AGEMA_signal_14544 ;
    wire new_AGEMA_signal_14545 ;
    wire new_AGEMA_signal_14546 ;
    wire new_AGEMA_signal_14547 ;
    wire new_AGEMA_signal_14548 ;
    wire new_AGEMA_signal_14549 ;
    wire new_AGEMA_signal_14550 ;
    wire new_AGEMA_signal_14551 ;
    wire new_AGEMA_signal_14552 ;
    wire new_AGEMA_signal_14553 ;
    wire new_AGEMA_signal_14554 ;
    wire new_AGEMA_signal_14555 ;
    wire new_AGEMA_signal_14556 ;
    wire new_AGEMA_signal_14557 ;
    wire new_AGEMA_signal_14558 ;
    wire new_AGEMA_signal_14559 ;
    wire new_AGEMA_signal_14560 ;
    wire new_AGEMA_signal_14561 ;
    wire new_AGEMA_signal_14562 ;
    wire new_AGEMA_signal_14563 ;
    wire new_AGEMA_signal_14564 ;
    wire new_AGEMA_signal_14565 ;
    wire new_AGEMA_signal_14566 ;
    wire new_AGEMA_signal_14567 ;
    wire new_AGEMA_signal_14568 ;
    wire new_AGEMA_signal_14569 ;
    wire new_AGEMA_signal_14570 ;
    wire new_AGEMA_signal_14571 ;
    wire new_AGEMA_signal_14572 ;
    wire new_AGEMA_signal_14573 ;
    wire new_AGEMA_signal_14574 ;
    wire new_AGEMA_signal_14575 ;
    wire new_AGEMA_signal_14576 ;
    wire new_AGEMA_signal_14577 ;
    wire new_AGEMA_signal_14578 ;
    wire new_AGEMA_signal_14579 ;
    wire new_AGEMA_signal_14580 ;
    wire new_AGEMA_signal_14581 ;
    wire new_AGEMA_signal_14582 ;
    wire new_AGEMA_signal_14583 ;
    wire new_AGEMA_signal_14584 ;
    wire new_AGEMA_signal_14585 ;
    wire new_AGEMA_signal_14586 ;
    wire new_AGEMA_signal_14587 ;
    wire new_AGEMA_signal_14588 ;
    wire new_AGEMA_signal_14589 ;
    wire new_AGEMA_signal_14590 ;
    wire new_AGEMA_signal_14591 ;
    wire new_AGEMA_signal_14592 ;
    wire new_AGEMA_signal_14593 ;
    wire new_AGEMA_signal_14594 ;
    wire new_AGEMA_signal_14595 ;
    wire new_AGEMA_signal_14596 ;
    wire new_AGEMA_signal_14597 ;
    wire new_AGEMA_signal_14598 ;
    wire new_AGEMA_signal_14599 ;
    wire new_AGEMA_signal_14600 ;
    wire new_AGEMA_signal_14601 ;
    wire new_AGEMA_signal_14602 ;
    wire new_AGEMA_signal_14603 ;
    wire new_AGEMA_signal_14604 ;
    wire new_AGEMA_signal_14605 ;
    wire new_AGEMA_signal_14606 ;
    wire new_AGEMA_signal_14607 ;
    wire new_AGEMA_signal_14608 ;
    wire new_AGEMA_signal_14609 ;
    wire new_AGEMA_signal_14610 ;
    wire new_AGEMA_signal_14611 ;
    wire new_AGEMA_signal_14612 ;
    wire new_AGEMA_signal_14613 ;
    wire new_AGEMA_signal_14614 ;
    wire new_AGEMA_signal_14615 ;
    wire new_AGEMA_signal_14616 ;
    wire new_AGEMA_signal_14617 ;
    wire new_AGEMA_signal_14618 ;
    wire new_AGEMA_signal_14619 ;
    wire new_AGEMA_signal_14620 ;
    wire new_AGEMA_signal_14621 ;
    wire new_AGEMA_signal_14622 ;
    wire new_AGEMA_signal_14623 ;
    wire new_AGEMA_signal_14624 ;
    wire new_AGEMA_signal_14625 ;
    wire new_AGEMA_signal_14626 ;
    wire new_AGEMA_signal_14627 ;
    wire new_AGEMA_signal_14628 ;
    wire new_AGEMA_signal_14629 ;
    wire new_AGEMA_signal_14630 ;
    wire new_AGEMA_signal_14631 ;
    wire new_AGEMA_signal_14632 ;
    wire new_AGEMA_signal_14633 ;
    wire new_AGEMA_signal_14634 ;
    wire new_AGEMA_signal_14635 ;
    wire new_AGEMA_signal_14636 ;
    wire new_AGEMA_signal_14637 ;
    wire new_AGEMA_signal_14638 ;
    wire new_AGEMA_signal_14639 ;
    wire new_AGEMA_signal_14640 ;
    wire new_AGEMA_signal_14641 ;
    wire new_AGEMA_signal_14642 ;
    wire new_AGEMA_signal_14643 ;
    wire new_AGEMA_signal_14644 ;
    wire new_AGEMA_signal_14645 ;
    wire new_AGEMA_signal_14646 ;
    wire new_AGEMA_signal_14647 ;
    wire new_AGEMA_signal_14648 ;
    wire new_AGEMA_signal_14649 ;
    wire new_AGEMA_signal_14650 ;
    wire new_AGEMA_signal_14651 ;
    wire new_AGEMA_signal_14652 ;
    wire new_AGEMA_signal_14653 ;
    wire new_AGEMA_signal_14654 ;
    wire new_AGEMA_signal_14655 ;
    wire new_AGEMA_signal_14656 ;
    wire new_AGEMA_signal_14657 ;
    wire new_AGEMA_signal_14658 ;
    wire new_AGEMA_signal_14659 ;
    wire new_AGEMA_signal_14660 ;
    wire new_AGEMA_signal_14661 ;
    wire new_AGEMA_signal_14662 ;
    wire new_AGEMA_signal_14663 ;
    wire new_AGEMA_signal_14664 ;
    wire new_AGEMA_signal_14665 ;
    wire new_AGEMA_signal_14666 ;
    wire new_AGEMA_signal_14667 ;
    wire new_AGEMA_signal_14668 ;
    wire new_AGEMA_signal_14669 ;
    wire new_AGEMA_signal_14670 ;
    wire new_AGEMA_signal_14671 ;
    wire new_AGEMA_signal_14672 ;
    wire new_AGEMA_signal_14673 ;
    wire new_AGEMA_signal_14674 ;
    wire new_AGEMA_signal_14675 ;
    wire new_AGEMA_signal_14676 ;
    wire new_AGEMA_signal_14677 ;
    wire new_AGEMA_signal_14678 ;
    wire new_AGEMA_signal_14679 ;
    wire new_AGEMA_signal_14680 ;
    wire new_AGEMA_signal_14681 ;
    wire new_AGEMA_signal_14682 ;
    wire new_AGEMA_signal_14683 ;
    wire new_AGEMA_signal_14684 ;
    wire new_AGEMA_signal_14685 ;
    wire new_AGEMA_signal_14686 ;
    wire new_AGEMA_signal_14687 ;
    wire new_AGEMA_signal_14688 ;
    wire new_AGEMA_signal_14689 ;
    wire new_AGEMA_signal_14690 ;
    wire new_AGEMA_signal_14691 ;
    wire new_AGEMA_signal_14692 ;
    wire new_AGEMA_signal_14693 ;
    wire new_AGEMA_signal_14694 ;
    wire new_AGEMA_signal_14695 ;
    wire new_AGEMA_signal_14696 ;
    wire new_AGEMA_signal_14697 ;
    wire new_AGEMA_signal_14698 ;
    wire new_AGEMA_signal_14699 ;
    wire new_AGEMA_signal_14700 ;
    wire new_AGEMA_signal_14701 ;
    wire new_AGEMA_signal_14702 ;
    wire new_AGEMA_signal_14703 ;
    wire new_AGEMA_signal_14704 ;
    wire new_AGEMA_signal_14705 ;
    wire new_AGEMA_signal_14706 ;
    wire new_AGEMA_signal_14707 ;
    wire new_AGEMA_signal_14708 ;
    wire new_AGEMA_signal_14709 ;
    wire new_AGEMA_signal_14710 ;
    wire new_AGEMA_signal_14711 ;
    wire new_AGEMA_signal_14712 ;
    wire new_AGEMA_signal_14713 ;
    wire new_AGEMA_signal_14714 ;
    wire new_AGEMA_signal_14715 ;
    wire new_AGEMA_signal_14716 ;
    wire new_AGEMA_signal_14717 ;
    wire new_AGEMA_signal_14718 ;
    wire new_AGEMA_signal_14719 ;
    wire new_AGEMA_signal_14720 ;
    wire new_AGEMA_signal_14721 ;
    wire new_AGEMA_signal_14722 ;
    wire new_AGEMA_signal_14723 ;
    wire new_AGEMA_signal_14724 ;
    wire new_AGEMA_signal_14725 ;
    wire new_AGEMA_signal_14726 ;
    wire new_AGEMA_signal_14727 ;
    wire new_AGEMA_signal_14728 ;
    wire new_AGEMA_signal_14729 ;
    wire new_AGEMA_signal_14730 ;
    wire new_AGEMA_signal_14731 ;
    wire new_AGEMA_signal_14732 ;
    wire new_AGEMA_signal_14733 ;
    wire new_AGEMA_signal_14734 ;
    wire new_AGEMA_signal_14735 ;
    wire new_AGEMA_signal_14736 ;
    wire new_AGEMA_signal_14737 ;
    wire new_AGEMA_signal_14738 ;
    wire new_AGEMA_signal_14739 ;
    wire new_AGEMA_signal_14740 ;
    wire new_AGEMA_signal_14741 ;
    wire new_AGEMA_signal_14742 ;
    wire new_AGEMA_signal_14743 ;
    wire new_AGEMA_signal_14744 ;
    wire new_AGEMA_signal_14745 ;
    wire new_AGEMA_signal_14746 ;
    wire new_AGEMA_signal_14747 ;
    wire new_AGEMA_signal_14748 ;
    wire new_AGEMA_signal_14749 ;
    wire new_AGEMA_signal_14750 ;
    wire new_AGEMA_signal_14751 ;
    wire new_AGEMA_signal_14752 ;
    wire new_AGEMA_signal_14753 ;
    wire new_AGEMA_signal_14754 ;
    wire new_AGEMA_signal_14755 ;
    wire new_AGEMA_signal_14756 ;
    wire new_AGEMA_signal_14757 ;
    wire new_AGEMA_signal_14758 ;
    wire new_AGEMA_signal_14759 ;
    wire new_AGEMA_signal_14760 ;
    wire new_AGEMA_signal_14761 ;
    wire new_AGEMA_signal_14762 ;
    wire new_AGEMA_signal_14763 ;
    wire new_AGEMA_signal_14764 ;
    wire new_AGEMA_signal_14765 ;
    wire new_AGEMA_signal_14766 ;
    wire new_AGEMA_signal_14767 ;
    wire new_AGEMA_signal_14768 ;
    wire new_AGEMA_signal_14769 ;
    wire new_AGEMA_signal_14770 ;
    wire new_AGEMA_signal_14771 ;
    wire new_AGEMA_signal_14772 ;
    wire new_AGEMA_signal_14773 ;
    wire new_AGEMA_signal_14774 ;
    wire new_AGEMA_signal_14775 ;
    wire new_AGEMA_signal_14776 ;
    wire new_AGEMA_signal_14777 ;
    wire new_AGEMA_signal_14778 ;
    wire new_AGEMA_signal_14779 ;
    wire new_AGEMA_signal_14780 ;
    wire new_AGEMA_signal_14781 ;
    wire new_AGEMA_signal_14782 ;
    wire new_AGEMA_signal_14783 ;
    wire new_AGEMA_signal_14784 ;
    wire new_AGEMA_signal_14785 ;
    wire new_AGEMA_signal_14786 ;
    wire new_AGEMA_signal_14787 ;
    wire new_AGEMA_signal_14788 ;
    wire new_AGEMA_signal_14789 ;
    wire new_AGEMA_signal_14790 ;
    wire new_AGEMA_signal_14791 ;
    wire new_AGEMA_signal_14792 ;
    wire new_AGEMA_signal_14793 ;
    wire new_AGEMA_signal_14794 ;
    wire new_AGEMA_signal_14795 ;
    wire new_AGEMA_signal_14796 ;
    wire new_AGEMA_signal_14797 ;
    wire new_AGEMA_signal_14798 ;
    wire new_AGEMA_signal_14799 ;
    wire new_AGEMA_signal_14800 ;
    wire new_AGEMA_signal_14801 ;
    wire new_AGEMA_signal_14802 ;
    wire new_AGEMA_signal_14803 ;
    wire new_AGEMA_signal_14804 ;
    wire new_AGEMA_signal_14805 ;
    wire new_AGEMA_signal_14806 ;
    wire new_AGEMA_signal_14807 ;
    wire new_AGEMA_signal_14808 ;
    wire new_AGEMA_signal_14809 ;
    wire new_AGEMA_signal_14810 ;
    wire new_AGEMA_signal_14811 ;
    wire new_AGEMA_signal_14812 ;
    wire new_AGEMA_signal_14813 ;
    wire new_AGEMA_signal_14814 ;
    wire new_AGEMA_signal_14815 ;
    wire new_AGEMA_signal_14816 ;
    wire new_AGEMA_signal_14817 ;
    wire new_AGEMA_signal_14818 ;
    wire new_AGEMA_signal_14819 ;
    wire new_AGEMA_signal_14820 ;
    wire new_AGEMA_signal_14821 ;
    wire new_AGEMA_signal_14822 ;
    wire new_AGEMA_signal_14823 ;
    wire new_AGEMA_signal_14824 ;
    wire new_AGEMA_signal_14825 ;
    wire new_AGEMA_signal_14826 ;
    wire new_AGEMA_signal_14827 ;
    wire new_AGEMA_signal_14828 ;
    wire new_AGEMA_signal_14829 ;
    wire new_AGEMA_signal_14830 ;
    wire new_AGEMA_signal_14831 ;
    wire new_AGEMA_signal_14832 ;
    wire new_AGEMA_signal_14833 ;
    wire new_AGEMA_signal_14834 ;
    wire new_AGEMA_signal_14835 ;
    wire new_AGEMA_signal_14836 ;
    wire new_AGEMA_signal_14837 ;
    wire new_AGEMA_signal_14838 ;
    wire new_AGEMA_signal_14839 ;
    wire new_AGEMA_signal_14840 ;
    wire new_AGEMA_signal_14841 ;
    wire new_AGEMA_signal_14842 ;
    wire new_AGEMA_signal_14843 ;
    wire new_AGEMA_signal_14844 ;
    wire new_AGEMA_signal_14845 ;
    wire new_AGEMA_signal_14846 ;
    wire new_AGEMA_signal_14847 ;
    wire new_AGEMA_signal_14848 ;
    wire new_AGEMA_signal_14849 ;
    wire new_AGEMA_signal_14850 ;
    wire new_AGEMA_signal_14851 ;
    wire new_AGEMA_signal_14852 ;
    wire new_AGEMA_signal_14853 ;
    wire new_AGEMA_signal_14854 ;
    wire new_AGEMA_signal_14855 ;
    wire new_AGEMA_signal_14856 ;
    wire new_AGEMA_signal_14857 ;
    wire new_AGEMA_signal_14858 ;
    wire new_AGEMA_signal_14859 ;
    wire new_AGEMA_signal_14860 ;
    wire new_AGEMA_signal_14861 ;
    wire new_AGEMA_signal_14862 ;
    wire new_AGEMA_signal_14863 ;
    wire new_AGEMA_signal_14864 ;
    wire new_AGEMA_signal_14865 ;
    wire new_AGEMA_signal_14866 ;
    wire new_AGEMA_signal_14867 ;
    wire new_AGEMA_signal_14868 ;
    wire new_AGEMA_signal_14869 ;
    wire new_AGEMA_signal_14870 ;
    wire new_AGEMA_signal_14871 ;
    wire new_AGEMA_signal_14872 ;
    wire new_AGEMA_signal_14873 ;
    wire new_AGEMA_signal_14874 ;
    wire new_AGEMA_signal_14875 ;
    wire new_AGEMA_signal_14876 ;
    wire new_AGEMA_signal_14877 ;
    wire new_AGEMA_signal_14878 ;
    wire new_AGEMA_signal_14879 ;
    wire new_AGEMA_signal_14880 ;
    wire new_AGEMA_signal_14881 ;
    wire new_AGEMA_signal_14882 ;
    wire new_AGEMA_signal_14883 ;
    wire new_AGEMA_signal_14884 ;
    wire new_AGEMA_signal_14885 ;
    wire new_AGEMA_signal_14886 ;
    wire new_AGEMA_signal_14887 ;
    wire new_AGEMA_signal_14888 ;
    wire new_AGEMA_signal_14889 ;
    wire new_AGEMA_signal_14890 ;
    wire new_AGEMA_signal_14891 ;
    wire new_AGEMA_signal_14892 ;
    wire new_AGEMA_signal_14893 ;
    wire new_AGEMA_signal_14894 ;
    wire new_AGEMA_signal_14895 ;
    wire new_AGEMA_signal_14896 ;
    wire new_AGEMA_signal_14897 ;
    wire new_AGEMA_signal_14898 ;
    wire new_AGEMA_signal_14899 ;
    wire new_AGEMA_signal_14900 ;
    wire new_AGEMA_signal_14901 ;
    wire new_AGEMA_signal_14902 ;
    wire new_AGEMA_signal_14903 ;
    wire new_AGEMA_signal_14904 ;
    wire new_AGEMA_signal_14905 ;
    wire new_AGEMA_signal_14906 ;
    wire new_AGEMA_signal_14907 ;
    wire new_AGEMA_signal_14908 ;
    wire new_AGEMA_signal_14909 ;
    wire new_AGEMA_signal_14910 ;
    wire new_AGEMA_signal_14911 ;
    wire new_AGEMA_signal_14912 ;
    wire new_AGEMA_signal_14913 ;
    wire new_AGEMA_signal_14914 ;
    wire new_AGEMA_signal_14915 ;
    wire new_AGEMA_signal_14916 ;
    wire new_AGEMA_signal_14917 ;
    wire new_AGEMA_signal_14918 ;
    wire new_AGEMA_signal_14919 ;
    wire new_AGEMA_signal_14920 ;
    wire new_AGEMA_signal_14921 ;
    wire new_AGEMA_signal_14922 ;
    wire new_AGEMA_signal_14923 ;
    wire new_AGEMA_signal_14924 ;
    wire new_AGEMA_signal_14925 ;
    wire new_AGEMA_signal_14926 ;
    wire new_AGEMA_signal_14927 ;
    wire new_AGEMA_signal_14928 ;
    wire new_AGEMA_signal_14929 ;
    wire new_AGEMA_signal_14930 ;
    wire new_AGEMA_signal_14931 ;
    wire new_AGEMA_signal_14932 ;
    wire new_AGEMA_signal_14933 ;
    wire new_AGEMA_signal_14934 ;
    wire new_AGEMA_signal_14935 ;
    wire new_AGEMA_signal_14936 ;
    wire new_AGEMA_signal_14937 ;
    wire new_AGEMA_signal_14938 ;
    wire new_AGEMA_signal_14939 ;
    wire new_AGEMA_signal_14940 ;
    wire new_AGEMA_signal_14941 ;
    wire new_AGEMA_signal_14942 ;
    wire new_AGEMA_signal_14943 ;
    wire new_AGEMA_signal_14944 ;
    wire new_AGEMA_signal_14945 ;
    wire new_AGEMA_signal_14946 ;
    wire new_AGEMA_signal_14947 ;
    wire new_AGEMA_signal_14948 ;
    wire new_AGEMA_signal_14949 ;
    wire new_AGEMA_signal_14950 ;
    wire new_AGEMA_signal_14951 ;
    wire new_AGEMA_signal_14952 ;
    wire new_AGEMA_signal_14953 ;
    wire new_AGEMA_signal_14954 ;
    wire new_AGEMA_signal_14955 ;
    wire new_AGEMA_signal_14956 ;
    wire new_AGEMA_signal_14957 ;
    wire new_AGEMA_signal_14958 ;
    wire new_AGEMA_signal_14959 ;
    wire new_AGEMA_signal_14960 ;
    wire new_AGEMA_signal_14961 ;
    wire new_AGEMA_signal_14962 ;
    wire new_AGEMA_signal_14963 ;
    wire new_AGEMA_signal_14964 ;
    wire new_AGEMA_signal_14965 ;
    wire new_AGEMA_signal_14966 ;
    wire new_AGEMA_signal_14967 ;
    wire new_AGEMA_signal_14968 ;
    wire new_AGEMA_signal_14969 ;
    wire new_AGEMA_signal_14970 ;
    wire new_AGEMA_signal_14971 ;
    wire new_AGEMA_signal_14972 ;
    wire new_AGEMA_signal_14973 ;
    wire new_AGEMA_signal_14974 ;
    wire new_AGEMA_signal_14975 ;
    wire new_AGEMA_signal_14976 ;
    wire new_AGEMA_signal_14977 ;
    wire new_AGEMA_signal_14978 ;
    wire new_AGEMA_signal_14979 ;
    wire new_AGEMA_signal_14980 ;
    wire new_AGEMA_signal_14981 ;
    wire new_AGEMA_signal_14982 ;
    wire new_AGEMA_signal_14983 ;
    wire new_AGEMA_signal_14984 ;
    wire new_AGEMA_signal_14985 ;
    wire new_AGEMA_signal_14986 ;
    wire new_AGEMA_signal_14987 ;
    wire new_AGEMA_signal_14988 ;
    wire new_AGEMA_signal_14989 ;
    wire new_AGEMA_signal_14990 ;
    wire new_AGEMA_signal_14991 ;
    wire new_AGEMA_signal_14992 ;
    wire new_AGEMA_signal_14993 ;
    wire new_AGEMA_signal_14994 ;
    wire new_AGEMA_signal_14995 ;
    wire new_AGEMA_signal_14996 ;
    wire new_AGEMA_signal_14997 ;
    wire new_AGEMA_signal_14998 ;
    wire new_AGEMA_signal_14999 ;
    wire new_AGEMA_signal_15000 ;
    wire new_AGEMA_signal_15001 ;
    wire new_AGEMA_signal_15002 ;
    wire new_AGEMA_signal_15003 ;
    wire new_AGEMA_signal_15004 ;
    wire new_AGEMA_signal_15005 ;
    wire new_AGEMA_signal_15006 ;
    wire new_AGEMA_signal_15007 ;
    wire new_AGEMA_signal_15008 ;
    wire new_AGEMA_signal_15009 ;
    wire new_AGEMA_signal_15010 ;
    wire new_AGEMA_signal_15011 ;
    wire new_AGEMA_signal_15012 ;
    wire new_AGEMA_signal_15013 ;
    wire new_AGEMA_signal_15014 ;
    wire new_AGEMA_signal_15015 ;
    wire new_AGEMA_signal_15016 ;
    wire new_AGEMA_signal_15017 ;
    wire new_AGEMA_signal_15018 ;
    wire new_AGEMA_signal_15019 ;
    wire new_AGEMA_signal_15020 ;
    wire new_AGEMA_signal_15021 ;
    wire new_AGEMA_signal_15022 ;
    wire new_AGEMA_signal_15023 ;
    wire new_AGEMA_signal_15024 ;
    wire new_AGEMA_signal_15025 ;
    wire new_AGEMA_signal_15026 ;
    wire new_AGEMA_signal_15027 ;
    wire new_AGEMA_signal_15028 ;
    wire new_AGEMA_signal_15029 ;
    wire new_AGEMA_signal_15030 ;
    wire new_AGEMA_signal_15031 ;
    wire new_AGEMA_signal_15032 ;
    wire new_AGEMA_signal_15033 ;
    wire new_AGEMA_signal_15034 ;
    wire new_AGEMA_signal_15035 ;
    wire new_AGEMA_signal_15036 ;
    wire new_AGEMA_signal_15037 ;
    wire new_AGEMA_signal_15038 ;
    wire new_AGEMA_signal_15039 ;
    wire new_AGEMA_signal_15040 ;
    wire new_AGEMA_signal_15041 ;
    wire new_AGEMA_signal_15042 ;
    wire new_AGEMA_signal_15043 ;
    wire new_AGEMA_signal_15044 ;
    wire new_AGEMA_signal_15045 ;
    wire new_AGEMA_signal_15046 ;
    wire new_AGEMA_signal_15047 ;
    wire new_AGEMA_signal_15048 ;
    wire new_AGEMA_signal_15049 ;
    wire new_AGEMA_signal_15050 ;
    wire new_AGEMA_signal_15051 ;
    wire new_AGEMA_signal_15052 ;
    wire new_AGEMA_signal_15053 ;
    wire new_AGEMA_signal_15054 ;
    wire new_AGEMA_signal_15055 ;
    wire new_AGEMA_signal_15056 ;
    wire new_AGEMA_signal_15057 ;
    wire new_AGEMA_signal_15058 ;
    wire new_AGEMA_signal_15059 ;
    wire new_AGEMA_signal_15060 ;
    wire new_AGEMA_signal_15061 ;
    wire new_AGEMA_signal_15062 ;
    wire new_AGEMA_signal_15063 ;
    wire new_AGEMA_signal_15064 ;
    wire new_AGEMA_signal_15065 ;
    wire new_AGEMA_signal_15066 ;
    wire new_AGEMA_signal_15067 ;
    wire new_AGEMA_signal_15068 ;
    wire new_AGEMA_signal_15069 ;
    wire new_AGEMA_signal_15070 ;
    wire new_AGEMA_signal_15071 ;
    wire new_AGEMA_signal_15072 ;
    wire new_AGEMA_signal_15073 ;
    wire new_AGEMA_signal_15074 ;
    wire new_AGEMA_signal_15075 ;
    wire new_AGEMA_signal_15076 ;
    wire new_AGEMA_signal_15077 ;
    wire new_AGEMA_signal_15078 ;
    wire new_AGEMA_signal_15079 ;
    wire new_AGEMA_signal_15080 ;
    wire new_AGEMA_signal_15081 ;
    wire new_AGEMA_signal_15082 ;
    wire new_AGEMA_signal_15083 ;
    wire new_AGEMA_signal_15084 ;
    wire new_AGEMA_signal_15085 ;
    wire new_AGEMA_signal_15086 ;
    wire new_AGEMA_signal_15087 ;
    wire new_AGEMA_signal_15088 ;
    wire new_AGEMA_signal_15089 ;
    wire new_AGEMA_signal_15090 ;
    wire new_AGEMA_signal_15091 ;
    wire new_AGEMA_signal_15092 ;
    wire new_AGEMA_signal_15093 ;
    wire new_AGEMA_signal_15094 ;
    wire new_AGEMA_signal_15095 ;
    wire new_AGEMA_signal_15096 ;
    wire new_AGEMA_signal_15097 ;
    wire new_AGEMA_signal_15098 ;
    wire new_AGEMA_signal_15099 ;
    wire new_AGEMA_signal_15100 ;
    wire new_AGEMA_signal_15101 ;
    wire new_AGEMA_signal_15102 ;
    wire new_AGEMA_signal_15103 ;
    wire new_AGEMA_signal_15104 ;
    wire new_AGEMA_signal_15105 ;
    wire new_AGEMA_signal_15106 ;
    wire new_AGEMA_signal_15107 ;
    wire new_AGEMA_signal_15108 ;
    wire new_AGEMA_signal_15109 ;
    wire new_AGEMA_signal_15110 ;
    wire new_AGEMA_signal_15111 ;
    wire new_AGEMA_signal_15112 ;
    wire new_AGEMA_signal_15113 ;
    wire new_AGEMA_signal_15114 ;
    wire new_AGEMA_signal_15115 ;
    wire new_AGEMA_signal_15116 ;
    wire new_AGEMA_signal_15117 ;
    wire new_AGEMA_signal_15118 ;
    wire new_AGEMA_signal_15119 ;
    wire new_AGEMA_signal_15120 ;
    wire new_AGEMA_signal_15121 ;
    wire new_AGEMA_signal_15122 ;
    wire new_AGEMA_signal_15123 ;
    wire new_AGEMA_signal_15124 ;
    wire new_AGEMA_signal_15125 ;
    wire new_AGEMA_signal_15126 ;
    wire new_AGEMA_signal_15127 ;
    wire new_AGEMA_signal_15128 ;
    wire new_AGEMA_signal_15129 ;
    wire new_AGEMA_signal_15130 ;
    wire new_AGEMA_signal_15131 ;
    wire new_AGEMA_signal_15132 ;
    wire new_AGEMA_signal_15133 ;
    wire new_AGEMA_signal_15134 ;
    wire new_AGEMA_signal_15135 ;
    wire new_AGEMA_signal_15136 ;
    wire new_AGEMA_signal_15137 ;
    wire new_AGEMA_signal_15138 ;
    wire new_AGEMA_signal_15139 ;
    wire new_AGEMA_signal_15140 ;
    wire new_AGEMA_signal_15141 ;
    wire new_AGEMA_signal_15142 ;
    wire new_AGEMA_signal_15143 ;
    wire new_AGEMA_signal_15144 ;
    wire new_AGEMA_signal_15145 ;
    wire new_AGEMA_signal_15146 ;
    wire new_AGEMA_signal_15147 ;
    wire new_AGEMA_signal_15148 ;
    wire new_AGEMA_signal_15149 ;
    wire new_AGEMA_signal_15150 ;
    wire new_AGEMA_signal_15151 ;
    wire new_AGEMA_signal_15152 ;
    wire new_AGEMA_signal_15153 ;
    wire new_AGEMA_signal_15154 ;
    wire new_AGEMA_signal_15155 ;
    wire new_AGEMA_signal_15156 ;
    wire new_AGEMA_signal_15157 ;
    wire new_AGEMA_signal_15158 ;
    wire new_AGEMA_signal_15159 ;
    wire new_AGEMA_signal_15160 ;
    wire new_AGEMA_signal_15161 ;
    wire new_AGEMA_signal_15162 ;
    wire new_AGEMA_signal_15163 ;
    wire new_AGEMA_signal_15164 ;
    wire new_AGEMA_signal_15165 ;
    wire new_AGEMA_signal_15166 ;
    wire new_AGEMA_signal_15167 ;
    wire new_AGEMA_signal_15168 ;
    wire new_AGEMA_signal_15169 ;
    wire new_AGEMA_signal_15170 ;
    wire new_AGEMA_signal_15171 ;
    wire new_AGEMA_signal_15172 ;
    wire new_AGEMA_signal_15173 ;
    wire new_AGEMA_signal_15174 ;
    wire new_AGEMA_signal_15175 ;
    wire new_AGEMA_signal_15176 ;
    wire new_AGEMA_signal_15177 ;
    wire new_AGEMA_signal_15178 ;
    wire new_AGEMA_signal_15179 ;
    wire new_AGEMA_signal_15180 ;
    wire new_AGEMA_signal_15181 ;
    wire new_AGEMA_signal_15182 ;
    wire new_AGEMA_signal_15183 ;
    wire new_AGEMA_signal_15184 ;
    wire new_AGEMA_signal_15185 ;
    wire new_AGEMA_signal_15186 ;
    wire new_AGEMA_signal_15187 ;
    wire new_AGEMA_signal_15188 ;
    wire new_AGEMA_signal_15189 ;
    wire new_AGEMA_signal_15190 ;
    wire new_AGEMA_signal_15191 ;
    wire new_AGEMA_signal_15192 ;
    wire new_AGEMA_signal_15193 ;
    wire new_AGEMA_signal_15194 ;
    wire new_AGEMA_signal_15195 ;
    wire new_AGEMA_signal_15196 ;
    wire new_AGEMA_signal_15197 ;
    wire new_AGEMA_signal_15198 ;
    wire new_AGEMA_signal_15199 ;
    wire new_AGEMA_signal_15200 ;
    wire new_AGEMA_signal_15201 ;
    wire new_AGEMA_signal_15202 ;
    wire new_AGEMA_signal_15203 ;
    wire new_AGEMA_signal_15204 ;
    wire new_AGEMA_signal_15205 ;
    wire new_AGEMA_signal_15206 ;
    wire new_AGEMA_signal_15207 ;
    wire new_AGEMA_signal_15208 ;
    wire new_AGEMA_signal_15209 ;
    wire new_AGEMA_signal_15210 ;
    wire new_AGEMA_signal_15211 ;
    wire new_AGEMA_signal_15212 ;
    wire new_AGEMA_signal_15213 ;
    wire new_AGEMA_signal_15214 ;
    wire new_AGEMA_signal_15215 ;
    wire new_AGEMA_signal_15216 ;
    wire new_AGEMA_signal_15217 ;
    wire new_AGEMA_signal_15218 ;
    wire new_AGEMA_signal_15219 ;
    wire new_AGEMA_signal_15220 ;
    wire new_AGEMA_signal_15221 ;
    wire new_AGEMA_signal_15222 ;
    wire new_AGEMA_signal_15223 ;
    wire new_AGEMA_signal_15224 ;
    wire new_AGEMA_signal_15225 ;
    wire new_AGEMA_signal_15226 ;
    wire new_AGEMA_signal_15227 ;
    wire new_AGEMA_signal_15228 ;
    wire new_AGEMA_signal_15229 ;
    wire new_AGEMA_signal_15230 ;
    wire new_AGEMA_signal_15231 ;
    wire new_AGEMA_signal_15232 ;
    wire new_AGEMA_signal_15233 ;
    wire new_AGEMA_signal_15234 ;
    wire new_AGEMA_signal_15235 ;
    wire new_AGEMA_signal_15236 ;
    wire new_AGEMA_signal_15237 ;
    wire new_AGEMA_signal_15238 ;
    wire new_AGEMA_signal_15239 ;
    wire new_AGEMA_signal_15240 ;
    wire new_AGEMA_signal_15241 ;
    wire new_AGEMA_signal_15242 ;
    wire new_AGEMA_signal_15243 ;
    wire new_AGEMA_signal_15244 ;
    wire new_AGEMA_signal_15245 ;
    wire new_AGEMA_signal_15246 ;
    wire new_AGEMA_signal_15247 ;
    wire new_AGEMA_signal_15248 ;
    wire new_AGEMA_signal_15249 ;
    wire new_AGEMA_signal_15250 ;
    wire new_AGEMA_signal_15251 ;
    wire new_AGEMA_signal_15252 ;
    wire new_AGEMA_signal_15253 ;
    wire new_AGEMA_signal_15254 ;
    wire new_AGEMA_signal_15255 ;
    wire new_AGEMA_signal_15256 ;
    wire new_AGEMA_signal_15257 ;
    wire new_AGEMA_signal_15258 ;
    wire new_AGEMA_signal_15259 ;
    wire new_AGEMA_signal_15260 ;
    wire new_AGEMA_signal_15261 ;
    wire new_AGEMA_signal_15262 ;
    wire new_AGEMA_signal_15263 ;
    wire new_AGEMA_signal_15264 ;
    wire new_AGEMA_signal_15265 ;
    wire new_AGEMA_signal_15266 ;
    wire new_AGEMA_signal_15267 ;
    wire new_AGEMA_signal_15268 ;
    wire new_AGEMA_signal_15269 ;
    wire new_AGEMA_signal_15270 ;
    wire new_AGEMA_signal_15271 ;
    wire new_AGEMA_signal_15272 ;
    wire new_AGEMA_signal_15273 ;
    wire new_AGEMA_signal_15274 ;
    wire new_AGEMA_signal_15275 ;
    wire new_AGEMA_signal_15276 ;
    wire new_AGEMA_signal_15277 ;
    wire new_AGEMA_signal_15278 ;
    wire new_AGEMA_signal_15279 ;
    wire new_AGEMA_signal_15280 ;
    wire new_AGEMA_signal_15281 ;
    wire new_AGEMA_signal_15282 ;
    wire new_AGEMA_signal_15283 ;
    wire new_AGEMA_signal_15284 ;
    wire new_AGEMA_signal_15285 ;
    wire new_AGEMA_signal_15286 ;
    wire new_AGEMA_signal_15287 ;
    wire new_AGEMA_signal_15288 ;
    wire new_AGEMA_signal_15289 ;
    wire new_AGEMA_signal_15290 ;
    wire new_AGEMA_signal_15291 ;
    wire new_AGEMA_signal_15292 ;
    wire new_AGEMA_signal_15293 ;
    wire new_AGEMA_signal_15294 ;
    wire new_AGEMA_signal_15295 ;
    wire new_AGEMA_signal_15296 ;
    wire new_AGEMA_signal_15297 ;
    wire new_AGEMA_signal_15298 ;
    wire new_AGEMA_signal_15299 ;
    wire new_AGEMA_signal_15300 ;
    wire new_AGEMA_signal_15301 ;
    wire new_AGEMA_signal_15302 ;
    wire new_AGEMA_signal_15303 ;
    wire new_AGEMA_signal_15304 ;
    wire new_AGEMA_signal_15305 ;
    wire new_AGEMA_signal_15306 ;
    wire new_AGEMA_signal_15307 ;
    wire new_AGEMA_signal_15308 ;
    wire new_AGEMA_signal_15309 ;
    wire new_AGEMA_signal_15310 ;
    wire new_AGEMA_signal_15311 ;
    wire new_AGEMA_signal_15312 ;
    wire new_AGEMA_signal_15313 ;
    wire new_AGEMA_signal_15314 ;
    wire new_AGEMA_signal_15315 ;
    wire new_AGEMA_signal_15316 ;
    wire new_AGEMA_signal_15317 ;
    wire new_AGEMA_signal_15318 ;
    wire new_AGEMA_signal_15319 ;
    wire new_AGEMA_signal_15320 ;
    wire new_AGEMA_signal_15321 ;
    wire new_AGEMA_signal_15322 ;
    wire new_AGEMA_signal_15323 ;
    wire new_AGEMA_signal_15324 ;
    wire new_AGEMA_signal_15325 ;
    wire new_AGEMA_signal_15326 ;
    wire new_AGEMA_signal_15327 ;
    wire new_AGEMA_signal_15328 ;
    wire new_AGEMA_signal_15329 ;
    wire new_AGEMA_signal_15330 ;
    wire new_AGEMA_signal_15331 ;
    wire new_AGEMA_signal_15332 ;
    wire new_AGEMA_signal_15333 ;
    wire new_AGEMA_signal_15334 ;
    wire new_AGEMA_signal_15335 ;
    wire new_AGEMA_signal_15336 ;
    wire new_AGEMA_signal_15337 ;
    wire new_AGEMA_signal_15338 ;
    wire new_AGEMA_signal_15339 ;
    wire new_AGEMA_signal_15340 ;
    wire new_AGEMA_signal_15341 ;
    wire new_AGEMA_signal_15342 ;
    wire new_AGEMA_signal_15343 ;
    wire new_AGEMA_signal_15344 ;
    wire new_AGEMA_signal_15345 ;
    wire new_AGEMA_signal_15346 ;
    wire new_AGEMA_signal_15347 ;
    wire new_AGEMA_signal_15348 ;
    wire new_AGEMA_signal_15349 ;
    wire new_AGEMA_signal_15350 ;
    wire new_AGEMA_signal_15351 ;
    wire new_AGEMA_signal_15352 ;
    wire new_AGEMA_signal_15353 ;
    wire new_AGEMA_signal_15354 ;
    wire new_AGEMA_signal_15355 ;
    wire new_AGEMA_signal_15356 ;
    wire new_AGEMA_signal_15357 ;
    wire new_AGEMA_signal_15358 ;
    wire new_AGEMA_signal_15359 ;
    wire new_AGEMA_signal_15360 ;
    wire new_AGEMA_signal_15361 ;
    wire new_AGEMA_signal_15362 ;
    wire new_AGEMA_signal_15363 ;
    wire new_AGEMA_signal_15364 ;
    wire new_AGEMA_signal_15365 ;
    wire new_AGEMA_signal_15366 ;
    wire new_AGEMA_signal_15367 ;
    wire new_AGEMA_signal_15368 ;
    wire new_AGEMA_signal_15369 ;
    wire new_AGEMA_signal_15370 ;
    wire new_AGEMA_signal_15371 ;
    wire new_AGEMA_signal_15372 ;
    wire new_AGEMA_signal_15373 ;
    wire new_AGEMA_signal_15374 ;
    wire new_AGEMA_signal_15375 ;
    wire new_AGEMA_signal_15376 ;
    wire new_AGEMA_signal_15377 ;
    wire new_AGEMA_signal_15378 ;
    wire new_AGEMA_signal_15379 ;
    wire new_AGEMA_signal_15380 ;
    wire new_AGEMA_signal_15381 ;
    wire new_AGEMA_signal_15382 ;
    wire new_AGEMA_signal_15383 ;
    wire new_AGEMA_signal_15384 ;
    wire new_AGEMA_signal_15385 ;
    wire new_AGEMA_signal_15386 ;
    wire new_AGEMA_signal_15387 ;
    wire new_AGEMA_signal_15388 ;
    wire new_AGEMA_signal_15389 ;
    wire new_AGEMA_signal_15390 ;
    wire new_AGEMA_signal_15391 ;
    wire new_AGEMA_signal_15392 ;
    wire new_AGEMA_signal_15393 ;
    wire new_AGEMA_signal_15394 ;
    wire new_AGEMA_signal_15395 ;
    wire new_AGEMA_signal_15396 ;
    wire new_AGEMA_signal_15397 ;
    wire new_AGEMA_signal_15398 ;
    wire new_AGEMA_signal_15399 ;
    wire new_AGEMA_signal_15400 ;
    wire new_AGEMA_signal_15401 ;
    wire new_AGEMA_signal_15402 ;
    wire new_AGEMA_signal_15403 ;
    wire new_AGEMA_signal_15404 ;
    wire new_AGEMA_signal_15405 ;
    wire new_AGEMA_signal_15406 ;
    wire new_AGEMA_signal_15407 ;
    wire new_AGEMA_signal_15408 ;
    wire new_AGEMA_signal_15409 ;
    wire new_AGEMA_signal_15410 ;
    wire new_AGEMA_signal_15411 ;
    wire new_AGEMA_signal_15412 ;
    wire new_AGEMA_signal_15413 ;
    wire new_AGEMA_signal_15414 ;
    wire new_AGEMA_signal_15415 ;
    wire new_AGEMA_signal_15416 ;
    wire new_AGEMA_signal_15417 ;
    wire new_AGEMA_signal_15418 ;
    wire new_AGEMA_signal_15419 ;
    wire new_AGEMA_signal_15420 ;
    wire new_AGEMA_signal_15421 ;
    wire new_AGEMA_signal_15422 ;
    wire new_AGEMA_signal_15423 ;
    wire new_AGEMA_signal_15424 ;
    wire new_AGEMA_signal_15425 ;
    wire new_AGEMA_signal_15426 ;
    wire new_AGEMA_signal_15427 ;
    wire new_AGEMA_signal_15428 ;
    wire new_AGEMA_signal_15429 ;
    wire new_AGEMA_signal_15430 ;
    wire new_AGEMA_signal_15431 ;
    wire new_AGEMA_signal_15432 ;
    wire new_AGEMA_signal_15433 ;
    wire new_AGEMA_signal_15434 ;
    wire new_AGEMA_signal_15435 ;
    wire new_AGEMA_signal_15436 ;
    wire new_AGEMA_signal_15437 ;
    wire new_AGEMA_signal_15438 ;
    wire new_AGEMA_signal_15439 ;
    wire new_AGEMA_signal_15440 ;
    wire new_AGEMA_signal_15441 ;
    wire new_AGEMA_signal_15442 ;
    wire new_AGEMA_signal_15443 ;
    wire new_AGEMA_signal_15444 ;
    wire new_AGEMA_signal_15445 ;
    wire new_AGEMA_signal_15446 ;
    wire new_AGEMA_signal_15447 ;
    wire new_AGEMA_signal_15448 ;
    wire new_AGEMA_signal_15449 ;
    wire new_AGEMA_signal_15450 ;
    wire new_AGEMA_signal_15451 ;
    wire new_AGEMA_signal_15452 ;
    wire new_AGEMA_signal_15453 ;
    wire new_AGEMA_signal_15454 ;
    wire new_AGEMA_signal_15455 ;
    wire new_AGEMA_signal_15456 ;
    wire new_AGEMA_signal_15457 ;
    wire new_AGEMA_signal_15458 ;
    wire new_AGEMA_signal_15459 ;
    wire new_AGEMA_signal_15460 ;
    wire new_AGEMA_signal_15461 ;
    wire new_AGEMA_signal_15462 ;
    wire new_AGEMA_signal_15463 ;
    wire new_AGEMA_signal_15464 ;
    wire new_AGEMA_signal_15465 ;
    wire new_AGEMA_signal_15466 ;
    wire new_AGEMA_signal_15467 ;
    wire new_AGEMA_signal_15468 ;
    wire new_AGEMA_signal_15469 ;
    wire new_AGEMA_signal_15470 ;
    wire new_AGEMA_signal_15471 ;
    wire new_AGEMA_signal_15472 ;
    wire new_AGEMA_signal_15473 ;
    wire new_AGEMA_signal_15474 ;
    wire new_AGEMA_signal_15475 ;
    wire new_AGEMA_signal_15476 ;
    wire new_AGEMA_signal_15477 ;
    wire new_AGEMA_signal_15478 ;
    wire new_AGEMA_signal_15479 ;
    wire new_AGEMA_signal_15480 ;
    wire new_AGEMA_signal_15481 ;
    wire new_AGEMA_signal_15482 ;
    wire new_AGEMA_signal_15483 ;
    wire new_AGEMA_signal_15484 ;
    wire new_AGEMA_signal_15485 ;
    wire new_AGEMA_signal_15486 ;
    wire new_AGEMA_signal_15487 ;
    wire new_AGEMA_signal_15488 ;
    wire new_AGEMA_signal_15489 ;
    wire new_AGEMA_signal_15490 ;
    wire new_AGEMA_signal_15491 ;
    wire new_AGEMA_signal_15492 ;
    wire new_AGEMA_signal_15493 ;
    wire new_AGEMA_signal_15494 ;
    wire new_AGEMA_signal_15495 ;
    wire new_AGEMA_signal_15496 ;
    wire new_AGEMA_signal_15497 ;
    wire new_AGEMA_signal_15498 ;
    wire new_AGEMA_signal_15499 ;
    wire new_AGEMA_signal_15500 ;
    wire new_AGEMA_signal_15501 ;
    wire new_AGEMA_signal_15502 ;
    wire new_AGEMA_signal_15503 ;
    wire new_AGEMA_signal_15504 ;
    wire new_AGEMA_signal_15505 ;
    wire new_AGEMA_signal_15506 ;
    wire new_AGEMA_signal_15507 ;
    wire new_AGEMA_signal_15508 ;
    wire new_AGEMA_signal_15509 ;
    wire new_AGEMA_signal_15510 ;
    wire new_AGEMA_signal_15511 ;
    wire new_AGEMA_signal_15512 ;
    wire new_AGEMA_signal_15513 ;
    wire new_AGEMA_signal_15514 ;
    wire new_AGEMA_signal_15515 ;
    wire new_AGEMA_signal_15516 ;
    wire new_AGEMA_signal_15517 ;
    wire new_AGEMA_signal_15518 ;
    wire new_AGEMA_signal_15519 ;
    wire new_AGEMA_signal_15520 ;
    wire new_AGEMA_signal_15521 ;
    wire new_AGEMA_signal_15522 ;
    wire new_AGEMA_signal_15523 ;
    wire new_AGEMA_signal_15524 ;
    wire new_AGEMA_signal_15525 ;
    wire new_AGEMA_signal_15526 ;
    wire new_AGEMA_signal_15527 ;
    wire new_AGEMA_signal_15528 ;
    wire new_AGEMA_signal_15529 ;
    wire new_AGEMA_signal_15530 ;
    wire new_AGEMA_signal_15531 ;
    wire new_AGEMA_signal_15532 ;
    wire new_AGEMA_signal_15533 ;
    wire new_AGEMA_signal_15534 ;
    wire new_AGEMA_signal_15535 ;
    wire new_AGEMA_signal_15536 ;
    wire new_AGEMA_signal_15537 ;
    wire new_AGEMA_signal_15538 ;
    wire new_AGEMA_signal_15539 ;
    wire new_AGEMA_signal_15540 ;
    wire new_AGEMA_signal_15541 ;
    wire new_AGEMA_signal_15542 ;
    wire new_AGEMA_signal_15543 ;
    wire new_AGEMA_signal_15544 ;
    wire new_AGEMA_signal_15545 ;
    wire new_AGEMA_signal_15546 ;
    wire new_AGEMA_signal_15547 ;
    wire new_AGEMA_signal_15548 ;
    wire new_AGEMA_signal_15549 ;
    wire new_AGEMA_signal_15550 ;
    wire new_AGEMA_signal_15551 ;
    wire new_AGEMA_signal_15552 ;
    wire new_AGEMA_signal_15553 ;
    wire new_AGEMA_signal_15554 ;
    wire new_AGEMA_signal_15555 ;
    wire new_AGEMA_signal_15556 ;
    wire new_AGEMA_signal_15557 ;
    wire new_AGEMA_signal_15558 ;
    wire new_AGEMA_signal_15559 ;
    wire new_AGEMA_signal_15560 ;
    wire new_AGEMA_signal_15561 ;
    wire new_AGEMA_signal_15562 ;
    wire new_AGEMA_signal_15563 ;
    wire new_AGEMA_signal_15564 ;
    wire new_AGEMA_signal_15565 ;
    wire new_AGEMA_signal_15566 ;
    wire new_AGEMA_signal_15567 ;
    wire new_AGEMA_signal_15568 ;
    wire new_AGEMA_signal_15569 ;
    wire new_AGEMA_signal_15570 ;
    wire new_AGEMA_signal_15571 ;
    wire new_AGEMA_signal_15572 ;
    wire new_AGEMA_signal_15573 ;
    wire new_AGEMA_signal_15574 ;
    wire new_AGEMA_signal_15575 ;
    wire new_AGEMA_signal_15576 ;
    wire new_AGEMA_signal_15577 ;
    wire new_AGEMA_signal_15578 ;
    wire new_AGEMA_signal_15579 ;
    wire new_AGEMA_signal_15580 ;
    wire new_AGEMA_signal_15581 ;
    wire new_AGEMA_signal_15582 ;
    wire new_AGEMA_signal_15583 ;
    wire new_AGEMA_signal_15584 ;
    wire new_AGEMA_signal_15585 ;
    wire new_AGEMA_signal_15586 ;
    wire new_AGEMA_signal_15587 ;
    wire new_AGEMA_signal_15588 ;
    wire new_AGEMA_signal_15589 ;
    wire new_AGEMA_signal_15590 ;
    wire new_AGEMA_signal_15591 ;
    wire new_AGEMA_signal_15592 ;
    wire new_AGEMA_signal_15593 ;
    wire new_AGEMA_signal_15594 ;
    wire new_AGEMA_signal_15595 ;
    wire new_AGEMA_signal_15596 ;
    wire new_AGEMA_signal_15597 ;
    wire new_AGEMA_signal_15598 ;
    wire new_AGEMA_signal_15599 ;
    wire new_AGEMA_signal_15600 ;
    wire new_AGEMA_signal_15601 ;
    wire new_AGEMA_signal_15602 ;
    wire new_AGEMA_signal_15603 ;
    wire new_AGEMA_signal_15604 ;
    wire new_AGEMA_signal_15605 ;
    wire new_AGEMA_signal_15606 ;
    wire new_AGEMA_signal_15607 ;
    wire new_AGEMA_signal_15608 ;
    wire new_AGEMA_signal_15609 ;
    wire new_AGEMA_signal_15610 ;
    wire new_AGEMA_signal_15611 ;
    wire new_AGEMA_signal_15612 ;
    wire new_AGEMA_signal_15613 ;
    wire new_AGEMA_signal_15614 ;
    wire new_AGEMA_signal_15615 ;
    wire new_AGEMA_signal_15616 ;
    wire new_AGEMA_signal_15617 ;
    wire new_AGEMA_signal_15618 ;
    wire new_AGEMA_signal_15619 ;
    wire new_AGEMA_signal_15620 ;
    wire new_AGEMA_signal_15621 ;
    wire new_AGEMA_signal_15622 ;
    wire new_AGEMA_signal_15623 ;
    wire new_AGEMA_signal_15624 ;
    wire new_AGEMA_signal_15625 ;
    wire new_AGEMA_signal_15626 ;
    wire new_AGEMA_signal_15627 ;
    wire new_AGEMA_signal_15628 ;
    wire new_AGEMA_signal_15629 ;
    wire new_AGEMA_signal_15630 ;
    wire new_AGEMA_signal_15631 ;
    wire new_AGEMA_signal_15632 ;
    wire new_AGEMA_signal_15633 ;
    wire new_AGEMA_signal_15634 ;
    wire new_AGEMA_signal_15635 ;
    wire new_AGEMA_signal_15636 ;
    wire new_AGEMA_signal_15637 ;
    wire new_AGEMA_signal_15638 ;
    wire new_AGEMA_signal_15639 ;
    wire new_AGEMA_signal_15640 ;
    wire new_AGEMA_signal_15641 ;
    wire new_AGEMA_signal_15642 ;
    wire new_AGEMA_signal_15643 ;
    wire new_AGEMA_signal_15644 ;
    wire new_AGEMA_signal_15645 ;
    wire new_AGEMA_signal_15646 ;
    wire new_AGEMA_signal_15647 ;
    wire new_AGEMA_signal_15648 ;
    wire new_AGEMA_signal_15649 ;
    wire new_AGEMA_signal_15650 ;
    wire new_AGEMA_signal_15651 ;
    wire new_AGEMA_signal_15652 ;
    wire new_AGEMA_signal_15653 ;
    wire new_AGEMA_signal_15654 ;
    wire new_AGEMA_signal_15655 ;
    wire new_AGEMA_signal_15656 ;
    wire new_AGEMA_signal_15657 ;
    wire new_AGEMA_signal_15658 ;
    wire new_AGEMA_signal_15659 ;
    wire new_AGEMA_signal_15660 ;
    wire new_AGEMA_signal_15661 ;
    wire new_AGEMA_signal_15662 ;
    wire new_AGEMA_signal_15663 ;
    wire new_AGEMA_signal_15664 ;
    wire new_AGEMA_signal_15665 ;
    wire new_AGEMA_signal_15666 ;
    wire new_AGEMA_signal_15667 ;
    wire new_AGEMA_signal_15668 ;
    wire new_AGEMA_signal_15669 ;
    wire new_AGEMA_signal_15670 ;
    wire new_AGEMA_signal_15671 ;
    wire new_AGEMA_signal_15672 ;
    wire new_AGEMA_signal_15673 ;
    wire new_AGEMA_signal_15674 ;
    wire new_AGEMA_signal_15675 ;
    wire new_AGEMA_signal_15676 ;
    wire new_AGEMA_signal_15677 ;
    wire new_AGEMA_signal_15678 ;
    wire new_AGEMA_signal_15679 ;
    wire new_AGEMA_signal_15680 ;
    wire new_AGEMA_signal_15681 ;
    wire new_AGEMA_signal_15682 ;
    wire new_AGEMA_signal_15683 ;
    wire new_AGEMA_signal_15684 ;
    wire new_AGEMA_signal_15685 ;
    wire new_AGEMA_signal_15686 ;
    wire new_AGEMA_signal_15687 ;
    wire new_AGEMA_signal_15688 ;
    wire new_AGEMA_signal_15689 ;
    wire new_AGEMA_signal_15690 ;
    wire new_AGEMA_signal_15691 ;
    wire new_AGEMA_signal_15692 ;
    wire new_AGEMA_signal_15693 ;
    wire new_AGEMA_signal_15694 ;
    wire new_AGEMA_signal_15695 ;
    wire new_AGEMA_signal_15696 ;
    wire new_AGEMA_signal_15697 ;
    wire new_AGEMA_signal_15698 ;
    wire new_AGEMA_signal_15699 ;
    wire new_AGEMA_signal_15700 ;
    wire new_AGEMA_signal_15701 ;
    wire new_AGEMA_signal_15702 ;
    wire new_AGEMA_signal_15703 ;
    wire new_AGEMA_signal_15704 ;
    wire new_AGEMA_signal_15705 ;
    wire new_AGEMA_signal_15706 ;
    wire new_AGEMA_signal_15707 ;
    wire new_AGEMA_signal_15708 ;
    wire new_AGEMA_signal_15709 ;
    wire new_AGEMA_signal_15710 ;
    wire new_AGEMA_signal_15711 ;
    wire new_AGEMA_signal_15712 ;
    wire new_AGEMA_signal_15713 ;
    wire new_AGEMA_signal_15714 ;
    wire new_AGEMA_signal_15715 ;
    wire new_AGEMA_signal_15716 ;
    wire new_AGEMA_signal_15717 ;
    wire new_AGEMA_signal_15718 ;
    wire new_AGEMA_signal_15719 ;
    wire new_AGEMA_signal_15720 ;
    wire new_AGEMA_signal_15721 ;
    wire new_AGEMA_signal_15722 ;
    wire new_AGEMA_signal_15723 ;
    wire new_AGEMA_signal_15724 ;
    wire new_AGEMA_signal_15725 ;
    wire new_AGEMA_signal_15726 ;
    wire new_AGEMA_signal_15727 ;
    wire new_AGEMA_signal_15728 ;
    wire new_AGEMA_signal_15729 ;
    wire new_AGEMA_signal_15730 ;
    wire new_AGEMA_signal_15731 ;
    wire new_AGEMA_signal_15732 ;
    wire new_AGEMA_signal_15733 ;
    wire new_AGEMA_signal_15734 ;
    wire new_AGEMA_signal_15735 ;
    wire new_AGEMA_signal_15736 ;
    wire new_AGEMA_signal_15737 ;
    wire new_AGEMA_signal_15738 ;
    wire new_AGEMA_signal_15739 ;
    wire new_AGEMA_signal_15740 ;
    wire new_AGEMA_signal_15741 ;
    wire new_AGEMA_signal_15742 ;
    wire new_AGEMA_signal_15743 ;
    wire new_AGEMA_signal_15744 ;
    wire new_AGEMA_signal_15745 ;
    wire new_AGEMA_signal_15746 ;
    wire new_AGEMA_signal_15747 ;
    wire new_AGEMA_signal_15748 ;
    wire new_AGEMA_signal_15749 ;
    wire new_AGEMA_signal_15750 ;
    wire new_AGEMA_signal_15751 ;
    wire new_AGEMA_signal_15752 ;
    wire new_AGEMA_signal_15753 ;
    wire new_AGEMA_signal_15754 ;
    wire new_AGEMA_signal_15755 ;
    wire new_AGEMA_signal_15756 ;
    wire new_AGEMA_signal_15757 ;
    wire new_AGEMA_signal_15758 ;
    wire new_AGEMA_signal_15759 ;
    wire new_AGEMA_signal_15760 ;
    wire new_AGEMA_signal_15761 ;
    wire new_AGEMA_signal_15762 ;
    wire new_AGEMA_signal_15763 ;
    wire new_AGEMA_signal_15764 ;
    wire new_AGEMA_signal_15765 ;
    wire new_AGEMA_signal_15766 ;
    wire new_AGEMA_signal_15767 ;
    wire new_AGEMA_signal_15768 ;
    wire new_AGEMA_signal_15769 ;
    wire new_AGEMA_signal_15770 ;
    wire new_AGEMA_signal_15771 ;
    wire new_AGEMA_signal_15772 ;
    wire new_AGEMA_signal_15773 ;
    wire new_AGEMA_signal_15774 ;
    wire new_AGEMA_signal_15775 ;
    wire new_AGEMA_signal_15776 ;
    wire new_AGEMA_signal_15777 ;
    wire new_AGEMA_signal_15778 ;
    wire new_AGEMA_signal_15779 ;
    wire new_AGEMA_signal_15780 ;
    wire new_AGEMA_signal_15781 ;
    wire new_AGEMA_signal_15782 ;
    wire new_AGEMA_signal_15783 ;
    wire new_AGEMA_signal_15784 ;
    wire new_AGEMA_signal_15785 ;
    wire new_AGEMA_signal_15786 ;
    wire new_AGEMA_signal_15787 ;
    wire new_AGEMA_signal_15788 ;
    wire new_AGEMA_signal_15789 ;
    wire new_AGEMA_signal_15790 ;
    wire new_AGEMA_signal_15791 ;
    wire new_AGEMA_signal_15792 ;
    wire new_AGEMA_signal_15793 ;
    wire new_AGEMA_signal_15794 ;
    wire new_AGEMA_signal_15795 ;
    wire new_AGEMA_signal_15796 ;
    wire new_AGEMA_signal_15797 ;
    wire new_AGEMA_signal_15798 ;
    wire new_AGEMA_signal_15799 ;
    wire new_AGEMA_signal_15800 ;
    wire new_AGEMA_signal_15801 ;
    wire new_AGEMA_signal_15802 ;
    wire new_AGEMA_signal_15803 ;
    wire new_AGEMA_signal_15804 ;
    wire new_AGEMA_signal_15805 ;
    wire new_AGEMA_signal_15806 ;
    wire new_AGEMA_signal_15807 ;
    wire new_AGEMA_signal_15808 ;
    wire new_AGEMA_signal_15809 ;
    wire new_AGEMA_signal_15810 ;
    wire new_AGEMA_signal_15811 ;
    wire new_AGEMA_signal_15812 ;
    wire new_AGEMA_signal_15813 ;
    wire new_AGEMA_signal_15814 ;
    wire new_AGEMA_signal_15815 ;
    wire new_AGEMA_signal_15816 ;
    wire new_AGEMA_signal_15817 ;
    wire new_AGEMA_signal_15818 ;
    wire new_AGEMA_signal_15819 ;
    wire new_AGEMA_signal_15820 ;
    wire new_AGEMA_signal_15821 ;
    wire new_AGEMA_signal_15822 ;
    wire new_AGEMA_signal_15823 ;
    wire new_AGEMA_signal_15824 ;
    wire new_AGEMA_signal_15825 ;
    wire new_AGEMA_signal_15826 ;
    wire new_AGEMA_signal_15827 ;
    wire new_AGEMA_signal_15828 ;
    wire new_AGEMA_signal_15829 ;
    wire new_AGEMA_signal_15830 ;
    wire new_AGEMA_signal_15831 ;
    wire new_AGEMA_signal_15832 ;
    wire new_AGEMA_signal_15833 ;
    wire new_AGEMA_signal_15834 ;
    wire new_AGEMA_signal_15835 ;
    wire new_AGEMA_signal_15836 ;
    wire new_AGEMA_signal_15837 ;
    wire new_AGEMA_signal_15838 ;
    wire new_AGEMA_signal_15839 ;
    wire new_AGEMA_signal_15840 ;
    wire new_AGEMA_signal_15841 ;
    wire new_AGEMA_signal_15842 ;
    wire new_AGEMA_signal_15843 ;
    wire new_AGEMA_signal_15844 ;
    wire new_AGEMA_signal_15845 ;
    wire new_AGEMA_signal_15846 ;
    wire new_AGEMA_signal_15847 ;
    wire new_AGEMA_signal_15848 ;
    wire new_AGEMA_signal_15849 ;
    wire new_AGEMA_signal_15850 ;
    wire new_AGEMA_signal_15851 ;
    wire new_AGEMA_signal_15852 ;
    wire new_AGEMA_signal_15853 ;
    wire new_AGEMA_signal_15854 ;
    wire new_AGEMA_signal_15855 ;
    wire new_AGEMA_signal_15856 ;
    wire new_AGEMA_signal_15857 ;
    wire new_AGEMA_signal_15858 ;
    wire new_AGEMA_signal_15859 ;
    wire new_AGEMA_signal_15860 ;
    wire new_AGEMA_signal_15861 ;
    wire new_AGEMA_signal_15862 ;
    wire new_AGEMA_signal_15863 ;
    wire new_AGEMA_signal_15864 ;
    wire new_AGEMA_signal_15865 ;
    wire new_AGEMA_signal_15866 ;
    wire new_AGEMA_signal_15867 ;
    wire new_AGEMA_signal_15868 ;
    wire new_AGEMA_signal_15869 ;
    wire new_AGEMA_signal_15870 ;
    wire new_AGEMA_signal_15871 ;
    wire new_AGEMA_signal_15872 ;
    wire new_AGEMA_signal_15873 ;
    wire new_AGEMA_signal_15874 ;
    wire new_AGEMA_signal_15875 ;
    wire new_AGEMA_signal_15876 ;
    wire new_AGEMA_signal_15877 ;
    wire new_AGEMA_signal_15878 ;
    wire new_AGEMA_signal_15879 ;
    wire new_AGEMA_signal_15880 ;
    wire new_AGEMA_signal_15881 ;
    wire new_AGEMA_signal_15882 ;
    wire new_AGEMA_signal_15883 ;
    wire new_AGEMA_signal_15884 ;
    wire new_AGEMA_signal_15885 ;
    wire new_AGEMA_signal_15886 ;
    wire new_AGEMA_signal_15887 ;
    wire new_AGEMA_signal_15888 ;
    wire new_AGEMA_signal_15889 ;
    wire new_AGEMA_signal_15890 ;
    wire new_AGEMA_signal_15891 ;
    wire new_AGEMA_signal_15892 ;
    wire new_AGEMA_signal_15893 ;
    wire new_AGEMA_signal_15894 ;
    wire new_AGEMA_signal_15895 ;
    wire new_AGEMA_signal_15896 ;
    wire new_AGEMA_signal_15897 ;
    wire new_AGEMA_signal_15898 ;
    wire new_AGEMA_signal_15899 ;
    wire new_AGEMA_signal_15900 ;
    wire new_AGEMA_signal_15901 ;
    wire new_AGEMA_signal_15902 ;
    wire new_AGEMA_signal_15903 ;
    wire new_AGEMA_signal_15904 ;
    wire new_AGEMA_signal_15905 ;
    wire new_AGEMA_signal_15906 ;
    wire new_AGEMA_signal_15907 ;
    wire new_AGEMA_signal_15908 ;
    wire new_AGEMA_signal_15909 ;
    wire new_AGEMA_signal_15910 ;
    wire new_AGEMA_signal_15911 ;
    wire new_AGEMA_signal_15912 ;
    wire new_AGEMA_signal_15913 ;
    wire new_AGEMA_signal_15914 ;
    wire new_AGEMA_signal_15915 ;
    wire new_AGEMA_signal_15916 ;
    wire new_AGEMA_signal_15917 ;
    wire new_AGEMA_signal_15918 ;
    wire new_AGEMA_signal_15919 ;
    wire new_AGEMA_signal_15920 ;
    wire new_AGEMA_signal_15921 ;
    wire new_AGEMA_signal_15922 ;
    wire new_AGEMA_signal_15923 ;
    wire new_AGEMA_signal_15924 ;
    wire new_AGEMA_signal_15925 ;
    wire new_AGEMA_signal_15926 ;
    wire new_AGEMA_signal_15927 ;
    wire new_AGEMA_signal_15928 ;
    wire new_AGEMA_signal_15929 ;
    wire new_AGEMA_signal_15930 ;
    wire new_AGEMA_signal_15931 ;
    wire new_AGEMA_signal_15932 ;
    wire new_AGEMA_signal_15933 ;
    wire new_AGEMA_signal_15934 ;
    wire new_AGEMA_signal_15935 ;
    wire new_AGEMA_signal_15936 ;
    wire new_AGEMA_signal_15937 ;
    wire new_AGEMA_signal_15938 ;
    wire new_AGEMA_signal_15939 ;
    wire new_AGEMA_signal_15940 ;
    wire new_AGEMA_signal_15941 ;
    wire new_AGEMA_signal_15942 ;
    wire new_AGEMA_signal_15943 ;
    wire new_AGEMA_signal_15944 ;
    wire new_AGEMA_signal_15945 ;
    wire new_AGEMA_signal_15946 ;
    wire new_AGEMA_signal_15947 ;
    wire new_AGEMA_signal_15948 ;
    wire new_AGEMA_signal_15949 ;
    wire new_AGEMA_signal_15950 ;
    wire new_AGEMA_signal_15951 ;
    wire new_AGEMA_signal_15952 ;
    wire new_AGEMA_signal_15953 ;
    wire new_AGEMA_signal_15954 ;
    wire new_AGEMA_signal_15955 ;
    wire new_AGEMA_signal_15956 ;
    wire new_AGEMA_signal_15957 ;
    wire new_AGEMA_signal_15958 ;
    wire new_AGEMA_signal_15959 ;
    wire new_AGEMA_signal_15960 ;
    wire new_AGEMA_signal_15961 ;
    wire new_AGEMA_signal_15962 ;
    wire new_AGEMA_signal_15963 ;
    wire new_AGEMA_signal_15964 ;
    wire new_AGEMA_signal_15965 ;
    wire new_AGEMA_signal_15966 ;
    wire new_AGEMA_signal_15967 ;
    wire new_AGEMA_signal_15968 ;
    wire new_AGEMA_signal_15969 ;
    wire new_AGEMA_signal_15970 ;
    wire new_AGEMA_signal_15971 ;
    wire new_AGEMA_signal_15972 ;
    wire new_AGEMA_signal_15973 ;
    wire new_AGEMA_signal_15974 ;
    wire new_AGEMA_signal_15975 ;
    wire new_AGEMA_signal_15976 ;
    wire new_AGEMA_signal_15977 ;
    wire new_AGEMA_signal_15978 ;
    wire new_AGEMA_signal_15979 ;
    wire new_AGEMA_signal_15980 ;
    wire new_AGEMA_signal_15981 ;
    wire new_AGEMA_signal_15982 ;
    wire new_AGEMA_signal_15983 ;
    wire new_AGEMA_signal_15984 ;
    wire new_AGEMA_signal_15985 ;
    wire new_AGEMA_signal_15986 ;
    wire new_AGEMA_signal_15987 ;
    wire new_AGEMA_signal_15988 ;
    wire new_AGEMA_signal_15989 ;
    wire new_AGEMA_signal_15990 ;
    wire new_AGEMA_signal_15991 ;
    wire new_AGEMA_signal_15992 ;
    wire new_AGEMA_signal_15993 ;
    wire new_AGEMA_signal_15994 ;
    wire new_AGEMA_signal_15995 ;
    wire new_AGEMA_signal_15996 ;
    wire new_AGEMA_signal_15997 ;
    wire new_AGEMA_signal_15998 ;
    wire new_AGEMA_signal_15999 ;
    wire new_AGEMA_signal_16000 ;
    wire new_AGEMA_signal_16001 ;
    wire new_AGEMA_signal_16002 ;
    wire new_AGEMA_signal_16003 ;
    wire new_AGEMA_signal_16004 ;
    wire new_AGEMA_signal_16005 ;
    wire new_AGEMA_signal_16006 ;
    wire new_AGEMA_signal_16007 ;
    wire new_AGEMA_signal_16008 ;
    wire new_AGEMA_signal_16009 ;
    wire new_AGEMA_signal_16010 ;
    wire new_AGEMA_signal_16011 ;
    wire new_AGEMA_signal_16012 ;
    wire new_AGEMA_signal_16013 ;
    wire new_AGEMA_signal_16014 ;
    wire new_AGEMA_signal_16015 ;
    wire new_AGEMA_signal_16016 ;
    wire new_AGEMA_signal_16017 ;
    wire new_AGEMA_signal_16018 ;
    wire new_AGEMA_signal_16019 ;
    wire new_AGEMA_signal_16020 ;
    wire new_AGEMA_signal_16021 ;
    wire new_AGEMA_signal_16022 ;
    wire new_AGEMA_signal_16023 ;
    wire new_AGEMA_signal_16024 ;
    wire new_AGEMA_signal_16025 ;
    wire new_AGEMA_signal_16026 ;
    wire new_AGEMA_signal_16027 ;
    wire new_AGEMA_signal_16028 ;
    wire new_AGEMA_signal_16029 ;
    wire new_AGEMA_signal_16030 ;
    wire new_AGEMA_signal_16031 ;
    wire new_AGEMA_signal_16032 ;
    wire new_AGEMA_signal_16033 ;
    wire new_AGEMA_signal_16034 ;
    wire new_AGEMA_signal_16035 ;
    wire new_AGEMA_signal_16036 ;
    wire new_AGEMA_signal_16037 ;
    wire new_AGEMA_signal_16038 ;
    wire new_AGEMA_signal_16039 ;
    wire new_AGEMA_signal_16040 ;
    wire new_AGEMA_signal_16041 ;
    wire new_AGEMA_signal_16042 ;
    wire new_AGEMA_signal_16043 ;
    wire new_AGEMA_signal_16044 ;
    wire new_AGEMA_signal_16045 ;
    wire new_AGEMA_signal_16046 ;
    wire new_AGEMA_signal_16047 ;
    wire new_AGEMA_signal_16048 ;
    wire new_AGEMA_signal_16049 ;
    wire new_AGEMA_signal_16050 ;
    wire new_AGEMA_signal_16051 ;
    wire new_AGEMA_signal_16052 ;
    wire new_AGEMA_signal_16053 ;
    wire new_AGEMA_signal_16054 ;
    wire new_AGEMA_signal_16055 ;
    wire new_AGEMA_signal_16056 ;
    wire new_AGEMA_signal_16057 ;
    wire new_AGEMA_signal_16058 ;
    wire new_AGEMA_signal_16059 ;
    wire new_AGEMA_signal_16060 ;
    wire new_AGEMA_signal_16061 ;
    wire new_AGEMA_signal_16062 ;
    wire new_AGEMA_signal_16063 ;
    wire new_AGEMA_signal_16064 ;
    wire new_AGEMA_signal_16065 ;
    wire new_AGEMA_signal_16066 ;
    wire new_AGEMA_signal_16067 ;
    wire new_AGEMA_signal_16068 ;
    wire new_AGEMA_signal_16069 ;
    wire new_AGEMA_signal_16070 ;
    wire new_AGEMA_signal_16071 ;
    wire new_AGEMA_signal_16072 ;
    wire new_AGEMA_signal_16073 ;
    wire new_AGEMA_signal_16074 ;
    wire new_AGEMA_signal_16075 ;
    wire new_AGEMA_signal_16076 ;
    wire new_AGEMA_signal_16077 ;
    wire new_AGEMA_signal_16078 ;
    wire new_AGEMA_signal_16079 ;
    wire new_AGEMA_signal_16080 ;
    wire new_AGEMA_signal_16081 ;
    wire new_AGEMA_signal_16082 ;
    wire new_AGEMA_signal_16083 ;
    wire new_AGEMA_signal_16084 ;
    wire new_AGEMA_signal_16085 ;
    wire new_AGEMA_signal_16086 ;
    wire new_AGEMA_signal_16087 ;
    wire new_AGEMA_signal_16088 ;
    wire new_AGEMA_signal_16089 ;
    wire new_AGEMA_signal_16090 ;
    wire new_AGEMA_signal_16091 ;
    wire new_AGEMA_signal_16092 ;
    wire new_AGEMA_signal_16093 ;
    wire new_AGEMA_signal_16094 ;
    wire new_AGEMA_signal_16095 ;
    wire new_AGEMA_signal_16096 ;
    wire new_AGEMA_signal_16097 ;
    wire new_AGEMA_signal_16098 ;
    wire new_AGEMA_signal_16099 ;
    wire new_AGEMA_signal_16100 ;
    wire new_AGEMA_signal_16101 ;
    wire new_AGEMA_signal_16102 ;
    wire new_AGEMA_signal_16103 ;
    wire new_AGEMA_signal_16104 ;
    wire new_AGEMA_signal_16105 ;
    wire new_AGEMA_signal_16106 ;
    wire new_AGEMA_signal_16107 ;
    wire new_AGEMA_signal_16108 ;
    wire new_AGEMA_signal_16109 ;
    wire new_AGEMA_signal_16110 ;
    wire new_AGEMA_signal_16111 ;
    wire new_AGEMA_signal_16112 ;
    wire new_AGEMA_signal_16113 ;
    wire new_AGEMA_signal_16114 ;
    wire new_AGEMA_signal_16115 ;
    wire new_AGEMA_signal_16116 ;
    wire new_AGEMA_signal_16117 ;
    wire new_AGEMA_signal_16118 ;
    wire new_AGEMA_signal_16119 ;
    wire new_AGEMA_signal_16120 ;
    wire new_AGEMA_signal_16121 ;
    wire new_AGEMA_signal_16122 ;
    wire new_AGEMA_signal_16123 ;
    wire new_AGEMA_signal_16124 ;
    wire new_AGEMA_signal_16125 ;
    wire new_AGEMA_signal_16126 ;
    wire new_AGEMA_signal_16127 ;
    wire new_AGEMA_signal_16128 ;
    wire new_AGEMA_signal_16129 ;
    wire new_AGEMA_signal_16130 ;
    wire new_AGEMA_signal_16131 ;
    wire new_AGEMA_signal_16132 ;
    wire new_AGEMA_signal_16133 ;
    wire new_AGEMA_signal_16134 ;
    wire new_AGEMA_signal_16135 ;
    wire new_AGEMA_signal_16136 ;
    wire new_AGEMA_signal_16137 ;
    wire new_AGEMA_signal_16138 ;
    wire new_AGEMA_signal_16139 ;
    wire new_AGEMA_signal_16140 ;
    wire new_AGEMA_signal_16141 ;
    wire new_AGEMA_signal_16142 ;
    wire new_AGEMA_signal_16143 ;
    wire new_AGEMA_signal_16144 ;
    wire new_AGEMA_signal_16145 ;
    wire new_AGEMA_signal_16146 ;
    wire new_AGEMA_signal_16147 ;
    wire new_AGEMA_signal_16148 ;
    wire new_AGEMA_signal_16149 ;
    wire new_AGEMA_signal_16150 ;
    wire new_AGEMA_signal_16151 ;
    wire new_AGEMA_signal_16152 ;
    wire new_AGEMA_signal_16153 ;
    wire new_AGEMA_signal_16154 ;
    wire new_AGEMA_signal_16155 ;
    wire new_AGEMA_signal_16156 ;
    wire new_AGEMA_signal_16157 ;
    wire new_AGEMA_signal_16158 ;
    wire new_AGEMA_signal_16159 ;
    wire new_AGEMA_signal_16160 ;
    wire new_AGEMA_signal_16161 ;
    wire new_AGEMA_signal_16162 ;
    wire new_AGEMA_signal_16163 ;
    wire new_AGEMA_signal_16164 ;
    wire new_AGEMA_signal_16165 ;
    wire new_AGEMA_signal_16166 ;
    wire new_AGEMA_signal_16167 ;
    wire new_AGEMA_signal_16168 ;
    wire new_AGEMA_signal_16169 ;
    wire new_AGEMA_signal_16170 ;
    wire new_AGEMA_signal_16171 ;
    wire new_AGEMA_signal_16172 ;
    wire new_AGEMA_signal_16173 ;
    wire new_AGEMA_signal_16174 ;
    wire new_AGEMA_signal_16175 ;
    wire new_AGEMA_signal_16176 ;
    wire new_AGEMA_signal_16177 ;
    wire new_AGEMA_signal_16178 ;
    wire new_AGEMA_signal_16179 ;
    wire new_AGEMA_signal_16180 ;
    wire new_AGEMA_signal_16181 ;
    wire new_AGEMA_signal_16182 ;
    wire new_AGEMA_signal_16183 ;
    wire new_AGEMA_signal_16184 ;
    wire new_AGEMA_signal_16185 ;
    wire new_AGEMA_signal_16186 ;
    wire new_AGEMA_signal_16187 ;
    wire new_AGEMA_signal_16188 ;
    wire new_AGEMA_signal_16189 ;
    wire new_AGEMA_signal_16190 ;
    wire new_AGEMA_signal_16191 ;
    wire new_AGEMA_signal_16192 ;
    wire new_AGEMA_signal_16193 ;
    wire new_AGEMA_signal_16194 ;
    wire new_AGEMA_signal_16195 ;
    wire new_AGEMA_signal_16196 ;
    wire new_AGEMA_signal_16197 ;
    wire new_AGEMA_signal_16198 ;
    wire new_AGEMA_signal_16199 ;
    wire new_AGEMA_signal_16200 ;
    wire new_AGEMA_signal_16201 ;
    wire new_AGEMA_signal_16202 ;
    wire new_AGEMA_signal_16203 ;
    wire new_AGEMA_signal_16204 ;
    wire new_AGEMA_signal_16205 ;
    wire new_AGEMA_signal_16206 ;
    wire new_AGEMA_signal_16207 ;
    wire new_AGEMA_signal_16208 ;
    wire new_AGEMA_signal_16209 ;
    wire new_AGEMA_signal_16210 ;
    wire new_AGEMA_signal_16211 ;
    wire new_AGEMA_signal_16212 ;
    wire new_AGEMA_signal_16213 ;
    wire new_AGEMA_signal_16214 ;
    wire new_AGEMA_signal_16215 ;
    wire new_AGEMA_signal_16216 ;
    wire new_AGEMA_signal_16217 ;
    wire new_AGEMA_signal_16218 ;
    wire new_AGEMA_signal_16219 ;
    wire new_AGEMA_signal_16220 ;
    wire new_AGEMA_signal_16221 ;
    wire new_AGEMA_signal_16222 ;
    wire new_AGEMA_signal_16223 ;
    wire new_AGEMA_signal_16224 ;
    wire new_AGEMA_signal_16225 ;
    wire new_AGEMA_signal_16226 ;
    wire new_AGEMA_signal_16227 ;
    wire new_AGEMA_signal_16228 ;
    wire new_AGEMA_signal_16229 ;
    wire new_AGEMA_signal_16230 ;
    wire new_AGEMA_signal_16231 ;
    wire new_AGEMA_signal_16232 ;
    wire new_AGEMA_signal_16233 ;
    wire new_AGEMA_signal_16234 ;
    wire new_AGEMA_signal_16235 ;
    wire new_AGEMA_signal_16236 ;
    wire new_AGEMA_signal_16237 ;
    wire new_AGEMA_signal_16238 ;
    wire new_AGEMA_signal_16239 ;
    wire new_AGEMA_signal_16240 ;
    wire new_AGEMA_signal_16241 ;
    wire new_AGEMA_signal_16242 ;
    wire new_AGEMA_signal_16243 ;
    wire new_AGEMA_signal_16244 ;
    wire new_AGEMA_signal_16245 ;
    wire new_AGEMA_signal_16246 ;
    wire new_AGEMA_signal_16247 ;
    wire new_AGEMA_signal_16248 ;
    wire new_AGEMA_signal_16249 ;
    wire new_AGEMA_signal_16250 ;
    wire new_AGEMA_signal_16251 ;
    wire new_AGEMA_signal_16252 ;
    wire new_AGEMA_signal_16253 ;
    wire new_AGEMA_signal_16254 ;
    wire new_AGEMA_signal_16255 ;
    wire new_AGEMA_signal_16256 ;
    wire new_AGEMA_signal_16257 ;
    wire new_AGEMA_signal_16258 ;
    wire new_AGEMA_signal_16259 ;
    wire new_AGEMA_signal_16260 ;
    wire new_AGEMA_signal_16261 ;
    wire new_AGEMA_signal_16262 ;
    wire new_AGEMA_signal_16263 ;
    wire new_AGEMA_signal_16264 ;
    wire new_AGEMA_signal_16265 ;
    wire new_AGEMA_signal_16266 ;
    wire new_AGEMA_signal_16267 ;
    wire new_AGEMA_signal_16268 ;
    wire new_AGEMA_signal_16269 ;
    wire new_AGEMA_signal_16270 ;
    wire new_AGEMA_signal_16271 ;
    wire new_AGEMA_signal_16272 ;
    wire new_AGEMA_signal_16273 ;
    wire new_AGEMA_signal_16274 ;
    wire new_AGEMA_signal_16275 ;
    wire new_AGEMA_signal_16276 ;
    wire new_AGEMA_signal_16277 ;
    wire new_AGEMA_signal_16278 ;
    wire new_AGEMA_signal_16279 ;
    wire new_AGEMA_signal_16280 ;
    wire new_AGEMA_signal_16281 ;
    wire new_AGEMA_signal_16282 ;
    wire new_AGEMA_signal_16283 ;
    wire new_AGEMA_signal_16284 ;
    wire new_AGEMA_signal_16285 ;
    wire new_AGEMA_signal_16286 ;
    wire new_AGEMA_signal_16287 ;
    wire new_AGEMA_signal_16288 ;
    wire new_AGEMA_signal_16289 ;
    wire new_AGEMA_signal_16290 ;
    wire new_AGEMA_signal_16291 ;
    wire new_AGEMA_signal_16292 ;
    wire new_AGEMA_signal_16293 ;
    wire new_AGEMA_signal_16294 ;
    wire new_AGEMA_signal_16295 ;
    wire new_AGEMA_signal_16296 ;
    wire new_AGEMA_signal_16297 ;
    wire new_AGEMA_signal_16298 ;
    wire new_AGEMA_signal_16299 ;
    wire new_AGEMA_signal_16300 ;
    wire new_AGEMA_signal_16301 ;
    wire new_AGEMA_signal_16302 ;
    wire new_AGEMA_signal_16303 ;
    wire new_AGEMA_signal_16304 ;
    wire new_AGEMA_signal_16305 ;
    wire new_AGEMA_signal_16306 ;
    wire new_AGEMA_signal_16307 ;
    wire new_AGEMA_signal_16308 ;
    wire new_AGEMA_signal_16309 ;
    wire new_AGEMA_signal_16310 ;
    wire new_AGEMA_signal_16311 ;
    wire new_AGEMA_signal_16312 ;
    wire new_AGEMA_signal_16313 ;
    wire new_AGEMA_signal_16314 ;
    wire new_AGEMA_signal_16315 ;
    wire new_AGEMA_signal_16316 ;
    wire new_AGEMA_signal_16317 ;
    wire new_AGEMA_signal_16318 ;
    wire new_AGEMA_signal_16319 ;
    wire new_AGEMA_signal_16320 ;
    wire new_AGEMA_signal_16321 ;
    wire new_AGEMA_signal_16322 ;
    wire new_AGEMA_signal_16323 ;
    wire new_AGEMA_signal_16324 ;
    wire new_AGEMA_signal_16325 ;
    wire new_AGEMA_signal_16326 ;
    wire new_AGEMA_signal_16327 ;
    wire new_AGEMA_signal_16328 ;
    wire new_AGEMA_signal_16329 ;
    wire new_AGEMA_signal_16330 ;
    wire new_AGEMA_signal_16331 ;
    wire new_AGEMA_signal_16332 ;
    wire new_AGEMA_signal_16333 ;
    wire new_AGEMA_signal_16334 ;
    wire new_AGEMA_signal_16335 ;
    wire new_AGEMA_signal_16336 ;
    wire new_AGEMA_signal_16337 ;
    wire new_AGEMA_signal_16338 ;
    wire new_AGEMA_signal_16339 ;
    wire new_AGEMA_signal_16340 ;
    wire new_AGEMA_signal_16341 ;
    wire new_AGEMA_signal_16342 ;
    wire new_AGEMA_signal_16343 ;
    wire new_AGEMA_signal_16344 ;
    wire new_AGEMA_signal_16345 ;
    wire new_AGEMA_signal_16346 ;
    wire new_AGEMA_signal_16347 ;
    wire new_AGEMA_signal_16348 ;
    wire new_AGEMA_signal_16349 ;
    wire new_AGEMA_signal_16350 ;
    wire new_AGEMA_signal_16351 ;
    wire new_AGEMA_signal_16352 ;
    wire new_AGEMA_signal_16353 ;
    wire new_AGEMA_signal_16354 ;
    wire new_AGEMA_signal_16355 ;
    wire new_AGEMA_signal_16356 ;
    wire new_AGEMA_signal_16357 ;
    wire new_AGEMA_signal_16358 ;
    wire new_AGEMA_signal_16359 ;
    wire new_AGEMA_signal_16360 ;
    wire new_AGEMA_signal_16361 ;
    wire new_AGEMA_signal_16362 ;
    wire new_AGEMA_signal_16363 ;
    wire new_AGEMA_signal_16364 ;
    wire new_AGEMA_signal_16365 ;
    wire new_AGEMA_signal_16366 ;
    wire new_AGEMA_signal_16367 ;
    wire new_AGEMA_signal_16368 ;
    wire new_AGEMA_signal_16369 ;
    wire new_AGEMA_signal_16370 ;
    wire new_AGEMA_signal_16371 ;
    wire new_AGEMA_signal_16372 ;
    wire new_AGEMA_signal_16373 ;
    wire new_AGEMA_signal_16374 ;
    wire new_AGEMA_signal_16375 ;
    wire new_AGEMA_signal_16376 ;
    wire new_AGEMA_signal_16377 ;
    wire new_AGEMA_signal_16378 ;
    wire new_AGEMA_signal_16379 ;
    wire new_AGEMA_signal_16380 ;
    wire new_AGEMA_signal_16381 ;
    wire new_AGEMA_signal_16382 ;
    wire new_AGEMA_signal_16383 ;
    wire new_AGEMA_signal_16384 ;
    wire new_AGEMA_signal_16385 ;
    wire new_AGEMA_signal_16386 ;
    wire new_AGEMA_signal_16387 ;
    wire new_AGEMA_signal_16388 ;
    wire new_AGEMA_signal_16389 ;
    wire new_AGEMA_signal_16390 ;
    wire new_AGEMA_signal_16391 ;
    wire new_AGEMA_signal_16392 ;
    wire new_AGEMA_signal_16393 ;
    wire new_AGEMA_signal_16394 ;
    wire new_AGEMA_signal_16395 ;
    wire new_AGEMA_signal_16396 ;
    wire new_AGEMA_signal_16397 ;
    wire new_AGEMA_signal_16398 ;
    wire new_AGEMA_signal_16399 ;
    wire new_AGEMA_signal_16400 ;
    wire new_AGEMA_signal_16401 ;
    wire new_AGEMA_signal_16402 ;
    wire new_AGEMA_signal_16403 ;
    wire new_AGEMA_signal_16404 ;
    wire new_AGEMA_signal_16405 ;
    wire new_AGEMA_signal_16406 ;
    wire new_AGEMA_signal_16407 ;
    wire new_AGEMA_signal_16408 ;
    wire new_AGEMA_signal_16409 ;
    wire new_AGEMA_signal_16410 ;
    wire new_AGEMA_signal_16411 ;
    wire new_AGEMA_signal_16412 ;
    wire new_AGEMA_signal_16413 ;
    wire new_AGEMA_signal_16414 ;
    wire new_AGEMA_signal_16415 ;
    wire new_AGEMA_signal_16416 ;
    wire new_AGEMA_signal_16417 ;
    wire new_AGEMA_signal_16418 ;
    wire new_AGEMA_signal_16419 ;
    wire new_AGEMA_signal_16420 ;
    wire new_AGEMA_signal_16421 ;
    wire new_AGEMA_signal_16422 ;
    wire new_AGEMA_signal_16423 ;
    wire new_AGEMA_signal_16424 ;
    wire new_AGEMA_signal_16425 ;
    wire new_AGEMA_signal_16426 ;
    wire new_AGEMA_signal_16427 ;
    wire new_AGEMA_signal_16428 ;
    wire new_AGEMA_signal_16429 ;
    wire new_AGEMA_signal_16430 ;
    wire new_AGEMA_signal_16431 ;
    wire new_AGEMA_signal_16432 ;
    wire new_AGEMA_signal_16433 ;
    wire new_AGEMA_signal_16434 ;
    wire new_AGEMA_signal_16435 ;
    wire new_AGEMA_signal_16436 ;
    wire new_AGEMA_signal_16437 ;
    wire new_AGEMA_signal_16438 ;
    wire new_AGEMA_signal_16439 ;
    wire new_AGEMA_signal_16440 ;
    wire new_AGEMA_signal_16441 ;
    wire new_AGEMA_signal_16442 ;
    wire new_AGEMA_signal_16443 ;
    wire new_AGEMA_signal_16444 ;
    wire new_AGEMA_signal_16445 ;
    wire new_AGEMA_signal_16446 ;
    wire new_AGEMA_signal_16447 ;
    wire new_AGEMA_signal_16448 ;
    wire new_AGEMA_signal_16449 ;
    wire new_AGEMA_signal_16450 ;
    wire new_AGEMA_signal_16451 ;
    wire new_AGEMA_signal_16452 ;
    wire new_AGEMA_signal_16453 ;
    wire new_AGEMA_signal_16454 ;
    wire new_AGEMA_signal_16455 ;
    wire new_AGEMA_signal_16456 ;
    wire new_AGEMA_signal_16457 ;
    wire new_AGEMA_signal_16458 ;
    wire new_AGEMA_signal_16459 ;
    wire new_AGEMA_signal_16460 ;
    wire new_AGEMA_signal_16461 ;
    wire new_AGEMA_signal_16462 ;
    wire new_AGEMA_signal_16463 ;
    wire new_AGEMA_signal_16464 ;
    wire new_AGEMA_signal_16465 ;
    wire new_AGEMA_signal_16466 ;
    wire new_AGEMA_signal_16467 ;
    wire new_AGEMA_signal_16468 ;
    wire new_AGEMA_signal_16469 ;
    wire new_AGEMA_signal_16470 ;
    wire new_AGEMA_signal_16471 ;
    wire new_AGEMA_signal_16472 ;
    wire new_AGEMA_signal_16473 ;
    wire new_AGEMA_signal_16474 ;
    wire new_AGEMA_signal_16475 ;
    wire new_AGEMA_signal_16476 ;
    wire new_AGEMA_signal_16477 ;
    wire new_AGEMA_signal_16478 ;
    wire new_AGEMA_signal_16479 ;
    wire new_AGEMA_signal_16480 ;
    wire new_AGEMA_signal_16481 ;
    wire new_AGEMA_signal_16482 ;
    wire new_AGEMA_signal_16483 ;
    wire new_AGEMA_signal_16484 ;
    wire new_AGEMA_signal_16485 ;
    wire new_AGEMA_signal_16486 ;
    wire new_AGEMA_signal_16487 ;
    wire new_AGEMA_signal_16488 ;
    wire new_AGEMA_signal_16489 ;
    wire new_AGEMA_signal_16490 ;
    wire new_AGEMA_signal_16491 ;
    wire new_AGEMA_signal_16492 ;
    wire new_AGEMA_signal_16493 ;
    wire new_AGEMA_signal_16494 ;
    wire new_AGEMA_signal_16495 ;
    wire new_AGEMA_signal_16496 ;
    wire new_AGEMA_signal_16497 ;
    wire new_AGEMA_signal_16498 ;
    wire new_AGEMA_signal_16499 ;
    wire new_AGEMA_signal_16500 ;
    wire new_AGEMA_signal_16501 ;
    wire new_AGEMA_signal_16502 ;
    wire new_AGEMA_signal_16503 ;
    wire new_AGEMA_signal_16504 ;
    wire new_AGEMA_signal_16505 ;
    wire new_AGEMA_signal_16506 ;
    wire new_AGEMA_signal_16507 ;
    wire new_AGEMA_signal_16508 ;
    wire new_AGEMA_signal_16509 ;
    wire new_AGEMA_signal_16510 ;
    wire new_AGEMA_signal_16511 ;
    wire new_AGEMA_signal_16512 ;
    wire new_AGEMA_signal_16513 ;
    wire new_AGEMA_signal_16514 ;
    wire new_AGEMA_signal_16515 ;
    wire new_AGEMA_signal_16516 ;
    wire new_AGEMA_signal_16517 ;
    wire new_AGEMA_signal_16518 ;
    wire new_AGEMA_signal_16519 ;
    wire new_AGEMA_signal_16520 ;
    wire new_AGEMA_signal_16521 ;
    wire new_AGEMA_signal_16522 ;
    wire new_AGEMA_signal_16523 ;
    wire new_AGEMA_signal_16524 ;
    wire new_AGEMA_signal_16525 ;
    wire new_AGEMA_signal_16526 ;
    wire new_AGEMA_signal_16527 ;
    wire new_AGEMA_signal_16528 ;
    wire new_AGEMA_signal_16529 ;
    wire new_AGEMA_signal_16530 ;
    wire new_AGEMA_signal_16531 ;
    wire new_AGEMA_signal_16532 ;
    wire new_AGEMA_signal_16533 ;
    wire new_AGEMA_signal_16534 ;
    wire new_AGEMA_signal_16535 ;
    wire new_AGEMA_signal_16536 ;
    wire new_AGEMA_signal_16537 ;
    wire new_AGEMA_signal_16538 ;
    wire new_AGEMA_signal_16539 ;
    wire new_AGEMA_signal_16540 ;
    wire new_AGEMA_signal_16541 ;
    wire new_AGEMA_signal_16542 ;
    wire new_AGEMA_signal_16543 ;
    wire new_AGEMA_signal_16544 ;
    wire new_AGEMA_signal_16545 ;
    wire new_AGEMA_signal_16546 ;
    wire new_AGEMA_signal_16547 ;
    wire new_AGEMA_signal_16548 ;
    wire new_AGEMA_signal_16549 ;
    wire new_AGEMA_signal_16550 ;
    wire new_AGEMA_signal_16551 ;
    wire new_AGEMA_signal_16552 ;
    wire new_AGEMA_signal_16553 ;
    wire new_AGEMA_signal_16554 ;
    wire new_AGEMA_signal_16555 ;
    wire new_AGEMA_signal_16556 ;
    wire new_AGEMA_signal_16557 ;
    wire new_AGEMA_signal_16558 ;
    wire new_AGEMA_signal_16559 ;
    wire new_AGEMA_signal_16560 ;
    wire new_AGEMA_signal_16561 ;
    wire new_AGEMA_signal_16562 ;
    wire new_AGEMA_signal_16563 ;
    wire new_AGEMA_signal_16564 ;
    wire new_AGEMA_signal_16565 ;
    wire new_AGEMA_signal_16566 ;
    wire new_AGEMA_signal_16567 ;
    wire new_AGEMA_signal_16568 ;
    wire new_AGEMA_signal_16569 ;
    wire new_AGEMA_signal_16570 ;
    wire new_AGEMA_signal_16571 ;
    wire new_AGEMA_signal_16572 ;
    wire new_AGEMA_signal_16573 ;
    wire new_AGEMA_signal_16574 ;
    wire new_AGEMA_signal_16575 ;
    wire new_AGEMA_signal_16576 ;
    wire new_AGEMA_signal_16577 ;
    wire new_AGEMA_signal_16578 ;
    wire new_AGEMA_signal_16579 ;
    wire new_AGEMA_signal_16580 ;
    wire new_AGEMA_signal_16581 ;
    wire new_AGEMA_signal_16582 ;
    wire new_AGEMA_signal_16583 ;
    wire new_AGEMA_signal_16584 ;
    wire new_AGEMA_signal_16585 ;
    wire new_AGEMA_signal_16586 ;
    wire new_AGEMA_signal_16587 ;
    wire new_AGEMA_signal_16588 ;
    wire new_AGEMA_signal_16589 ;
    wire new_AGEMA_signal_16590 ;
    wire new_AGEMA_signal_16591 ;
    wire new_AGEMA_signal_16592 ;
    wire new_AGEMA_signal_16593 ;
    wire new_AGEMA_signal_16594 ;
    wire new_AGEMA_signal_16595 ;
    wire new_AGEMA_signal_16596 ;
    wire new_AGEMA_signal_16597 ;
    wire new_AGEMA_signal_16598 ;
    wire new_AGEMA_signal_16599 ;
    wire new_AGEMA_signal_16600 ;
    wire new_AGEMA_signal_16601 ;
    wire new_AGEMA_signal_16602 ;
    wire new_AGEMA_signal_16603 ;
    wire new_AGEMA_signal_16604 ;
    wire new_AGEMA_signal_16605 ;
    wire new_AGEMA_signal_16606 ;
    wire new_AGEMA_signal_16607 ;
    wire new_AGEMA_signal_16608 ;
    wire new_AGEMA_signal_16609 ;
    wire new_AGEMA_signal_16610 ;
    wire new_AGEMA_signal_16611 ;
    wire new_AGEMA_signal_16612 ;
    wire new_AGEMA_signal_16613 ;
    wire new_AGEMA_signal_16614 ;
    wire new_AGEMA_signal_16615 ;
    wire new_AGEMA_signal_16616 ;
    wire new_AGEMA_signal_16617 ;
    wire new_AGEMA_signal_16618 ;
    wire new_AGEMA_signal_16619 ;
    wire new_AGEMA_signal_16620 ;
    wire new_AGEMA_signal_16621 ;
    wire new_AGEMA_signal_16622 ;
    wire new_AGEMA_signal_16623 ;
    wire new_AGEMA_signal_16624 ;
    wire new_AGEMA_signal_16625 ;
    wire new_AGEMA_signal_16626 ;
    wire new_AGEMA_signal_16627 ;
    wire new_AGEMA_signal_16628 ;
    wire new_AGEMA_signal_16629 ;
    wire new_AGEMA_signal_16630 ;
    wire new_AGEMA_signal_16631 ;
    wire new_AGEMA_signal_16632 ;
    wire new_AGEMA_signal_16633 ;
    wire new_AGEMA_signal_16634 ;
    wire new_AGEMA_signal_16635 ;
    wire new_AGEMA_signal_16636 ;
    wire new_AGEMA_signal_16637 ;
    wire new_AGEMA_signal_16638 ;
    wire new_AGEMA_signal_16639 ;
    wire new_AGEMA_signal_16640 ;
    wire new_AGEMA_signal_16641 ;
    wire new_AGEMA_signal_16642 ;
    wire new_AGEMA_signal_16643 ;
    wire new_AGEMA_signal_16644 ;
    wire new_AGEMA_signal_16645 ;
    wire new_AGEMA_signal_16646 ;
    wire new_AGEMA_signal_16647 ;
    wire new_AGEMA_signal_16648 ;
    wire new_AGEMA_signal_16649 ;
    wire new_AGEMA_signal_16650 ;
    wire new_AGEMA_signal_16651 ;
    wire new_AGEMA_signal_16652 ;
    wire new_AGEMA_signal_16653 ;
    wire new_AGEMA_signal_16654 ;
    wire new_AGEMA_signal_16655 ;
    wire new_AGEMA_signal_16656 ;
    wire new_AGEMA_signal_16657 ;
    wire new_AGEMA_signal_16658 ;
    wire new_AGEMA_signal_16659 ;
    wire new_AGEMA_signal_16660 ;
    wire new_AGEMA_signal_16661 ;
    wire new_AGEMA_signal_16662 ;
    wire new_AGEMA_signal_16663 ;
    wire new_AGEMA_signal_16664 ;
    wire new_AGEMA_signal_16665 ;
    wire new_AGEMA_signal_16666 ;
    wire new_AGEMA_signal_16667 ;
    wire new_AGEMA_signal_16668 ;
    wire new_AGEMA_signal_16669 ;
    wire new_AGEMA_signal_16670 ;
    wire new_AGEMA_signal_16671 ;
    wire new_AGEMA_signal_16672 ;
    wire new_AGEMA_signal_16673 ;
    wire new_AGEMA_signal_16674 ;
    wire new_AGEMA_signal_16675 ;
    wire new_AGEMA_signal_16676 ;
    wire new_AGEMA_signal_16677 ;
    wire new_AGEMA_signal_16678 ;
    wire new_AGEMA_signal_16679 ;
    wire new_AGEMA_signal_16680 ;
    wire new_AGEMA_signal_16681 ;
    wire new_AGEMA_signal_16682 ;
    wire new_AGEMA_signal_16683 ;
    wire new_AGEMA_signal_16684 ;
    wire new_AGEMA_signal_16685 ;
    wire new_AGEMA_signal_16686 ;
    wire new_AGEMA_signal_16687 ;
    wire new_AGEMA_signal_16688 ;
    wire new_AGEMA_signal_16689 ;
    wire new_AGEMA_signal_16690 ;
    wire new_AGEMA_signal_16691 ;
    wire new_AGEMA_signal_16692 ;
    wire new_AGEMA_signal_16693 ;
    wire new_AGEMA_signal_16694 ;
    wire new_AGEMA_signal_16695 ;
    wire new_AGEMA_signal_16696 ;
    wire new_AGEMA_signal_16697 ;
    wire new_AGEMA_signal_16698 ;
    wire new_AGEMA_signal_16699 ;
    wire new_AGEMA_signal_16700 ;
    wire new_AGEMA_signal_16701 ;
    wire new_AGEMA_signal_16702 ;
    wire new_AGEMA_signal_16703 ;
    wire new_AGEMA_signal_16704 ;
    wire new_AGEMA_signal_16705 ;
    wire new_AGEMA_signal_16706 ;
    wire new_AGEMA_signal_16707 ;
    wire new_AGEMA_signal_16708 ;
    wire new_AGEMA_signal_16709 ;
    wire new_AGEMA_signal_16710 ;
    wire new_AGEMA_signal_16711 ;
    wire new_AGEMA_signal_16712 ;
    wire new_AGEMA_signal_16713 ;
    wire new_AGEMA_signal_16714 ;
    wire new_AGEMA_signal_16715 ;
    wire new_AGEMA_signal_16716 ;
    wire new_AGEMA_signal_16717 ;
    wire new_AGEMA_signal_16718 ;
    wire new_AGEMA_signal_16719 ;
    wire new_AGEMA_signal_16720 ;
    wire new_AGEMA_signal_16721 ;
    wire new_AGEMA_signal_16722 ;
    wire new_AGEMA_signal_16723 ;
    wire new_AGEMA_signal_16724 ;
    wire new_AGEMA_signal_16725 ;
    wire new_AGEMA_signal_16726 ;
    wire new_AGEMA_signal_16727 ;
    wire new_AGEMA_signal_16728 ;
    wire new_AGEMA_signal_16729 ;
    wire new_AGEMA_signal_16730 ;
    wire new_AGEMA_signal_16731 ;
    wire new_AGEMA_signal_16732 ;
    wire new_AGEMA_signal_16733 ;
    wire new_AGEMA_signal_16734 ;
    wire new_AGEMA_signal_16735 ;
    wire new_AGEMA_signal_16736 ;
    wire new_AGEMA_signal_16737 ;
    wire new_AGEMA_signal_16738 ;
    wire new_AGEMA_signal_16739 ;
    wire new_AGEMA_signal_16740 ;
    wire new_AGEMA_signal_16741 ;
    wire new_AGEMA_signal_16742 ;
    wire new_AGEMA_signal_16743 ;
    wire new_AGEMA_signal_16744 ;
    wire new_AGEMA_signal_16745 ;
    wire new_AGEMA_signal_16746 ;
    wire new_AGEMA_signal_16747 ;
    wire new_AGEMA_signal_16748 ;
    wire new_AGEMA_signal_16749 ;
    wire new_AGEMA_signal_16750 ;
    wire new_AGEMA_signal_16751 ;
    wire new_AGEMA_signal_16752 ;
    wire new_AGEMA_signal_16753 ;
    wire new_AGEMA_signal_16754 ;
    wire new_AGEMA_signal_16755 ;
    wire new_AGEMA_signal_16756 ;
    wire new_AGEMA_signal_16757 ;
    wire new_AGEMA_signal_16758 ;
    wire new_AGEMA_signal_16759 ;
    wire new_AGEMA_signal_16760 ;
    wire new_AGEMA_signal_16761 ;
    wire new_AGEMA_signal_16762 ;
    wire new_AGEMA_signal_16763 ;
    wire new_AGEMA_signal_16764 ;
    wire new_AGEMA_signal_16765 ;
    wire new_AGEMA_signal_16766 ;
    wire new_AGEMA_signal_16767 ;
    wire new_AGEMA_signal_16768 ;
    wire new_AGEMA_signal_16769 ;
    wire new_AGEMA_signal_16770 ;
    wire new_AGEMA_signal_16771 ;
    wire new_AGEMA_signal_16772 ;
    wire new_AGEMA_signal_16773 ;
    wire new_AGEMA_signal_16774 ;
    wire new_AGEMA_signal_16775 ;
    wire new_AGEMA_signal_16776 ;
    wire new_AGEMA_signal_16777 ;
    wire new_AGEMA_signal_16778 ;
    wire new_AGEMA_signal_16779 ;
    wire new_AGEMA_signal_16780 ;
    wire new_AGEMA_signal_16781 ;
    wire new_AGEMA_signal_16782 ;
    wire new_AGEMA_signal_16783 ;
    wire new_AGEMA_signal_16784 ;
    wire new_AGEMA_signal_16785 ;
    wire new_AGEMA_signal_16786 ;
    wire new_AGEMA_signal_16787 ;
    wire new_AGEMA_signal_16788 ;
    wire new_AGEMA_signal_16789 ;
    wire new_AGEMA_signal_16790 ;
    wire new_AGEMA_signal_16791 ;
    wire new_AGEMA_signal_16792 ;
    wire new_AGEMA_signal_16793 ;
    wire new_AGEMA_signal_16794 ;
    wire new_AGEMA_signal_16795 ;
    wire new_AGEMA_signal_16796 ;
    wire new_AGEMA_signal_16797 ;
    wire new_AGEMA_signal_16798 ;
    wire new_AGEMA_signal_16799 ;
    wire new_AGEMA_signal_16800 ;
    wire new_AGEMA_signal_16801 ;
    wire new_AGEMA_signal_16802 ;
    wire new_AGEMA_signal_16803 ;
    wire new_AGEMA_signal_16804 ;
    wire new_AGEMA_signal_16805 ;
    wire new_AGEMA_signal_16806 ;
    wire new_AGEMA_signal_16807 ;
    wire new_AGEMA_signal_16808 ;
    wire new_AGEMA_signal_16809 ;
    wire new_AGEMA_signal_16810 ;
    wire new_AGEMA_signal_16811 ;
    wire new_AGEMA_signal_16812 ;
    wire new_AGEMA_signal_16813 ;
    wire new_AGEMA_signal_16814 ;
    wire new_AGEMA_signal_16815 ;
    wire new_AGEMA_signal_16816 ;
    wire new_AGEMA_signal_16817 ;
    wire new_AGEMA_signal_16818 ;
    wire new_AGEMA_signal_16819 ;
    wire new_AGEMA_signal_16820 ;
    wire new_AGEMA_signal_16821 ;
    wire new_AGEMA_signal_16822 ;
    wire new_AGEMA_signal_16823 ;
    wire new_AGEMA_signal_16824 ;
    wire new_AGEMA_signal_16825 ;
    wire new_AGEMA_signal_16826 ;
    wire new_AGEMA_signal_16827 ;
    wire new_AGEMA_signal_16828 ;
    wire new_AGEMA_signal_16829 ;
    wire new_AGEMA_signal_16830 ;
    wire new_AGEMA_signal_16831 ;
    wire new_AGEMA_signal_16832 ;
    wire new_AGEMA_signal_16833 ;
    wire new_AGEMA_signal_16834 ;
    wire new_AGEMA_signal_16835 ;
    wire new_AGEMA_signal_16836 ;
    wire new_AGEMA_signal_16837 ;
    wire new_AGEMA_signal_16838 ;
    wire new_AGEMA_signal_16839 ;
    wire new_AGEMA_signal_16840 ;
    wire new_AGEMA_signal_16841 ;
    wire new_AGEMA_signal_16842 ;
    wire new_AGEMA_signal_16843 ;
    wire new_AGEMA_signal_16844 ;
    wire new_AGEMA_signal_16845 ;
    wire new_AGEMA_signal_16846 ;
    wire new_AGEMA_signal_16847 ;
    wire new_AGEMA_signal_16848 ;
    wire new_AGEMA_signal_16849 ;
    wire new_AGEMA_signal_16850 ;
    wire new_AGEMA_signal_16851 ;
    wire new_AGEMA_signal_16852 ;
    wire new_AGEMA_signal_16853 ;
    wire new_AGEMA_signal_16854 ;
    wire new_AGEMA_signal_16855 ;
    wire new_AGEMA_signal_16856 ;
    wire new_AGEMA_signal_16857 ;
    wire new_AGEMA_signal_16858 ;
    wire new_AGEMA_signal_16859 ;
    wire new_AGEMA_signal_16860 ;
    wire new_AGEMA_signal_16861 ;
    wire new_AGEMA_signal_16862 ;
    wire new_AGEMA_signal_16863 ;
    wire new_AGEMA_signal_16864 ;
    wire new_AGEMA_signal_16865 ;
    wire new_AGEMA_signal_16866 ;
    wire new_AGEMA_signal_16867 ;
    wire new_AGEMA_signal_16868 ;
    wire new_AGEMA_signal_16869 ;
    wire new_AGEMA_signal_16870 ;
    wire new_AGEMA_signal_16871 ;
    wire new_AGEMA_signal_16872 ;
    wire new_AGEMA_signal_16873 ;
    wire new_AGEMA_signal_16874 ;
    wire new_AGEMA_signal_16875 ;
    wire new_AGEMA_signal_16876 ;
    wire new_AGEMA_signal_16877 ;
    wire new_AGEMA_signal_16878 ;
    wire new_AGEMA_signal_16879 ;
    wire new_AGEMA_signal_16880 ;
    wire new_AGEMA_signal_16881 ;
    wire new_AGEMA_signal_16882 ;
    wire new_AGEMA_signal_16883 ;
    wire new_AGEMA_signal_16884 ;
    wire new_AGEMA_signal_16885 ;
    wire new_AGEMA_signal_16886 ;
    wire new_AGEMA_signal_16887 ;
    wire new_AGEMA_signal_16888 ;
    wire new_AGEMA_signal_16889 ;
    wire new_AGEMA_signal_16890 ;
    wire new_AGEMA_signal_16891 ;
    wire new_AGEMA_signal_16892 ;
    wire new_AGEMA_signal_16893 ;
    wire new_AGEMA_signal_16894 ;
    wire new_AGEMA_signal_16895 ;
    wire new_AGEMA_signal_16896 ;
    wire new_AGEMA_signal_16897 ;
    wire new_AGEMA_signal_16898 ;
    wire new_AGEMA_signal_16899 ;
    wire new_AGEMA_signal_16900 ;
    wire new_AGEMA_signal_16901 ;
    wire new_AGEMA_signal_16902 ;
    wire new_AGEMA_signal_16903 ;
    wire new_AGEMA_signal_16904 ;
    wire new_AGEMA_signal_16905 ;
    wire new_AGEMA_signal_16906 ;
    wire new_AGEMA_signal_16907 ;
    wire new_AGEMA_signal_16908 ;
    wire new_AGEMA_signal_16909 ;
    wire new_AGEMA_signal_16910 ;
    wire new_AGEMA_signal_16911 ;
    wire new_AGEMA_signal_16912 ;
    wire new_AGEMA_signal_16913 ;
    wire new_AGEMA_signal_16914 ;
    wire new_AGEMA_signal_16915 ;
    wire new_AGEMA_signal_16916 ;
    wire new_AGEMA_signal_16917 ;
    wire new_AGEMA_signal_16918 ;
    wire new_AGEMA_signal_16919 ;
    wire new_AGEMA_signal_16920 ;
    wire new_AGEMA_signal_16921 ;
    wire new_AGEMA_signal_16922 ;
    wire new_AGEMA_signal_16923 ;
    wire new_AGEMA_signal_16924 ;
    wire new_AGEMA_signal_16925 ;
    wire new_AGEMA_signal_16926 ;
    wire new_AGEMA_signal_16927 ;
    wire new_AGEMA_signal_16928 ;
    wire new_AGEMA_signal_16929 ;
    wire new_AGEMA_signal_16930 ;
    wire new_AGEMA_signal_16931 ;
    wire new_AGEMA_signal_16932 ;
    wire new_AGEMA_signal_16933 ;
    wire new_AGEMA_signal_16934 ;
    wire new_AGEMA_signal_16935 ;
    wire new_AGEMA_signal_16936 ;
    wire new_AGEMA_signal_16937 ;
    wire new_AGEMA_signal_16938 ;
    wire new_AGEMA_signal_16939 ;
    wire new_AGEMA_signal_16940 ;
    wire new_AGEMA_signal_16941 ;
    wire new_AGEMA_signal_16942 ;
    wire new_AGEMA_signal_16943 ;
    wire new_AGEMA_signal_16944 ;
    wire new_AGEMA_signal_16945 ;
    wire new_AGEMA_signal_16946 ;
    wire new_AGEMA_signal_16947 ;
    wire new_AGEMA_signal_16948 ;
    wire new_AGEMA_signal_16949 ;
    wire new_AGEMA_signal_16950 ;
    wire new_AGEMA_signal_16951 ;
    wire new_AGEMA_signal_16952 ;
    wire new_AGEMA_signal_16953 ;
    wire new_AGEMA_signal_16954 ;
    wire new_AGEMA_signal_16955 ;
    wire new_AGEMA_signal_16956 ;
    wire new_AGEMA_signal_16957 ;
    wire new_AGEMA_signal_16958 ;
    wire new_AGEMA_signal_16959 ;
    wire new_AGEMA_signal_16960 ;
    wire new_AGEMA_signal_16961 ;
    wire new_AGEMA_signal_16962 ;
    wire new_AGEMA_signal_16963 ;
    wire new_AGEMA_signal_16964 ;
    wire new_AGEMA_signal_16965 ;
    wire new_AGEMA_signal_16966 ;
    wire new_AGEMA_signal_16967 ;
    wire new_AGEMA_signal_16968 ;
    wire new_AGEMA_signal_16969 ;
    wire new_AGEMA_signal_16970 ;
    wire new_AGEMA_signal_16971 ;
    wire new_AGEMA_signal_16972 ;
    wire new_AGEMA_signal_16973 ;
    wire new_AGEMA_signal_16974 ;
    wire new_AGEMA_signal_16975 ;
    wire new_AGEMA_signal_16976 ;
    wire new_AGEMA_signal_16977 ;
    wire new_AGEMA_signal_16978 ;
    wire new_AGEMA_signal_16979 ;
    wire new_AGEMA_signal_16980 ;
    wire new_AGEMA_signal_16981 ;
    wire new_AGEMA_signal_16982 ;
    wire new_AGEMA_signal_16983 ;
    wire new_AGEMA_signal_16984 ;
    wire new_AGEMA_signal_16985 ;
    wire new_AGEMA_signal_16986 ;
    wire new_AGEMA_signal_16987 ;
    wire new_AGEMA_signal_16988 ;
    wire new_AGEMA_signal_16989 ;
    wire new_AGEMA_signal_16990 ;
    wire new_AGEMA_signal_16991 ;
    wire new_AGEMA_signal_16992 ;
    wire new_AGEMA_signal_16993 ;
    wire new_AGEMA_signal_16994 ;
    wire new_AGEMA_signal_16995 ;
    wire new_AGEMA_signal_16996 ;
    wire new_AGEMA_signal_16997 ;
    wire new_AGEMA_signal_16998 ;
    wire new_AGEMA_signal_16999 ;
    wire new_AGEMA_signal_17000 ;
    wire new_AGEMA_signal_17001 ;
    wire new_AGEMA_signal_17002 ;
    wire new_AGEMA_signal_17003 ;
    wire new_AGEMA_signal_17004 ;
    wire new_AGEMA_signal_17005 ;
    wire new_AGEMA_signal_17006 ;
    wire new_AGEMA_signal_17007 ;
    wire new_AGEMA_signal_17008 ;
    wire new_AGEMA_signal_17009 ;
    wire new_AGEMA_signal_17010 ;
    wire new_AGEMA_signal_17011 ;
    wire new_AGEMA_signal_17012 ;
    wire new_AGEMA_signal_17013 ;
    wire new_AGEMA_signal_17014 ;
    wire new_AGEMA_signal_17015 ;
    wire new_AGEMA_signal_17016 ;
    wire new_AGEMA_signal_17017 ;
    wire new_AGEMA_signal_17018 ;
    wire new_AGEMA_signal_17019 ;
    wire new_AGEMA_signal_17020 ;
    wire new_AGEMA_signal_17021 ;
    wire new_AGEMA_signal_17022 ;
    wire new_AGEMA_signal_17023 ;
    wire new_AGEMA_signal_17024 ;
    wire new_AGEMA_signal_17025 ;
    wire new_AGEMA_signal_17026 ;
    wire new_AGEMA_signal_17027 ;
    wire new_AGEMA_signal_17028 ;
    wire new_AGEMA_signal_17029 ;
    wire new_AGEMA_signal_17030 ;
    wire new_AGEMA_signal_17031 ;
    wire new_AGEMA_signal_17032 ;
    wire new_AGEMA_signal_17033 ;
    wire new_AGEMA_signal_17034 ;
    wire new_AGEMA_signal_17035 ;
    wire new_AGEMA_signal_17036 ;
    wire new_AGEMA_signal_17037 ;
    wire new_AGEMA_signal_17038 ;
    wire new_AGEMA_signal_17039 ;
    wire new_AGEMA_signal_17040 ;
    wire new_AGEMA_signal_17041 ;
    wire new_AGEMA_signal_17042 ;
    wire new_AGEMA_signal_17043 ;
    wire new_AGEMA_signal_17044 ;
    wire new_AGEMA_signal_17045 ;
    wire new_AGEMA_signal_17046 ;
    wire new_AGEMA_signal_17047 ;
    wire new_AGEMA_signal_17048 ;
    wire new_AGEMA_signal_17049 ;
    wire new_AGEMA_signal_17050 ;
    wire new_AGEMA_signal_17051 ;
    wire new_AGEMA_signal_17052 ;
    wire new_AGEMA_signal_17053 ;
    wire new_AGEMA_signal_17054 ;
    wire new_AGEMA_signal_17055 ;
    wire new_AGEMA_signal_17056 ;
    wire new_AGEMA_signal_17057 ;
    wire new_AGEMA_signal_17058 ;
    wire new_AGEMA_signal_17059 ;
    wire new_AGEMA_signal_17060 ;
    wire new_AGEMA_signal_17061 ;
    wire new_AGEMA_signal_17062 ;
    wire new_AGEMA_signal_17063 ;
    wire new_AGEMA_signal_17064 ;
    wire new_AGEMA_signal_17065 ;
    wire new_AGEMA_signal_17066 ;
    wire new_AGEMA_signal_17067 ;
    wire new_AGEMA_signal_17068 ;
    wire new_AGEMA_signal_17069 ;
    wire new_AGEMA_signal_17070 ;
    wire new_AGEMA_signal_17071 ;
    wire new_AGEMA_signal_17072 ;
    wire new_AGEMA_signal_17073 ;
    wire new_AGEMA_signal_17074 ;
    wire new_AGEMA_signal_17075 ;
    wire new_AGEMA_signal_17076 ;
    wire new_AGEMA_signal_17077 ;
    wire new_AGEMA_signal_17078 ;
    wire new_AGEMA_signal_17079 ;
    wire new_AGEMA_signal_17080 ;
    wire new_AGEMA_signal_17081 ;
    wire new_AGEMA_signal_17082 ;
    wire new_AGEMA_signal_17083 ;
    wire new_AGEMA_signal_17084 ;
    wire new_AGEMA_signal_17085 ;
    wire new_AGEMA_signal_17086 ;
    wire new_AGEMA_signal_17087 ;
    wire new_AGEMA_signal_17088 ;
    wire new_AGEMA_signal_17089 ;
    wire new_AGEMA_signal_17090 ;
    wire new_AGEMA_signal_17091 ;
    wire new_AGEMA_signal_17092 ;
    wire new_AGEMA_signal_17093 ;
    wire new_AGEMA_signal_17094 ;
    wire new_AGEMA_signal_17095 ;
    wire new_AGEMA_signal_17096 ;
    wire new_AGEMA_signal_17097 ;
    wire new_AGEMA_signal_17098 ;
    wire new_AGEMA_signal_17099 ;
    wire new_AGEMA_signal_17100 ;
    wire new_AGEMA_signal_17101 ;
    wire new_AGEMA_signal_17102 ;
    wire new_AGEMA_signal_17103 ;
    wire new_AGEMA_signal_17104 ;
    wire new_AGEMA_signal_17105 ;
    wire new_AGEMA_signal_17106 ;
    wire new_AGEMA_signal_17107 ;
    wire new_AGEMA_signal_17108 ;
    wire new_AGEMA_signal_17109 ;
    wire new_AGEMA_signal_17110 ;
    wire new_AGEMA_signal_17111 ;
    wire new_AGEMA_signal_17112 ;
    wire new_AGEMA_signal_17113 ;
    wire new_AGEMA_signal_17114 ;
    wire new_AGEMA_signal_17115 ;
    wire new_AGEMA_signal_17116 ;
    wire new_AGEMA_signal_17117 ;
    wire new_AGEMA_signal_17118 ;
    wire new_AGEMA_signal_17119 ;
    wire new_AGEMA_signal_17120 ;
    wire new_AGEMA_signal_17121 ;
    wire new_AGEMA_signal_17122 ;
    wire new_AGEMA_signal_17123 ;
    wire new_AGEMA_signal_17124 ;
    wire new_AGEMA_signal_17125 ;
    wire new_AGEMA_signal_17126 ;
    wire new_AGEMA_signal_17127 ;
    wire new_AGEMA_signal_17128 ;
    wire new_AGEMA_signal_17129 ;
    wire new_AGEMA_signal_17130 ;
    wire new_AGEMA_signal_17131 ;
    wire new_AGEMA_signal_17132 ;
    wire new_AGEMA_signal_17133 ;
    wire new_AGEMA_signal_17134 ;
    wire new_AGEMA_signal_17135 ;
    wire new_AGEMA_signal_17136 ;
    wire new_AGEMA_signal_17137 ;
    wire new_AGEMA_signal_17138 ;
    wire new_AGEMA_signal_17139 ;
    wire new_AGEMA_signal_17140 ;
    wire new_AGEMA_signal_17141 ;
    wire new_AGEMA_signal_17142 ;
    wire new_AGEMA_signal_17143 ;
    wire new_AGEMA_signal_17144 ;
    wire new_AGEMA_signal_17145 ;
    wire new_AGEMA_signal_17146 ;
    wire new_AGEMA_signal_17147 ;
    wire new_AGEMA_signal_17148 ;
    wire new_AGEMA_signal_17149 ;
    wire new_AGEMA_signal_17150 ;
    wire new_AGEMA_signal_17151 ;
    wire new_AGEMA_signal_17152 ;
    wire new_AGEMA_signal_17153 ;
    wire new_AGEMA_signal_17154 ;
    wire new_AGEMA_signal_17155 ;
    wire new_AGEMA_signal_17156 ;
    wire new_AGEMA_signal_17157 ;
    wire new_AGEMA_signal_17158 ;
    wire new_AGEMA_signal_17159 ;
    wire new_AGEMA_signal_17160 ;
    wire new_AGEMA_signal_17161 ;
    wire new_AGEMA_signal_17162 ;
    wire new_AGEMA_signal_17163 ;
    wire new_AGEMA_signal_17164 ;
    wire new_AGEMA_signal_17165 ;
    wire new_AGEMA_signal_17166 ;
    wire new_AGEMA_signal_17167 ;
    wire new_AGEMA_signal_17168 ;
    wire new_AGEMA_signal_17169 ;
    wire new_AGEMA_signal_17170 ;
    wire new_AGEMA_signal_17171 ;
    wire new_AGEMA_signal_17172 ;
    wire new_AGEMA_signal_17173 ;
    wire new_AGEMA_signal_17174 ;
    wire new_AGEMA_signal_17175 ;
    wire new_AGEMA_signal_17176 ;
    wire new_AGEMA_signal_17177 ;
    wire new_AGEMA_signal_17178 ;
    wire new_AGEMA_signal_17179 ;
    wire new_AGEMA_signal_17180 ;
    wire new_AGEMA_signal_17181 ;
    wire new_AGEMA_signal_17182 ;
    wire new_AGEMA_signal_17183 ;
    wire new_AGEMA_signal_17184 ;
    wire new_AGEMA_signal_17185 ;
    wire new_AGEMA_signal_17186 ;
    wire new_AGEMA_signal_17187 ;
    wire new_AGEMA_signal_17188 ;
    wire new_AGEMA_signal_17189 ;
    wire new_AGEMA_signal_17190 ;
    wire new_AGEMA_signal_17191 ;
    wire new_AGEMA_signal_17192 ;
    wire new_AGEMA_signal_17193 ;
    wire new_AGEMA_signal_17194 ;
    wire new_AGEMA_signal_17195 ;
    wire new_AGEMA_signal_17196 ;
    wire new_AGEMA_signal_17197 ;
    wire new_AGEMA_signal_17198 ;
    wire new_AGEMA_signal_17199 ;
    wire new_AGEMA_signal_17200 ;
    wire new_AGEMA_signal_17201 ;
    wire new_AGEMA_signal_17202 ;
    wire new_AGEMA_signal_17203 ;
    wire new_AGEMA_signal_17204 ;
    wire new_AGEMA_signal_17205 ;
    wire new_AGEMA_signal_17206 ;
    wire new_AGEMA_signal_17207 ;
    wire new_AGEMA_signal_17208 ;
    wire new_AGEMA_signal_17209 ;
    wire new_AGEMA_signal_17210 ;
    wire new_AGEMA_signal_17211 ;
    wire new_AGEMA_signal_17212 ;
    wire new_AGEMA_signal_17213 ;
    wire new_AGEMA_signal_17214 ;
    wire new_AGEMA_signal_17215 ;
    wire new_AGEMA_signal_17216 ;
    wire new_AGEMA_signal_17217 ;
    wire new_AGEMA_signal_17218 ;
    wire new_AGEMA_signal_17219 ;
    wire new_AGEMA_signal_17220 ;
    wire new_AGEMA_signal_17221 ;
    wire new_AGEMA_signal_17222 ;
    wire new_AGEMA_signal_17223 ;
    wire new_AGEMA_signal_17224 ;
    wire new_AGEMA_signal_17225 ;
    wire new_AGEMA_signal_17226 ;
    wire new_AGEMA_signal_17227 ;
    wire new_AGEMA_signal_17228 ;
    wire new_AGEMA_signal_17229 ;
    wire new_AGEMA_signal_17230 ;
    wire new_AGEMA_signal_17231 ;
    wire new_AGEMA_signal_17232 ;
    wire new_AGEMA_signal_17233 ;
    wire new_AGEMA_signal_17234 ;
    wire new_AGEMA_signal_17235 ;
    wire new_AGEMA_signal_17236 ;
    wire new_AGEMA_signal_17237 ;
    wire new_AGEMA_signal_17238 ;
    wire new_AGEMA_signal_17239 ;
    wire new_AGEMA_signal_17240 ;
    wire new_AGEMA_signal_17241 ;
    wire new_AGEMA_signal_17242 ;
    wire new_AGEMA_signal_17243 ;
    wire new_AGEMA_signal_17244 ;
    wire new_AGEMA_signal_17245 ;
    wire new_AGEMA_signal_17246 ;
    wire new_AGEMA_signal_17247 ;
    wire new_AGEMA_signal_17248 ;
    wire new_AGEMA_signal_17249 ;
    wire new_AGEMA_signal_17250 ;
    wire new_AGEMA_signal_17251 ;
    wire new_AGEMA_signal_17252 ;
    wire new_AGEMA_signal_17253 ;
    wire new_AGEMA_signal_17254 ;
    wire new_AGEMA_signal_17255 ;
    wire new_AGEMA_signal_17256 ;
    wire new_AGEMA_signal_17257 ;
    wire new_AGEMA_signal_17258 ;
    wire new_AGEMA_signal_17259 ;
    wire new_AGEMA_signal_17260 ;
    wire new_AGEMA_signal_17261 ;
    wire new_AGEMA_signal_17262 ;
    wire new_AGEMA_signal_17263 ;
    wire new_AGEMA_signal_17264 ;
    wire new_AGEMA_signal_17265 ;
    wire new_AGEMA_signal_17266 ;
    wire new_AGEMA_signal_17267 ;
    wire new_AGEMA_signal_17268 ;
    wire new_AGEMA_signal_17269 ;
    wire new_AGEMA_signal_17270 ;
    wire new_AGEMA_signal_17271 ;
    wire new_AGEMA_signal_17272 ;
    wire new_AGEMA_signal_17273 ;
    wire new_AGEMA_signal_17274 ;
    wire new_AGEMA_signal_17275 ;
    wire new_AGEMA_signal_17276 ;
    wire new_AGEMA_signal_17277 ;
    wire new_AGEMA_signal_17278 ;
    wire new_AGEMA_signal_17279 ;
    wire new_AGEMA_signal_17280 ;
    wire new_AGEMA_signal_17281 ;
    wire new_AGEMA_signal_17282 ;
    wire new_AGEMA_signal_17283 ;
    wire new_AGEMA_signal_17284 ;
    wire new_AGEMA_signal_17285 ;
    wire new_AGEMA_signal_17286 ;
    wire new_AGEMA_signal_17287 ;
    wire new_AGEMA_signal_17288 ;
    wire new_AGEMA_signal_17289 ;
    wire new_AGEMA_signal_17290 ;
    wire new_AGEMA_signal_17291 ;
    wire new_AGEMA_signal_17292 ;
    wire new_AGEMA_signal_17293 ;
    wire new_AGEMA_signal_17294 ;
    wire new_AGEMA_signal_17295 ;
    wire new_AGEMA_signal_17296 ;
    wire new_AGEMA_signal_17297 ;
    wire new_AGEMA_signal_17298 ;
    wire new_AGEMA_signal_17299 ;
    wire new_AGEMA_signal_17300 ;
    wire new_AGEMA_signal_17301 ;
    wire new_AGEMA_signal_17302 ;
    wire new_AGEMA_signal_17303 ;
    wire new_AGEMA_signal_17304 ;
    wire new_AGEMA_signal_17305 ;
    wire new_AGEMA_signal_17306 ;
    wire new_AGEMA_signal_17307 ;
    wire new_AGEMA_signal_17308 ;
    wire new_AGEMA_signal_17309 ;
    wire new_AGEMA_signal_17310 ;
    wire new_AGEMA_signal_17311 ;
    wire new_AGEMA_signal_17312 ;
    wire new_AGEMA_signal_17313 ;
    wire new_AGEMA_signal_17314 ;
    wire new_AGEMA_signal_17315 ;
    wire new_AGEMA_signal_17316 ;
    wire new_AGEMA_signal_17317 ;
    wire new_AGEMA_signal_17318 ;
    wire new_AGEMA_signal_17319 ;
    wire new_AGEMA_signal_17320 ;
    wire new_AGEMA_signal_17321 ;
    wire new_AGEMA_signal_17322 ;
    wire new_AGEMA_signal_17323 ;
    wire new_AGEMA_signal_17324 ;
    wire new_AGEMA_signal_17325 ;
    wire new_AGEMA_signal_17326 ;
    wire new_AGEMA_signal_17327 ;
    wire new_AGEMA_signal_17328 ;
    wire new_AGEMA_signal_17329 ;
    wire new_AGEMA_signal_17330 ;
    wire new_AGEMA_signal_17331 ;
    wire new_AGEMA_signal_17332 ;
    wire new_AGEMA_signal_17333 ;
    wire new_AGEMA_signal_17334 ;
    wire new_AGEMA_signal_17335 ;
    wire new_AGEMA_signal_17336 ;
    wire new_AGEMA_signal_17337 ;
    wire new_AGEMA_signal_17338 ;
    wire new_AGEMA_signal_17339 ;
    wire new_AGEMA_signal_17340 ;
    wire new_AGEMA_signal_17341 ;
    wire new_AGEMA_signal_17342 ;
    wire new_AGEMA_signal_17343 ;
    wire new_AGEMA_signal_17344 ;
    wire new_AGEMA_signal_17345 ;
    wire new_AGEMA_signal_17346 ;
    wire new_AGEMA_signal_17347 ;
    wire new_AGEMA_signal_17348 ;
    wire new_AGEMA_signal_17349 ;
    wire new_AGEMA_signal_17350 ;
    wire new_AGEMA_signal_17351 ;
    wire new_AGEMA_signal_17352 ;
    wire new_AGEMA_signal_17353 ;
    wire new_AGEMA_signal_17354 ;
    wire new_AGEMA_signal_17355 ;
    wire new_AGEMA_signal_17356 ;
    wire new_AGEMA_signal_17357 ;
    wire new_AGEMA_signal_17358 ;
    wire new_AGEMA_signal_17359 ;
    wire new_AGEMA_signal_17360 ;
    wire new_AGEMA_signal_17361 ;
    wire new_AGEMA_signal_17362 ;
    wire new_AGEMA_signal_17363 ;
    wire new_AGEMA_signal_17364 ;
    wire new_AGEMA_signal_17365 ;
    wire new_AGEMA_signal_17366 ;
    wire new_AGEMA_signal_17367 ;
    wire new_AGEMA_signal_17368 ;
    wire new_AGEMA_signal_17369 ;
    wire new_AGEMA_signal_17370 ;
    wire new_AGEMA_signal_17371 ;
    wire new_AGEMA_signal_17372 ;
    wire new_AGEMA_signal_17373 ;
    wire new_AGEMA_signal_17374 ;
    wire new_AGEMA_signal_17375 ;
    wire new_AGEMA_signal_17376 ;
    wire new_AGEMA_signal_17377 ;
    wire new_AGEMA_signal_17378 ;
    wire new_AGEMA_signal_17379 ;
    wire new_AGEMA_signal_17380 ;
    wire new_AGEMA_signal_17381 ;
    wire new_AGEMA_signal_17382 ;
    wire new_AGEMA_signal_17383 ;
    wire new_AGEMA_signal_17384 ;
    wire new_AGEMA_signal_17385 ;
    wire new_AGEMA_signal_17386 ;
    wire new_AGEMA_signal_17387 ;
    wire new_AGEMA_signal_17388 ;
    wire new_AGEMA_signal_17389 ;
    wire new_AGEMA_signal_17390 ;
    wire new_AGEMA_signal_17391 ;
    wire new_AGEMA_signal_17392 ;
    wire new_AGEMA_signal_17393 ;
    wire new_AGEMA_signal_17394 ;
    wire new_AGEMA_signal_17395 ;
    wire new_AGEMA_signal_17396 ;
    wire new_AGEMA_signal_17397 ;
    wire new_AGEMA_signal_17398 ;
    wire new_AGEMA_signal_17399 ;
    wire new_AGEMA_signal_17400 ;
    wire new_AGEMA_signal_17401 ;
    wire new_AGEMA_signal_17402 ;
    wire new_AGEMA_signal_17403 ;
    wire new_AGEMA_signal_17404 ;
    wire new_AGEMA_signal_17405 ;
    wire new_AGEMA_signal_17406 ;
    wire new_AGEMA_signal_17407 ;
    wire new_AGEMA_signal_17408 ;
    wire new_AGEMA_signal_17409 ;
    wire new_AGEMA_signal_17410 ;
    wire new_AGEMA_signal_17411 ;
    wire new_AGEMA_signal_17412 ;
    wire new_AGEMA_signal_17413 ;
    wire new_AGEMA_signal_17414 ;
    wire new_AGEMA_signal_17415 ;
    wire new_AGEMA_signal_17416 ;
    wire new_AGEMA_signal_17417 ;
    wire new_AGEMA_signal_17418 ;
    wire new_AGEMA_signal_17419 ;
    wire new_AGEMA_signal_17420 ;
    wire new_AGEMA_signal_17421 ;
    wire new_AGEMA_signal_17422 ;
    wire new_AGEMA_signal_17423 ;
    wire new_AGEMA_signal_17424 ;
    wire new_AGEMA_signal_17425 ;
    wire new_AGEMA_signal_17426 ;
    wire new_AGEMA_signal_17427 ;
    wire new_AGEMA_signal_17428 ;
    wire new_AGEMA_signal_17429 ;
    wire new_AGEMA_signal_17430 ;
    wire new_AGEMA_signal_17431 ;
    wire new_AGEMA_signal_17432 ;
    wire new_AGEMA_signal_17433 ;
    wire new_AGEMA_signal_17434 ;
    wire new_AGEMA_signal_17435 ;
    wire new_AGEMA_signal_17436 ;
    wire new_AGEMA_signal_17437 ;
    wire new_AGEMA_signal_17438 ;
    wire new_AGEMA_signal_17439 ;
    wire new_AGEMA_signal_17440 ;
    wire new_AGEMA_signal_17441 ;
    wire new_AGEMA_signal_17442 ;
    wire new_AGEMA_signal_17443 ;
    wire new_AGEMA_signal_17444 ;
    wire new_AGEMA_signal_17445 ;
    wire new_AGEMA_signal_17446 ;
    wire new_AGEMA_signal_17447 ;
    wire new_AGEMA_signal_17448 ;
    wire new_AGEMA_signal_17449 ;
    wire new_AGEMA_signal_17450 ;
    wire new_AGEMA_signal_17451 ;
    wire new_AGEMA_signal_17452 ;
    wire new_AGEMA_signal_17453 ;
    wire new_AGEMA_signal_17454 ;
    wire new_AGEMA_signal_17455 ;
    wire new_AGEMA_signal_17456 ;
    wire new_AGEMA_signal_17457 ;
    wire new_AGEMA_signal_17458 ;
    wire new_AGEMA_signal_17459 ;
    wire new_AGEMA_signal_17460 ;
    wire new_AGEMA_signal_17461 ;
    wire new_AGEMA_signal_17462 ;
    wire new_AGEMA_signal_17463 ;
    wire new_AGEMA_signal_17464 ;
    wire new_AGEMA_signal_17465 ;
    wire new_AGEMA_signal_17466 ;
    wire new_AGEMA_signal_17467 ;
    wire new_AGEMA_signal_17471 ;
    wire new_AGEMA_signal_17472 ;
    wire new_AGEMA_signal_17473 ;
    wire new_AGEMA_signal_17474 ;
    wire new_AGEMA_signal_17475 ;
    wire new_AGEMA_signal_17476 ;
    wire new_AGEMA_signal_17483 ;
    wire new_AGEMA_signal_17484 ;
    wire new_AGEMA_signal_17485 ;
    wire new_AGEMA_signal_17486 ;
    wire new_AGEMA_signal_17487 ;
    wire new_AGEMA_signal_17488 ;
    wire new_AGEMA_signal_17489 ;
    wire new_AGEMA_signal_17490 ;
    wire new_AGEMA_signal_17491 ;
    wire new_AGEMA_signal_17492 ;
    wire new_AGEMA_signal_17493 ;
    wire new_AGEMA_signal_17494 ;
    wire new_AGEMA_signal_17495 ;
    wire new_AGEMA_signal_17496 ;
    wire new_AGEMA_signal_17497 ;
    wire new_AGEMA_signal_17498 ;
    wire new_AGEMA_signal_17499 ;
    wire new_AGEMA_signal_17500 ;
    wire new_AGEMA_signal_17501 ;
    wire new_AGEMA_signal_17502 ;
    wire new_AGEMA_signal_17503 ;
    wire new_AGEMA_signal_17504 ;
    wire new_AGEMA_signal_17505 ;
    wire new_AGEMA_signal_17506 ;
    wire new_AGEMA_signal_17507 ;
    wire new_AGEMA_signal_17508 ;
    wire new_AGEMA_signal_17509 ;
    wire new_AGEMA_signal_17510 ;
    wire new_AGEMA_signal_17511 ;
    wire new_AGEMA_signal_17512 ;
    wire new_AGEMA_signal_17513 ;
    wire new_AGEMA_signal_17514 ;
    wire new_AGEMA_signal_17515 ;
    wire new_AGEMA_signal_17516 ;
    wire new_AGEMA_signal_17517 ;
    wire new_AGEMA_signal_17518 ;
    wire new_AGEMA_signal_17519 ;
    wire new_AGEMA_signal_17520 ;
    wire new_AGEMA_signal_17521 ;
    wire new_AGEMA_signal_17522 ;
    wire new_AGEMA_signal_17523 ;
    wire new_AGEMA_signal_17524 ;
    wire new_AGEMA_signal_17525 ;
    wire new_AGEMA_signal_17526 ;
    wire new_AGEMA_signal_17527 ;
    wire new_AGEMA_signal_17528 ;
    wire new_AGEMA_signal_17529 ;
    wire new_AGEMA_signal_17530 ;
    wire new_AGEMA_signal_17531 ;
    wire new_AGEMA_signal_17532 ;
    wire new_AGEMA_signal_17533 ;
    wire new_AGEMA_signal_17534 ;
    wire new_AGEMA_signal_17535 ;
    wire new_AGEMA_signal_17536 ;
    wire new_AGEMA_signal_17537 ;
    wire new_AGEMA_signal_17538 ;
    wire new_AGEMA_signal_17539 ;
    wire new_AGEMA_signal_17540 ;
    wire new_AGEMA_signal_17541 ;
    wire new_AGEMA_signal_17542 ;
    wire new_AGEMA_signal_17543 ;
    wire new_AGEMA_signal_17544 ;
    wire new_AGEMA_signal_17545 ;
    wire new_AGEMA_signal_17546 ;
    wire new_AGEMA_signal_17547 ;
    wire new_AGEMA_signal_17548 ;
    wire new_AGEMA_signal_17549 ;
    wire new_AGEMA_signal_17550 ;
    wire new_AGEMA_signal_17551 ;
    wire new_AGEMA_signal_17552 ;
    wire new_AGEMA_signal_17553 ;
    wire new_AGEMA_signal_17554 ;
    wire new_AGEMA_signal_17555 ;
    wire new_AGEMA_signal_17556 ;
    wire new_AGEMA_signal_17557 ;
    wire new_AGEMA_signal_17558 ;
    wire new_AGEMA_signal_17559 ;
    wire new_AGEMA_signal_17560 ;
    wire new_AGEMA_signal_17561 ;
    wire new_AGEMA_signal_17562 ;
    wire new_AGEMA_signal_17563 ;
    wire new_AGEMA_signal_17564 ;
    wire new_AGEMA_signal_17565 ;
    wire new_AGEMA_signal_17566 ;
    wire new_AGEMA_signal_17567 ;
    wire new_AGEMA_signal_17568 ;
    wire new_AGEMA_signal_17569 ;
    wire new_AGEMA_signal_17570 ;
    wire new_AGEMA_signal_17571 ;
    wire new_AGEMA_signal_17572 ;
    wire new_AGEMA_signal_17573 ;
    wire new_AGEMA_signal_17574 ;
    wire new_AGEMA_signal_17575 ;
    wire new_AGEMA_signal_17576 ;
    wire new_AGEMA_signal_17577 ;
    wire new_AGEMA_signal_17578 ;
    wire new_AGEMA_signal_17579 ;
    wire new_AGEMA_signal_17580 ;
    wire new_AGEMA_signal_17581 ;
    wire new_AGEMA_signal_17582 ;
    wire new_AGEMA_signal_17583 ;
    wire new_AGEMA_signal_17584 ;
    wire new_AGEMA_signal_17585 ;
    wire new_AGEMA_signal_17586 ;
    wire new_AGEMA_signal_17587 ;
    wire new_AGEMA_signal_17588 ;
    wire new_AGEMA_signal_17589 ;
    wire new_AGEMA_signal_17590 ;
    wire new_AGEMA_signal_17591 ;
    wire new_AGEMA_signal_17592 ;
    wire new_AGEMA_signal_17593 ;
    wire new_AGEMA_signal_17594 ;
    wire new_AGEMA_signal_17595 ;
    wire new_AGEMA_signal_17596 ;
    wire new_AGEMA_signal_17597 ;
    wire new_AGEMA_signal_17598 ;
    wire new_AGEMA_signal_17599 ;
    wire new_AGEMA_signal_17600 ;
    wire new_AGEMA_signal_17601 ;
    wire new_AGEMA_signal_17602 ;
    wire new_AGEMA_signal_17603 ;
    wire new_AGEMA_signal_17604 ;
    wire new_AGEMA_signal_17605 ;
    wire new_AGEMA_signal_17606 ;
    wire new_AGEMA_signal_17607 ;
    wire new_AGEMA_signal_17608 ;
    wire new_AGEMA_signal_17609 ;
    wire new_AGEMA_signal_17610 ;
    wire new_AGEMA_signal_17611 ;
    wire new_AGEMA_signal_17612 ;
    wire new_AGEMA_signal_17613 ;
    wire new_AGEMA_signal_17614 ;
    wire new_AGEMA_signal_17615 ;
    wire new_AGEMA_signal_17616 ;
    wire new_AGEMA_signal_17617 ;
    wire new_AGEMA_signal_17618 ;
    wire new_AGEMA_signal_17619 ;
    wire new_AGEMA_signal_17620 ;
    wire new_AGEMA_signal_17621 ;
    wire new_AGEMA_signal_17622 ;
    wire new_AGEMA_signal_17623 ;
    wire new_AGEMA_signal_17624 ;
    wire new_AGEMA_signal_17625 ;
    wire new_AGEMA_signal_17626 ;
    wire new_AGEMA_signal_17627 ;
    wire new_AGEMA_signal_17628 ;
    wire new_AGEMA_signal_17629 ;
    wire new_AGEMA_signal_17630 ;
    wire new_AGEMA_signal_17631 ;
    wire new_AGEMA_signal_17632 ;
    wire new_AGEMA_signal_17633 ;
    wire new_AGEMA_signal_17634 ;
    wire new_AGEMA_signal_17635 ;
    wire new_AGEMA_signal_17636 ;
    wire new_AGEMA_signal_17637 ;
    wire new_AGEMA_signal_17638 ;
    wire new_AGEMA_signal_17639 ;
    wire new_AGEMA_signal_17640 ;
    wire new_AGEMA_signal_17641 ;
    wire new_AGEMA_signal_17642 ;
    wire new_AGEMA_signal_17643 ;
    wire new_AGEMA_signal_17644 ;
    wire new_AGEMA_signal_17645 ;
    wire new_AGEMA_signal_17646 ;
    wire new_AGEMA_signal_17647 ;
    wire new_AGEMA_signal_17648 ;
    wire new_AGEMA_signal_17649 ;
    wire new_AGEMA_signal_17650 ;
    wire new_AGEMA_signal_17651 ;
    wire new_AGEMA_signal_17652 ;
    wire new_AGEMA_signal_17653 ;
    wire new_AGEMA_signal_17654 ;
    wire new_AGEMA_signal_17655 ;
    wire new_AGEMA_signal_17656 ;
    wire new_AGEMA_signal_17657 ;
    wire new_AGEMA_signal_17658 ;
    wire new_AGEMA_signal_17659 ;
    wire new_AGEMA_signal_17660 ;
    wire new_AGEMA_signal_17661 ;
    wire new_AGEMA_signal_17662 ;
    wire new_AGEMA_signal_17663 ;
    wire new_AGEMA_signal_17664 ;
    wire new_AGEMA_signal_17665 ;
    wire new_AGEMA_signal_17666 ;
    wire new_AGEMA_signal_17667 ;
    wire new_AGEMA_signal_17668 ;
    wire new_AGEMA_signal_17669 ;
    wire new_AGEMA_signal_17670 ;
    wire new_AGEMA_signal_17671 ;
    wire new_AGEMA_signal_17672 ;
    wire new_AGEMA_signal_17673 ;
    wire new_AGEMA_signal_17674 ;
    wire new_AGEMA_signal_17675 ;
    wire new_AGEMA_signal_17676 ;
    wire new_AGEMA_signal_17677 ;
    wire new_AGEMA_signal_17678 ;
    wire new_AGEMA_signal_17679 ;
    wire new_AGEMA_signal_17680 ;
    wire new_AGEMA_signal_17681 ;
    wire new_AGEMA_signal_17682 ;
    wire new_AGEMA_signal_17683 ;
    wire new_AGEMA_signal_17684 ;
    wire new_AGEMA_signal_17685 ;
    wire new_AGEMA_signal_17686 ;
    wire new_AGEMA_signal_17687 ;
    wire new_AGEMA_signal_17688 ;
    wire new_AGEMA_signal_17689 ;
    wire new_AGEMA_signal_17690 ;
    wire new_AGEMA_signal_17691 ;
    wire new_AGEMA_signal_17692 ;
    wire new_AGEMA_signal_17693 ;
    wire new_AGEMA_signal_17694 ;
    wire new_AGEMA_signal_17695 ;
    wire new_AGEMA_signal_17696 ;
    wire new_AGEMA_signal_17697 ;
    wire new_AGEMA_signal_17698 ;
    wire new_AGEMA_signal_17699 ;
    wire new_AGEMA_signal_17700 ;
    wire new_AGEMA_signal_17701 ;
    wire new_AGEMA_signal_17702 ;
    wire new_AGEMA_signal_17703 ;
    wire new_AGEMA_signal_17704 ;
    wire new_AGEMA_signal_17705 ;
    wire new_AGEMA_signal_17706 ;
    wire new_AGEMA_signal_17707 ;
    wire new_AGEMA_signal_17708 ;
    wire new_AGEMA_signal_17709 ;
    wire new_AGEMA_signal_17710 ;
    wire new_AGEMA_signal_17711 ;
    wire new_AGEMA_signal_17712 ;
    wire new_AGEMA_signal_17713 ;
    wire new_AGEMA_signal_17714 ;
    wire new_AGEMA_signal_17715 ;
    wire new_AGEMA_signal_17716 ;
    wire new_AGEMA_signal_17717 ;
    wire new_AGEMA_signal_17718 ;
    wire new_AGEMA_signal_17719 ;
    wire new_AGEMA_signal_17720 ;
    wire new_AGEMA_signal_17721 ;
    wire new_AGEMA_signal_17722 ;
    wire new_AGEMA_signal_17723 ;
    wire new_AGEMA_signal_17724 ;
    wire new_AGEMA_signal_17725 ;
    wire new_AGEMA_signal_17726 ;
    wire new_AGEMA_signal_17727 ;
    wire new_AGEMA_signal_17728 ;
    wire new_AGEMA_signal_17729 ;
    wire new_AGEMA_signal_17730 ;
    wire new_AGEMA_signal_17731 ;
    wire new_AGEMA_signal_17732 ;
    wire new_AGEMA_signal_17733 ;
    wire new_AGEMA_signal_17734 ;
    wire new_AGEMA_signal_17735 ;
    wire new_AGEMA_signal_17736 ;
    wire new_AGEMA_signal_17737 ;
    wire new_AGEMA_signal_17738 ;
    wire new_AGEMA_signal_17739 ;
    wire new_AGEMA_signal_17740 ;
    wire new_AGEMA_signal_17741 ;
    wire new_AGEMA_signal_17742 ;
    wire new_AGEMA_signal_17743 ;
    wire new_AGEMA_signal_17744 ;
    wire new_AGEMA_signal_17745 ;
    wire new_AGEMA_signal_17746 ;
    wire new_AGEMA_signal_17747 ;
    wire new_AGEMA_signal_17748 ;
    wire new_AGEMA_signal_17749 ;
    wire new_AGEMA_signal_17750 ;
    wire new_AGEMA_signal_17751 ;
    wire new_AGEMA_signal_17752 ;
    wire new_AGEMA_signal_17753 ;
    wire new_AGEMA_signal_17754 ;
    wire new_AGEMA_signal_17755 ;
    wire new_AGEMA_signal_17756 ;
    wire new_AGEMA_signal_17757 ;
    wire new_AGEMA_signal_17758 ;
    wire new_AGEMA_signal_17759 ;
    wire new_AGEMA_signal_17760 ;
    wire new_AGEMA_signal_17761 ;
    wire new_AGEMA_signal_17762 ;
    wire new_AGEMA_signal_17763 ;
    wire new_AGEMA_signal_17764 ;
    wire new_AGEMA_signal_17765 ;
    wire new_AGEMA_signal_17766 ;
    wire new_AGEMA_signal_17767 ;
    wire new_AGEMA_signal_17768 ;
    wire new_AGEMA_signal_17769 ;
    wire new_AGEMA_signal_17770 ;
    wire new_AGEMA_signal_17771 ;
    wire new_AGEMA_signal_17772 ;
    wire new_AGEMA_signal_17773 ;
    wire new_AGEMA_signal_17774 ;
    wire new_AGEMA_signal_17775 ;
    wire new_AGEMA_signal_17776 ;
    wire new_AGEMA_signal_17777 ;
    wire new_AGEMA_signal_17778 ;
    wire new_AGEMA_signal_17779 ;
    wire new_AGEMA_signal_17780 ;
    wire new_AGEMA_signal_17781 ;
    wire new_AGEMA_signal_17782 ;
    wire new_AGEMA_signal_17783 ;
    wire new_AGEMA_signal_17784 ;
    wire new_AGEMA_signal_17785 ;
    wire new_AGEMA_signal_17786 ;
    wire new_AGEMA_signal_17787 ;
    wire new_AGEMA_signal_17788 ;
    wire new_AGEMA_signal_17789 ;
    wire new_AGEMA_signal_17790 ;
    wire new_AGEMA_signal_17791 ;
    wire new_AGEMA_signal_17792 ;
    wire new_AGEMA_signal_17793 ;
    wire new_AGEMA_signal_17794 ;
    wire new_AGEMA_signal_17798 ;
    wire new_AGEMA_signal_17799 ;
    wire new_AGEMA_signal_17800 ;
    wire new_AGEMA_signal_17801 ;
    wire new_AGEMA_signal_17802 ;
    wire new_AGEMA_signal_17803 ;
    wire new_AGEMA_signal_17810 ;
    wire new_AGEMA_signal_17811 ;
    wire new_AGEMA_signal_17812 ;
    wire new_AGEMA_signal_17813 ;
    wire new_AGEMA_signal_17814 ;
    wire new_AGEMA_signal_17815 ;
    wire new_AGEMA_signal_17816 ;
    wire new_AGEMA_signal_17817 ;
    wire new_AGEMA_signal_17818 ;
    wire new_AGEMA_signal_17819 ;
    wire new_AGEMA_signal_17820 ;
    wire new_AGEMA_signal_17821 ;
    wire new_AGEMA_signal_17822 ;
    wire new_AGEMA_signal_17823 ;
    wire new_AGEMA_signal_17824 ;
    wire new_AGEMA_signal_17825 ;
    wire new_AGEMA_signal_17826 ;
    wire new_AGEMA_signal_17827 ;
    wire new_AGEMA_signal_17828 ;
    wire new_AGEMA_signal_17829 ;
    wire new_AGEMA_signal_17830 ;
    wire new_AGEMA_signal_17831 ;
    wire new_AGEMA_signal_17832 ;
    wire new_AGEMA_signal_17833 ;
    wire new_AGEMA_signal_17834 ;
    wire new_AGEMA_signal_17835 ;
    wire new_AGEMA_signal_17836 ;
    wire new_AGEMA_signal_17837 ;
    wire new_AGEMA_signal_17838 ;
    wire new_AGEMA_signal_17839 ;
    wire new_AGEMA_signal_17840 ;
    wire new_AGEMA_signal_17841 ;
    wire new_AGEMA_signal_17842 ;
    wire new_AGEMA_signal_17843 ;
    wire new_AGEMA_signal_17844 ;
    wire new_AGEMA_signal_17845 ;
    wire new_AGEMA_signal_17846 ;
    wire new_AGEMA_signal_17847 ;
    wire new_AGEMA_signal_17848 ;
    wire new_AGEMA_signal_17849 ;
    wire new_AGEMA_signal_17850 ;
    wire new_AGEMA_signal_17851 ;
    wire new_AGEMA_signal_17852 ;
    wire new_AGEMA_signal_17853 ;
    wire new_AGEMA_signal_17854 ;
    wire new_AGEMA_signal_17855 ;
    wire new_AGEMA_signal_17856 ;
    wire new_AGEMA_signal_17857 ;
    wire new_AGEMA_signal_17858 ;
    wire new_AGEMA_signal_17859 ;
    wire new_AGEMA_signal_17860 ;
    wire new_AGEMA_signal_17861 ;
    wire new_AGEMA_signal_17862 ;
    wire new_AGEMA_signal_17863 ;
    wire new_AGEMA_signal_17864 ;
    wire new_AGEMA_signal_17865 ;
    wire new_AGEMA_signal_17866 ;
    wire new_AGEMA_signal_17867 ;
    wire new_AGEMA_signal_17868 ;
    wire new_AGEMA_signal_17869 ;
    wire new_AGEMA_signal_17870 ;
    wire new_AGEMA_signal_17871 ;
    wire new_AGEMA_signal_17872 ;
    wire new_AGEMA_signal_17873 ;
    wire new_AGEMA_signal_17874 ;
    wire new_AGEMA_signal_17875 ;
    wire new_AGEMA_signal_17876 ;
    wire new_AGEMA_signal_17877 ;
    wire new_AGEMA_signal_17878 ;
    wire new_AGEMA_signal_17879 ;
    wire new_AGEMA_signal_17880 ;
    wire new_AGEMA_signal_17881 ;
    wire new_AGEMA_signal_17882 ;
    wire new_AGEMA_signal_17883 ;
    wire new_AGEMA_signal_17884 ;
    wire new_AGEMA_signal_17885 ;
    wire new_AGEMA_signal_17886 ;
    wire new_AGEMA_signal_17887 ;
    wire new_AGEMA_signal_17888 ;
    wire new_AGEMA_signal_17889 ;
    wire new_AGEMA_signal_17890 ;
    wire new_AGEMA_signal_17891 ;
    wire new_AGEMA_signal_17892 ;
    wire new_AGEMA_signal_17893 ;
    wire new_AGEMA_signal_17894 ;
    wire new_AGEMA_signal_17895 ;
    wire new_AGEMA_signal_17896 ;
    wire new_AGEMA_signal_17897 ;
    wire new_AGEMA_signal_17898 ;
    wire new_AGEMA_signal_17899 ;
    wire new_AGEMA_signal_17900 ;
    wire new_AGEMA_signal_17901 ;
    wire new_AGEMA_signal_17902 ;
    wire new_AGEMA_signal_17903 ;
    wire new_AGEMA_signal_17904 ;
    wire new_AGEMA_signal_17905 ;
    wire new_AGEMA_signal_17906 ;
    wire new_AGEMA_signal_17907 ;
    wire new_AGEMA_signal_17908 ;
    wire new_AGEMA_signal_17909 ;
    wire new_AGEMA_signal_17910 ;
    wire new_AGEMA_signal_17911 ;
    wire new_AGEMA_signal_17912 ;
    wire new_AGEMA_signal_17913 ;
    wire new_AGEMA_signal_17914 ;
    wire new_AGEMA_signal_17915 ;
    wire new_AGEMA_signal_17916 ;
    wire new_AGEMA_signal_17917 ;
    wire new_AGEMA_signal_17918 ;
    wire new_AGEMA_signal_17919 ;
    wire new_AGEMA_signal_17920 ;
    wire new_AGEMA_signal_17921 ;
    wire new_AGEMA_signal_17922 ;
    wire new_AGEMA_signal_17923 ;
    wire new_AGEMA_signal_17924 ;
    wire new_AGEMA_signal_17925 ;
    wire new_AGEMA_signal_17926 ;
    wire new_AGEMA_signal_17927 ;
    wire new_AGEMA_signal_17928 ;
    wire new_AGEMA_signal_17929 ;
    wire new_AGEMA_signal_17930 ;
    wire new_AGEMA_signal_17931 ;
    wire new_AGEMA_signal_17932 ;
    wire new_AGEMA_signal_17933 ;
    wire new_AGEMA_signal_17934 ;
    wire new_AGEMA_signal_17935 ;
    wire new_AGEMA_signal_17936 ;
    wire new_AGEMA_signal_17937 ;
    wire new_AGEMA_signal_17938 ;
    wire new_AGEMA_signal_17939 ;
    wire new_AGEMA_signal_17940 ;
    wire new_AGEMA_signal_17941 ;
    wire new_AGEMA_signal_17942 ;
    wire new_AGEMA_signal_17943 ;
    wire new_AGEMA_signal_17944 ;
    wire new_AGEMA_signal_17945 ;
    wire new_AGEMA_signal_17946 ;
    wire new_AGEMA_signal_17947 ;
    wire new_AGEMA_signal_17948 ;
    wire new_AGEMA_signal_17949 ;
    wire new_AGEMA_signal_17950 ;
    wire new_AGEMA_signal_17951 ;
    wire new_AGEMA_signal_17952 ;
    wire new_AGEMA_signal_17953 ;
    wire new_AGEMA_signal_17954 ;
    wire new_AGEMA_signal_17955 ;
    wire new_AGEMA_signal_17956 ;
    wire new_AGEMA_signal_17957 ;
    wire new_AGEMA_signal_17958 ;
    wire new_AGEMA_signal_17959 ;
    wire new_AGEMA_signal_17960 ;
    wire new_AGEMA_signal_17961 ;
    wire new_AGEMA_signal_17962 ;
    wire new_AGEMA_signal_17963 ;
    wire new_AGEMA_signal_17964 ;
    wire new_AGEMA_signal_17965 ;
    wire new_AGEMA_signal_17966 ;
    wire new_AGEMA_signal_17967 ;
    wire new_AGEMA_signal_17968 ;
    wire new_AGEMA_signal_17969 ;
    wire new_AGEMA_signal_17970 ;
    wire new_AGEMA_signal_17971 ;
    wire new_AGEMA_signal_17972 ;
    wire new_AGEMA_signal_17973 ;
    wire new_AGEMA_signal_17974 ;
    wire new_AGEMA_signal_17975 ;
    wire new_AGEMA_signal_17976 ;
    wire new_AGEMA_signal_17977 ;
    wire new_AGEMA_signal_17978 ;
    wire new_AGEMA_signal_17979 ;
    wire new_AGEMA_signal_17980 ;
    wire new_AGEMA_signal_17981 ;
    wire new_AGEMA_signal_17982 ;
    wire new_AGEMA_signal_17983 ;
    wire new_AGEMA_signal_17984 ;
    wire new_AGEMA_signal_17985 ;
    wire new_AGEMA_signal_17986 ;
    wire new_AGEMA_signal_17987 ;
    wire new_AGEMA_signal_17988 ;
    wire new_AGEMA_signal_17989 ;
    wire new_AGEMA_signal_17990 ;
    wire new_AGEMA_signal_17991 ;
    wire new_AGEMA_signal_17992 ;
    wire new_AGEMA_signal_17993 ;
    wire new_AGEMA_signal_17994 ;
    wire new_AGEMA_signal_17995 ;
    wire new_AGEMA_signal_17996 ;
    wire new_AGEMA_signal_17997 ;
    wire new_AGEMA_signal_17998 ;
    wire new_AGEMA_signal_17999 ;
    wire new_AGEMA_signal_18000 ;
    wire new_AGEMA_signal_18001 ;
    wire new_AGEMA_signal_18002 ;
    wire new_AGEMA_signal_18003 ;
    wire new_AGEMA_signal_18004 ;
    wire new_AGEMA_signal_18005 ;
    wire new_AGEMA_signal_18006 ;
    wire new_AGEMA_signal_18007 ;
    wire new_AGEMA_signal_18008 ;
    wire new_AGEMA_signal_18009 ;
    wire new_AGEMA_signal_18010 ;
    wire new_AGEMA_signal_18011 ;
    wire new_AGEMA_signal_18012 ;
    wire new_AGEMA_signal_18013 ;
    wire new_AGEMA_signal_18014 ;
    wire new_AGEMA_signal_18015 ;
    wire new_AGEMA_signal_18016 ;
    wire new_AGEMA_signal_18017 ;
    wire new_AGEMA_signal_18018 ;
    wire new_AGEMA_signal_18019 ;
    wire new_AGEMA_signal_18020 ;
    wire new_AGEMA_signal_18021 ;
    wire new_AGEMA_signal_18022 ;
    wire new_AGEMA_signal_18023 ;
    wire new_AGEMA_signal_18024 ;
    wire new_AGEMA_signal_18025 ;
    wire new_AGEMA_signal_18026 ;
    wire new_AGEMA_signal_18027 ;
    wire new_AGEMA_signal_18028 ;
    wire new_AGEMA_signal_18029 ;
    wire new_AGEMA_signal_18030 ;
    wire new_AGEMA_signal_18031 ;
    wire new_AGEMA_signal_18032 ;
    wire new_AGEMA_signal_18033 ;
    wire new_AGEMA_signal_18034 ;
    wire new_AGEMA_signal_18035 ;
    wire new_AGEMA_signal_18036 ;
    wire new_AGEMA_signal_18037 ;
    wire new_AGEMA_signal_18038 ;
    wire new_AGEMA_signal_18039 ;
    wire new_AGEMA_signal_18040 ;
    wire new_AGEMA_signal_18041 ;
    wire new_AGEMA_signal_18042 ;
    wire new_AGEMA_signal_18043 ;
    wire new_AGEMA_signal_18050 ;
    wire new_AGEMA_signal_18051 ;
    wire new_AGEMA_signal_18052 ;
    wire new_AGEMA_signal_18053 ;
    wire new_AGEMA_signal_18054 ;
    wire new_AGEMA_signal_18055 ;
    wire new_AGEMA_signal_18056 ;
    wire new_AGEMA_signal_18057 ;
    wire new_AGEMA_signal_18058 ;
    wire new_AGEMA_signal_18059 ;
    wire new_AGEMA_signal_18060 ;
    wire new_AGEMA_signal_18061 ;
    wire new_AGEMA_signal_18062 ;
    wire new_AGEMA_signal_18063 ;
    wire new_AGEMA_signal_18064 ;
    wire new_AGEMA_signal_18065 ;
    wire new_AGEMA_signal_18066 ;
    wire new_AGEMA_signal_18067 ;
    wire new_AGEMA_signal_18068 ;
    wire new_AGEMA_signal_18069 ;
    wire new_AGEMA_signal_18070 ;
    wire new_AGEMA_signal_18071 ;
    wire new_AGEMA_signal_18072 ;
    wire new_AGEMA_signal_18073 ;
    wire new_AGEMA_signal_18074 ;
    wire new_AGEMA_signal_18075 ;
    wire new_AGEMA_signal_18076 ;
    wire new_AGEMA_signal_18077 ;
    wire new_AGEMA_signal_18078 ;
    wire new_AGEMA_signal_18079 ;
    wire new_AGEMA_signal_18116 ;
    wire new_AGEMA_signal_18117 ;
    wire new_AGEMA_signal_18118 ;
    wire new_AGEMA_signal_18119 ;
    wire new_AGEMA_signal_18120 ;
    wire new_AGEMA_signal_18121 ;
    wire new_AGEMA_signal_18122 ;
    wire new_AGEMA_signal_18123 ;
    wire new_AGEMA_signal_18124 ;
    wire new_AGEMA_signal_18125 ;
    wire new_AGEMA_signal_18126 ;
    wire new_AGEMA_signal_18127 ;
    wire new_AGEMA_signal_18128 ;
    wire new_AGEMA_signal_18129 ;
    wire new_AGEMA_signal_18130 ;
    wire new_AGEMA_signal_18131 ;
    wire new_AGEMA_signal_18132 ;
    wire new_AGEMA_signal_18133 ;
    wire new_AGEMA_signal_18137 ;
    wire new_AGEMA_signal_18138 ;
    wire new_AGEMA_signal_18139 ;
    wire new_AGEMA_signal_18140 ;
    wire new_AGEMA_signal_18141 ;
    wire new_AGEMA_signal_18142 ;
    wire new_AGEMA_signal_18143 ;
    wire new_AGEMA_signal_18144 ;
    wire new_AGEMA_signal_18145 ;
    wire new_AGEMA_signal_18146 ;
    wire new_AGEMA_signal_18147 ;
    wire new_AGEMA_signal_18148 ;
    wire new_AGEMA_signal_18149 ;
    wire new_AGEMA_signal_18150 ;
    wire new_AGEMA_signal_18151 ;
    wire new_AGEMA_signal_18152 ;
    wire new_AGEMA_signal_18153 ;
    wire new_AGEMA_signal_18154 ;
    wire new_AGEMA_signal_18155 ;
    wire new_AGEMA_signal_18156 ;
    wire new_AGEMA_signal_18157 ;
    wire new_AGEMA_signal_18158 ;
    wire new_AGEMA_signal_18159 ;
    wire new_AGEMA_signal_18160 ;
    wire new_AGEMA_signal_18161 ;
    wire new_AGEMA_signal_18162 ;
    wire new_AGEMA_signal_18163 ;
    wire new_AGEMA_signal_18164 ;
    wire new_AGEMA_signal_18165 ;
    wire new_AGEMA_signal_18166 ;
    wire new_AGEMA_signal_18167 ;
    wire new_AGEMA_signal_18168 ;
    wire new_AGEMA_signal_18169 ;
    wire new_AGEMA_signal_18170 ;
    wire new_AGEMA_signal_18171 ;
    wire new_AGEMA_signal_18172 ;
    wire new_AGEMA_signal_18173 ;
    wire new_AGEMA_signal_18174 ;
    wire new_AGEMA_signal_18175 ;
    wire new_AGEMA_signal_18176 ;
    wire new_AGEMA_signal_18177 ;
    wire new_AGEMA_signal_18178 ;
    wire new_AGEMA_signal_18179 ;
    wire new_AGEMA_signal_18180 ;
    wire new_AGEMA_signal_18181 ;
    wire new_AGEMA_signal_18182 ;
    wire new_AGEMA_signal_18183 ;
    wire new_AGEMA_signal_18184 ;
    wire new_AGEMA_signal_18185 ;
    wire new_AGEMA_signal_18186 ;
    wire new_AGEMA_signal_18187 ;
    wire new_AGEMA_signal_18188 ;
    wire new_AGEMA_signal_18189 ;
    wire new_AGEMA_signal_18190 ;
    wire new_AGEMA_signal_18191 ;
    wire new_AGEMA_signal_18192 ;
    wire new_AGEMA_signal_18193 ;
    wire new_AGEMA_signal_18194 ;
    wire new_AGEMA_signal_18195 ;
    wire new_AGEMA_signal_18196 ;
    wire new_AGEMA_signal_18197 ;
    wire new_AGEMA_signal_18198 ;
    wire new_AGEMA_signal_18199 ;
    wire new_AGEMA_signal_18200 ;
    wire new_AGEMA_signal_18201 ;
    wire new_AGEMA_signal_18202 ;
    wire new_AGEMA_signal_18203 ;
    wire new_AGEMA_signal_18204 ;
    wire new_AGEMA_signal_18205 ;
    wire new_AGEMA_signal_18206 ;
    wire new_AGEMA_signal_18207 ;
    wire new_AGEMA_signal_18208 ;
    wire new_AGEMA_signal_18209 ;
    wire new_AGEMA_signal_18210 ;
    wire new_AGEMA_signal_18211 ;
    wire new_AGEMA_signal_18212 ;
    wire new_AGEMA_signal_18213 ;
    wire new_AGEMA_signal_18214 ;
    wire new_AGEMA_signal_18215 ;
    wire new_AGEMA_signal_18216 ;
    wire new_AGEMA_signal_18217 ;
    wire new_AGEMA_signal_18218 ;
    wire new_AGEMA_signal_18219 ;
    wire new_AGEMA_signal_18220 ;
    wire new_AGEMA_signal_18221 ;
    wire new_AGEMA_signal_18222 ;
    wire new_AGEMA_signal_18223 ;
    wire new_AGEMA_signal_18224 ;
    wire new_AGEMA_signal_18225 ;
    wire new_AGEMA_signal_18226 ;
    wire new_AGEMA_signal_18227 ;
    wire new_AGEMA_signal_18228 ;
    wire new_AGEMA_signal_18229 ;
    wire new_AGEMA_signal_18230 ;
    wire new_AGEMA_signal_18231 ;
    wire new_AGEMA_signal_18232 ;
    wire new_AGEMA_signal_18233 ;
    wire new_AGEMA_signal_18234 ;
    wire new_AGEMA_signal_18235 ;
    wire new_AGEMA_signal_18236 ;
    wire new_AGEMA_signal_18237 ;
    wire new_AGEMA_signal_18238 ;
    wire new_AGEMA_signal_18239 ;
    wire new_AGEMA_signal_18240 ;
    wire new_AGEMA_signal_18241 ;
    wire new_AGEMA_signal_18242 ;
    wire new_AGEMA_signal_18243 ;
    wire new_AGEMA_signal_18244 ;
    wire new_AGEMA_signal_18245 ;
    wire new_AGEMA_signal_18246 ;
    wire new_AGEMA_signal_18247 ;
    wire new_AGEMA_signal_18248 ;
    wire new_AGEMA_signal_18249 ;
    wire new_AGEMA_signal_18250 ;
    wire new_AGEMA_signal_18251 ;
    wire new_AGEMA_signal_18252 ;
    wire new_AGEMA_signal_18253 ;
    wire new_AGEMA_signal_18254 ;
    wire new_AGEMA_signal_18255 ;
    wire new_AGEMA_signal_18256 ;
    wire new_AGEMA_signal_18257 ;
    wire new_AGEMA_signal_18258 ;
    wire new_AGEMA_signal_18259 ;
    wire new_AGEMA_signal_18260 ;
    wire new_AGEMA_signal_18261 ;
    wire new_AGEMA_signal_18262 ;
    wire new_AGEMA_signal_18266 ;
    wire new_AGEMA_signal_18267 ;
    wire new_AGEMA_signal_18268 ;
    wire new_AGEMA_signal_18269 ;
    wire new_AGEMA_signal_18270 ;
    wire new_AGEMA_signal_18271 ;
    wire new_AGEMA_signal_18272 ;
    wire new_AGEMA_signal_18273 ;
    wire new_AGEMA_signal_18274 ;
    wire new_AGEMA_signal_18275 ;
    wire new_AGEMA_signal_18276 ;
    wire new_AGEMA_signal_18277 ;
    wire new_AGEMA_signal_18278 ;
    wire new_AGEMA_signal_18279 ;
    wire new_AGEMA_signal_18280 ;
    wire new_AGEMA_signal_18281 ;
    wire new_AGEMA_signal_18282 ;
    wire new_AGEMA_signal_18283 ;
    wire new_AGEMA_signal_18284 ;
    wire new_AGEMA_signal_18285 ;
    wire new_AGEMA_signal_18286 ;
    wire new_AGEMA_signal_18287 ;
    wire new_AGEMA_signal_18288 ;
    wire new_AGEMA_signal_18289 ;
    wire new_AGEMA_signal_18290 ;
    wire new_AGEMA_signal_18291 ;
    wire new_AGEMA_signal_18292 ;
    wire new_AGEMA_signal_18293 ;
    wire new_AGEMA_signal_18294 ;
    wire new_AGEMA_signal_18295 ;
    wire new_AGEMA_signal_18296 ;
    wire new_AGEMA_signal_18297 ;
    wire new_AGEMA_signal_18298 ;
    wire new_AGEMA_signal_18299 ;
    wire new_AGEMA_signal_18300 ;
    wire new_AGEMA_signal_18301 ;
    wire new_AGEMA_signal_18302 ;
    wire new_AGEMA_signal_18303 ;
    wire new_AGEMA_signal_18304 ;
    wire new_AGEMA_signal_18305 ;
    wire new_AGEMA_signal_18306 ;
    wire new_AGEMA_signal_18307 ;
    wire new_AGEMA_signal_18308 ;
    wire new_AGEMA_signal_18309 ;
    wire new_AGEMA_signal_18310 ;
    wire new_AGEMA_signal_18311 ;
    wire new_AGEMA_signal_18312 ;
    wire new_AGEMA_signal_18313 ;
    wire new_AGEMA_signal_18314 ;
    wire new_AGEMA_signal_18315 ;
    wire new_AGEMA_signal_18316 ;
    wire new_AGEMA_signal_18320 ;
    wire new_AGEMA_signal_18321 ;
    wire new_AGEMA_signal_18322 ;
    wire new_AGEMA_signal_18323 ;
    wire new_AGEMA_signal_18324 ;
    wire new_AGEMA_signal_18325 ;
    wire new_AGEMA_signal_18326 ;
    wire new_AGEMA_signal_18327 ;
    wire new_AGEMA_signal_18328 ;
    wire new_AGEMA_signal_18329 ;
    wire new_AGEMA_signal_18330 ;
    wire new_AGEMA_signal_18331 ;
    wire new_AGEMA_signal_18332 ;
    wire new_AGEMA_signal_18333 ;
    wire new_AGEMA_signal_18334 ;
    wire new_AGEMA_signal_18335 ;
    wire new_AGEMA_signal_18336 ;
    wire new_AGEMA_signal_18337 ;
    wire new_AGEMA_signal_18338 ;
    wire new_AGEMA_signal_18339 ;
    wire new_AGEMA_signal_18340 ;
    wire new_AGEMA_signal_18341 ;
    wire new_AGEMA_signal_18342 ;
    wire new_AGEMA_signal_18343 ;
    wire new_AGEMA_signal_18344 ;
    wire new_AGEMA_signal_18345 ;
    wire new_AGEMA_signal_18346 ;
    wire new_AGEMA_signal_18347 ;
    wire new_AGEMA_signal_18348 ;
    wire new_AGEMA_signal_18349 ;
    wire new_AGEMA_signal_18350 ;
    wire new_AGEMA_signal_18351 ;
    wire new_AGEMA_signal_18352 ;
    wire new_AGEMA_signal_18353 ;
    wire new_AGEMA_signal_18354 ;
    wire new_AGEMA_signal_18355 ;
    wire new_AGEMA_signal_18356 ;
    wire new_AGEMA_signal_18357 ;
    wire new_AGEMA_signal_18358 ;
    wire new_AGEMA_signal_18359 ;
    wire new_AGEMA_signal_18360 ;
    wire new_AGEMA_signal_18361 ;
    wire new_AGEMA_signal_18362 ;
    wire new_AGEMA_signal_18363 ;
    wire new_AGEMA_signal_18364 ;
    wire new_AGEMA_signal_18365 ;
    wire new_AGEMA_signal_18366 ;
    wire new_AGEMA_signal_18367 ;
    wire new_AGEMA_signal_18368 ;
    wire new_AGEMA_signal_18369 ;
    wire new_AGEMA_signal_18370 ;
    wire new_AGEMA_signal_18371 ;
    wire new_AGEMA_signal_18372 ;
    wire new_AGEMA_signal_18373 ;
    wire new_AGEMA_signal_18374 ;
    wire new_AGEMA_signal_18375 ;
    wire new_AGEMA_signal_18376 ;
    wire new_AGEMA_signal_18377 ;
    wire new_AGEMA_signal_18378 ;
    wire new_AGEMA_signal_18379 ;
    wire new_AGEMA_signal_18380 ;
    wire new_AGEMA_signal_18381 ;
    wire new_AGEMA_signal_18382 ;
    wire new_AGEMA_signal_18383 ;
    wire new_AGEMA_signal_18384 ;
    wire new_AGEMA_signal_18385 ;
    wire new_AGEMA_signal_18386 ;
    wire new_AGEMA_signal_18387 ;
    wire new_AGEMA_signal_18388 ;
    wire new_AGEMA_signal_18389 ;
    wire new_AGEMA_signal_18390 ;
    wire new_AGEMA_signal_18391 ;
    wire new_AGEMA_signal_18392 ;
    wire new_AGEMA_signal_18393 ;
    wire new_AGEMA_signal_18394 ;
    wire new_AGEMA_signal_18395 ;
    wire new_AGEMA_signal_18396 ;
    wire new_AGEMA_signal_18397 ;
    wire new_AGEMA_signal_18398 ;
    wire new_AGEMA_signal_18399 ;
    wire new_AGEMA_signal_18400 ;
    wire new_AGEMA_signal_18401 ;
    wire new_AGEMA_signal_18402 ;
    wire new_AGEMA_signal_18403 ;
    wire new_AGEMA_signal_18404 ;
    wire new_AGEMA_signal_18405 ;
    wire new_AGEMA_signal_18406 ;
    wire new_AGEMA_signal_18407 ;
    wire new_AGEMA_signal_18408 ;
    wire new_AGEMA_signal_18409 ;
    wire new_AGEMA_signal_18410 ;
    wire new_AGEMA_signal_18411 ;
    wire new_AGEMA_signal_18412 ;
    wire new_AGEMA_signal_18416 ;
    wire new_AGEMA_signal_18417 ;
    wire new_AGEMA_signal_18418 ;
    wire new_AGEMA_signal_18419 ;
    wire new_AGEMA_signal_18420 ;
    wire new_AGEMA_signal_18421 ;
    wire new_AGEMA_signal_18422 ;
    wire new_AGEMA_signal_18423 ;
    wire new_AGEMA_signal_18424 ;
    wire new_AGEMA_signal_18425 ;
    wire new_AGEMA_signal_18426 ;
    wire new_AGEMA_signal_18427 ;
    wire new_AGEMA_signal_18428 ;
    wire new_AGEMA_signal_18429 ;
    wire new_AGEMA_signal_18430 ;
    wire new_AGEMA_signal_18431 ;
    wire new_AGEMA_signal_18432 ;
    wire new_AGEMA_signal_18433 ;
    wire new_AGEMA_signal_18434 ;
    wire new_AGEMA_signal_18435 ;
    wire new_AGEMA_signal_18436 ;
    wire new_AGEMA_signal_18437 ;
    wire new_AGEMA_signal_18438 ;
    wire new_AGEMA_signal_18439 ;
    wire new_AGEMA_signal_18440 ;
    wire new_AGEMA_signal_18441 ;
    wire new_AGEMA_signal_18442 ;
    wire new_AGEMA_signal_18443 ;
    wire new_AGEMA_signal_18444 ;
    wire new_AGEMA_signal_18445 ;
    wire new_AGEMA_signal_18446 ;
    wire new_AGEMA_signal_18447 ;
    wire new_AGEMA_signal_18448 ;
    wire new_AGEMA_signal_18449 ;
    wire new_AGEMA_signal_18450 ;
    wire new_AGEMA_signal_18451 ;
    wire new_AGEMA_signal_18452 ;
    wire new_AGEMA_signal_18453 ;
    wire new_AGEMA_signal_18454 ;
    wire new_AGEMA_signal_18455 ;
    wire new_AGEMA_signal_18456 ;
    wire new_AGEMA_signal_18457 ;
    wire new_AGEMA_signal_18458 ;
    wire new_AGEMA_signal_18459 ;
    wire new_AGEMA_signal_18460 ;
    wire new_AGEMA_signal_18461 ;
    wire new_AGEMA_signal_18462 ;
    wire new_AGEMA_signal_18463 ;
    wire new_AGEMA_signal_18464 ;
    wire new_AGEMA_signal_18465 ;
    wire new_AGEMA_signal_18466 ;
    wire new_AGEMA_signal_18467 ;
    wire new_AGEMA_signal_18468 ;
    wire new_AGEMA_signal_18469 ;
    wire new_AGEMA_signal_18470 ;
    wire new_AGEMA_signal_18471 ;
    wire new_AGEMA_signal_18472 ;
    wire new_AGEMA_signal_18473 ;
    wire new_AGEMA_signal_18474 ;
    wire new_AGEMA_signal_18475 ;
    wire new_AGEMA_signal_18476 ;
    wire new_AGEMA_signal_18477 ;
    wire new_AGEMA_signal_18478 ;
    wire new_AGEMA_signal_18479 ;
    wire new_AGEMA_signal_18480 ;
    wire new_AGEMA_signal_18481 ;
    wire new_AGEMA_signal_18482 ;
    wire new_AGEMA_signal_18483 ;
    wire new_AGEMA_signal_18484 ;
    wire new_AGEMA_signal_18485 ;
    wire new_AGEMA_signal_18486 ;
    wire new_AGEMA_signal_18487 ;
    wire new_AGEMA_signal_18488 ;
    wire new_AGEMA_signal_18489 ;
    wire new_AGEMA_signal_18490 ;
    wire new_AGEMA_signal_18491 ;
    wire new_AGEMA_signal_18492 ;
    wire new_AGEMA_signal_18493 ;
    wire new_AGEMA_signal_18494 ;
    wire new_AGEMA_signal_18495 ;
    wire new_AGEMA_signal_18496 ;
    wire new_AGEMA_signal_18497 ;
    wire new_AGEMA_signal_18498 ;
    wire new_AGEMA_signal_18499 ;
    wire new_AGEMA_signal_18500 ;
    wire new_AGEMA_signal_18501 ;
    wire new_AGEMA_signal_18502 ;
    wire new_AGEMA_signal_18503 ;
    wire new_AGEMA_signal_18504 ;
    wire new_AGEMA_signal_18505 ;
    wire new_AGEMA_signal_18506 ;
    wire new_AGEMA_signal_18507 ;
    wire new_AGEMA_signal_18508 ;
    wire new_AGEMA_signal_18509 ;
    wire new_AGEMA_signal_18510 ;
    wire new_AGEMA_signal_18511 ;
    wire new_AGEMA_signal_18512 ;
    wire new_AGEMA_signal_18513 ;
    wire new_AGEMA_signal_18514 ;
    wire new_AGEMA_signal_18515 ;
    wire new_AGEMA_signal_18516 ;
    wire new_AGEMA_signal_18517 ;
    wire new_AGEMA_signal_18518 ;
    wire new_AGEMA_signal_18519 ;
    wire new_AGEMA_signal_18520 ;
    wire new_AGEMA_signal_18521 ;
    wire new_AGEMA_signal_18522 ;
    wire new_AGEMA_signal_18523 ;
    wire new_AGEMA_signal_18524 ;
    wire new_AGEMA_signal_18525 ;
    wire new_AGEMA_signal_18526 ;
    wire new_AGEMA_signal_18527 ;
    wire new_AGEMA_signal_18528 ;
    wire new_AGEMA_signal_18529 ;
    wire new_AGEMA_signal_18530 ;
    wire new_AGEMA_signal_18531 ;
    wire new_AGEMA_signal_18532 ;
    wire new_AGEMA_signal_18533 ;
    wire new_AGEMA_signal_18534 ;
    wire new_AGEMA_signal_18535 ;
    wire new_AGEMA_signal_18536 ;
    wire new_AGEMA_signal_18537 ;
    wire new_AGEMA_signal_18538 ;
    wire new_AGEMA_signal_18539 ;
    wire new_AGEMA_signal_18540 ;
    wire new_AGEMA_signal_18541 ;
    wire new_AGEMA_signal_18545 ;
    wire new_AGEMA_signal_18546 ;
    wire new_AGEMA_signal_18547 ;
    wire new_AGEMA_signal_18548 ;
    wire new_AGEMA_signal_18549 ;
    wire new_AGEMA_signal_18550 ;
    wire new_AGEMA_signal_18551 ;
    wire new_AGEMA_signal_18552 ;
    wire new_AGEMA_signal_18553 ;
    wire new_AGEMA_signal_18554 ;
    wire new_AGEMA_signal_18555 ;
    wire new_AGEMA_signal_18556 ;
    wire new_AGEMA_signal_18557 ;
    wire new_AGEMA_signal_18558 ;
    wire new_AGEMA_signal_18559 ;
    wire new_AGEMA_signal_18560 ;
    wire new_AGEMA_signal_18561 ;
    wire new_AGEMA_signal_18562 ;
    wire new_AGEMA_signal_18563 ;
    wire new_AGEMA_signal_18564 ;
    wire new_AGEMA_signal_18565 ;
    wire new_AGEMA_signal_18566 ;
    wire new_AGEMA_signal_18567 ;
    wire new_AGEMA_signal_18568 ;
    wire new_AGEMA_signal_18569 ;
    wire new_AGEMA_signal_18570 ;
    wire new_AGEMA_signal_18571 ;
    wire new_AGEMA_signal_18572 ;
    wire new_AGEMA_signal_18573 ;
    wire new_AGEMA_signal_18574 ;
    wire new_AGEMA_signal_18575 ;
    wire new_AGEMA_signal_18576 ;
    wire new_AGEMA_signal_18577 ;
    wire new_AGEMA_signal_18578 ;
    wire new_AGEMA_signal_18579 ;
    wire new_AGEMA_signal_18580 ;
    wire new_AGEMA_signal_18581 ;
    wire new_AGEMA_signal_18582 ;
    wire new_AGEMA_signal_18583 ;
    wire new_AGEMA_signal_18584 ;
    wire new_AGEMA_signal_18585 ;
    wire new_AGEMA_signal_18586 ;
    wire new_AGEMA_signal_18587 ;
    wire new_AGEMA_signal_18588 ;
    wire new_AGEMA_signal_18589 ;
    wire new_AGEMA_signal_18590 ;
    wire new_AGEMA_signal_18591 ;
    wire new_AGEMA_signal_18592 ;
    wire new_AGEMA_signal_18593 ;
    wire new_AGEMA_signal_18594 ;
    wire new_AGEMA_signal_18595 ;
    wire new_AGEMA_signal_18599 ;
    wire new_AGEMA_signal_18600 ;
    wire new_AGEMA_signal_18601 ;
    wire new_AGEMA_signal_18602 ;
    wire new_AGEMA_signal_18603 ;
    wire new_AGEMA_signal_18604 ;
    wire new_AGEMA_signal_18605 ;
    wire new_AGEMA_signal_18606 ;
    wire new_AGEMA_signal_18607 ;
    wire new_AGEMA_signal_18608 ;
    wire new_AGEMA_signal_18609 ;
    wire new_AGEMA_signal_18610 ;
    wire new_AGEMA_signal_18611 ;
    wire new_AGEMA_signal_18612 ;
    wire new_AGEMA_signal_18613 ;
    wire new_AGEMA_signal_18614 ;
    wire new_AGEMA_signal_18615 ;
    wire new_AGEMA_signal_18616 ;
    wire new_AGEMA_signal_18617 ;
    wire new_AGEMA_signal_18618 ;
    wire new_AGEMA_signal_18619 ;
    wire new_AGEMA_signal_18620 ;
    wire new_AGEMA_signal_18621 ;
    wire new_AGEMA_signal_18622 ;
    wire new_AGEMA_signal_18623 ;
    wire new_AGEMA_signal_18624 ;
    wire new_AGEMA_signal_18625 ;
    wire new_AGEMA_signal_18626 ;
    wire new_AGEMA_signal_18627 ;
    wire new_AGEMA_signal_18628 ;
    wire new_AGEMA_signal_18629 ;
    wire new_AGEMA_signal_18630 ;
    wire new_AGEMA_signal_18631 ;
    wire new_AGEMA_signal_18632 ;
    wire new_AGEMA_signal_18633 ;
    wire new_AGEMA_signal_18634 ;
    wire new_AGEMA_signal_18635 ;
    wire new_AGEMA_signal_18636 ;
    wire new_AGEMA_signal_18637 ;
    wire new_AGEMA_signal_18638 ;
    wire new_AGEMA_signal_18639 ;
    wire new_AGEMA_signal_18640 ;
    wire new_AGEMA_signal_18641 ;
    wire new_AGEMA_signal_18642 ;
    wire new_AGEMA_signal_18643 ;
    wire new_AGEMA_signal_18644 ;
    wire new_AGEMA_signal_18645 ;
    wire new_AGEMA_signal_18646 ;
    wire new_AGEMA_signal_18647 ;
    wire new_AGEMA_signal_18648 ;
    wire new_AGEMA_signal_18649 ;
    wire new_AGEMA_signal_18650 ;
    wire new_AGEMA_signal_18651 ;
    wire new_AGEMA_signal_18652 ;
    wire new_AGEMA_signal_18653 ;
    wire new_AGEMA_signal_18654 ;
    wire new_AGEMA_signal_18655 ;
    wire new_AGEMA_signal_18656 ;
    wire new_AGEMA_signal_18657 ;
    wire new_AGEMA_signal_18658 ;
    wire new_AGEMA_signal_18659 ;
    wire new_AGEMA_signal_18660 ;
    wire new_AGEMA_signal_18661 ;
    wire new_AGEMA_signal_18662 ;
    wire new_AGEMA_signal_18663 ;
    wire new_AGEMA_signal_18664 ;
    wire new_AGEMA_signal_18665 ;
    wire new_AGEMA_signal_18666 ;
    wire new_AGEMA_signal_18667 ;
    wire new_AGEMA_signal_18668 ;
    wire new_AGEMA_signal_18669 ;
    wire new_AGEMA_signal_18670 ;
    wire new_AGEMA_signal_18671 ;
    wire new_AGEMA_signal_18672 ;
    wire new_AGEMA_signal_18673 ;
    wire new_AGEMA_signal_18674 ;
    wire new_AGEMA_signal_18675 ;
    wire new_AGEMA_signal_18676 ;
    wire new_AGEMA_signal_18677 ;
    wire new_AGEMA_signal_18678 ;
    wire new_AGEMA_signal_18679 ;
    wire new_AGEMA_signal_18680 ;
    wire new_AGEMA_signal_18681 ;
    wire new_AGEMA_signal_18682 ;
    wire new_AGEMA_signal_18683 ;
    wire new_AGEMA_signal_18684 ;
    wire new_AGEMA_signal_18685 ;
    wire new_AGEMA_signal_18686 ;
    wire new_AGEMA_signal_18687 ;
    wire new_AGEMA_signal_18688 ;
    wire new_AGEMA_signal_18689 ;
    wire new_AGEMA_signal_18690 ;
    wire new_AGEMA_signal_18691 ;
    wire new_AGEMA_signal_18692 ;
    wire new_AGEMA_signal_18693 ;
    wire new_AGEMA_signal_18694 ;
    wire new_AGEMA_signal_18695 ;
    wire new_AGEMA_signal_18696 ;
    wire new_AGEMA_signal_18697 ;
    wire new_AGEMA_signal_18698 ;
    wire new_AGEMA_signal_18699 ;
    wire new_AGEMA_signal_18700 ;
    wire new_AGEMA_signal_18701 ;
    wire new_AGEMA_signal_18702 ;
    wire new_AGEMA_signal_18703 ;
    wire new_AGEMA_signal_18704 ;
    wire new_AGEMA_signal_18705 ;
    wire new_AGEMA_signal_18706 ;
    wire new_AGEMA_signal_18707 ;
    wire new_AGEMA_signal_18708 ;
    wire new_AGEMA_signal_18709 ;
    wire new_AGEMA_signal_18749 ;
    wire new_AGEMA_signal_18750 ;
    wire new_AGEMA_signal_18751 ;
    wire new_AGEMA_signal_18752 ;
    wire new_AGEMA_signal_18753 ;
    wire new_AGEMA_signal_18754 ;
    wire new_AGEMA_signal_18755 ;
    wire new_AGEMA_signal_18756 ;
    wire new_AGEMA_signal_18757 ;
    wire new_AGEMA_signal_18758 ;
    wire new_AGEMA_signal_18759 ;
    wire new_AGEMA_signal_18760 ;
    wire new_AGEMA_signal_18761 ;
    wire new_AGEMA_signal_18762 ;
    wire new_AGEMA_signal_18763 ;
    wire new_AGEMA_signal_18764 ;
    wire new_AGEMA_signal_18765 ;
    wire new_AGEMA_signal_18766 ;
    wire new_AGEMA_signal_18767 ;
    wire new_AGEMA_signal_18768 ;
    wire new_AGEMA_signal_18769 ;
    wire new_AGEMA_signal_18770 ;
    wire new_AGEMA_signal_18771 ;
    wire new_AGEMA_signal_18772 ;
    wire new_AGEMA_signal_18773 ;
    wire new_AGEMA_signal_18774 ;
    wire new_AGEMA_signal_18775 ;
    wire new_AGEMA_signal_18776 ;
    wire new_AGEMA_signal_18777 ;
    wire new_AGEMA_signal_18778 ;
    wire new_AGEMA_signal_18779 ;
    wire new_AGEMA_signal_18780 ;
    wire new_AGEMA_signal_18781 ;
    wire new_AGEMA_signal_18782 ;
    wire new_AGEMA_signal_18783 ;
    wire new_AGEMA_signal_18784 ;
    wire new_AGEMA_signal_18785 ;
    wire new_AGEMA_signal_18786 ;
    wire new_AGEMA_signal_18787 ;
    wire new_AGEMA_signal_18788 ;
    wire new_AGEMA_signal_18789 ;
    wire new_AGEMA_signal_18790 ;
    wire new_AGEMA_signal_18791 ;
    wire new_AGEMA_signal_18792 ;
    wire new_AGEMA_signal_18793 ;
    wire new_AGEMA_signal_18794 ;
    wire new_AGEMA_signal_18795 ;
    wire new_AGEMA_signal_18796 ;
    wire new_AGEMA_signal_18797 ;
    wire new_AGEMA_signal_18798 ;
    wire new_AGEMA_signal_18799 ;
    wire new_AGEMA_signal_18800 ;
    wire new_AGEMA_signal_18801 ;
    wire new_AGEMA_signal_18802 ;
    wire new_AGEMA_signal_18803 ;
    wire new_AGEMA_signal_18804 ;
    wire new_AGEMA_signal_18805 ;
    wire new_AGEMA_signal_18806 ;
    wire new_AGEMA_signal_18807 ;
    wire new_AGEMA_signal_18808 ;
    wire new_AGEMA_signal_18809 ;
    wire new_AGEMA_signal_18810 ;
    wire new_AGEMA_signal_18811 ;
    wire new_AGEMA_signal_18812 ;
    wire new_AGEMA_signal_18813 ;
    wire new_AGEMA_signal_18814 ;
    wire new_AGEMA_signal_18815 ;
    wire new_AGEMA_signal_18816 ;
    wire new_AGEMA_signal_18817 ;
    wire new_AGEMA_signal_18818 ;
    wire new_AGEMA_signal_18819 ;
    wire new_AGEMA_signal_18820 ;
    wire new_AGEMA_signal_18821 ;
    wire new_AGEMA_signal_18822 ;
    wire new_AGEMA_signal_18823 ;
    wire new_AGEMA_signal_18824 ;
    wire new_AGEMA_signal_18825 ;
    wire new_AGEMA_signal_18826 ;
    wire new_AGEMA_signal_18827 ;
    wire new_AGEMA_signal_18828 ;
    wire new_AGEMA_signal_18829 ;
    wire new_AGEMA_signal_18830 ;
    wire new_AGEMA_signal_18831 ;
    wire new_AGEMA_signal_18832 ;
    wire new_AGEMA_signal_18833 ;
    wire new_AGEMA_signal_18834 ;
    wire new_AGEMA_signal_18835 ;
    wire new_AGEMA_signal_18836 ;
    wire new_AGEMA_signal_18837 ;
    wire new_AGEMA_signal_18838 ;
    wire new_AGEMA_signal_18839 ;
    wire new_AGEMA_signal_18840 ;
    wire new_AGEMA_signal_18841 ;
    wire new_AGEMA_signal_18842 ;
    wire new_AGEMA_signal_18843 ;
    wire new_AGEMA_signal_18844 ;
    wire new_AGEMA_signal_18848 ;
    wire new_AGEMA_signal_18849 ;
    wire new_AGEMA_signal_18850 ;
    wire new_AGEMA_signal_18851 ;
    wire new_AGEMA_signal_18852 ;
    wire new_AGEMA_signal_18853 ;
    wire new_AGEMA_signal_18854 ;
    wire new_AGEMA_signal_18855 ;
    wire new_AGEMA_signal_18856 ;
    wire new_AGEMA_signal_18857 ;
    wire new_AGEMA_signal_18858 ;
    wire new_AGEMA_signal_18859 ;
    wire new_AGEMA_signal_18860 ;
    wire new_AGEMA_signal_18861 ;
    wire new_AGEMA_signal_18862 ;
    wire new_AGEMA_signal_18863 ;
    wire new_AGEMA_signal_18864 ;
    wire new_AGEMA_signal_18865 ;
    wire new_AGEMA_signal_18866 ;
    wire new_AGEMA_signal_18867 ;
    wire new_AGEMA_signal_18868 ;
    wire new_AGEMA_signal_18869 ;
    wire new_AGEMA_signal_18870 ;
    wire new_AGEMA_signal_18871 ;
    wire new_AGEMA_signal_18872 ;
    wire new_AGEMA_signal_18873 ;
    wire new_AGEMA_signal_18874 ;
    wire new_AGEMA_signal_18875 ;
    wire new_AGEMA_signal_18876 ;
    wire new_AGEMA_signal_18877 ;
    wire new_AGEMA_signal_18878 ;
    wire new_AGEMA_signal_18879 ;
    wire new_AGEMA_signal_18880 ;
    wire new_AGEMA_signal_18881 ;
    wire new_AGEMA_signal_18882 ;
    wire new_AGEMA_signal_18883 ;
    wire new_AGEMA_signal_18884 ;
    wire new_AGEMA_signal_18885 ;
    wire new_AGEMA_signal_18886 ;
    wire new_AGEMA_signal_18887 ;
    wire new_AGEMA_signal_18888 ;
    wire new_AGEMA_signal_18889 ;
    wire new_AGEMA_signal_18890 ;
    wire new_AGEMA_signal_18891 ;
    wire new_AGEMA_signal_18892 ;
    wire new_AGEMA_signal_18893 ;
    wire new_AGEMA_signal_18894 ;
    wire new_AGEMA_signal_18895 ;
    wire new_AGEMA_signal_18896 ;
    wire new_AGEMA_signal_18897 ;
    wire new_AGEMA_signal_18898 ;
    wire new_AGEMA_signal_18899 ;
    wire new_AGEMA_signal_18900 ;
    wire new_AGEMA_signal_18901 ;
    wire new_AGEMA_signal_18902 ;
    wire new_AGEMA_signal_18903 ;
    wire new_AGEMA_signal_18904 ;
    wire new_AGEMA_signal_18905 ;
    wire new_AGEMA_signal_18906 ;
    wire new_AGEMA_signal_18907 ;
    wire new_AGEMA_signal_18908 ;
    wire new_AGEMA_signal_18909 ;
    wire new_AGEMA_signal_18910 ;
    wire new_AGEMA_signal_18911 ;
    wire new_AGEMA_signal_18912 ;
    wire new_AGEMA_signal_18913 ;
    wire new_AGEMA_signal_18917 ;
    wire new_AGEMA_signal_18918 ;
    wire new_AGEMA_signal_18919 ;
    wire new_AGEMA_signal_18920 ;
    wire new_AGEMA_signal_18921 ;
    wire new_AGEMA_signal_18922 ;
    wire new_AGEMA_signal_18923 ;
    wire new_AGEMA_signal_18924 ;
    wire new_AGEMA_signal_18925 ;
    wire new_AGEMA_signal_18926 ;
    wire new_AGEMA_signal_18927 ;
    wire new_AGEMA_signal_18928 ;
    wire new_AGEMA_signal_18929 ;
    wire new_AGEMA_signal_18930 ;
    wire new_AGEMA_signal_18931 ;
    wire new_AGEMA_signal_18932 ;
    wire new_AGEMA_signal_18933 ;
    wire new_AGEMA_signal_18934 ;
    wire new_AGEMA_signal_18935 ;
    wire new_AGEMA_signal_18936 ;
    wire new_AGEMA_signal_18937 ;
    wire new_AGEMA_signal_18938 ;
    wire new_AGEMA_signal_18939 ;
    wire new_AGEMA_signal_18940 ;
    wire new_AGEMA_signal_18941 ;
    wire new_AGEMA_signal_18942 ;
    wire new_AGEMA_signal_18943 ;
    wire new_AGEMA_signal_18944 ;
    wire new_AGEMA_signal_18945 ;
    wire new_AGEMA_signal_18946 ;
    wire new_AGEMA_signal_18947 ;
    wire new_AGEMA_signal_18948 ;
    wire new_AGEMA_signal_18949 ;
    wire new_AGEMA_signal_18950 ;
    wire new_AGEMA_signal_18951 ;
    wire new_AGEMA_signal_18952 ;
    wire new_AGEMA_signal_18953 ;
    wire new_AGEMA_signal_18954 ;
    wire new_AGEMA_signal_18955 ;
    wire new_AGEMA_signal_18956 ;
    wire new_AGEMA_signal_18957 ;
    wire new_AGEMA_signal_18958 ;
    wire new_AGEMA_signal_18959 ;
    wire new_AGEMA_signal_18960 ;
    wire new_AGEMA_signal_18961 ;
    wire new_AGEMA_signal_18962 ;
    wire new_AGEMA_signal_18963 ;
    wire new_AGEMA_signal_18964 ;
    wire new_AGEMA_signal_18965 ;
    wire new_AGEMA_signal_18966 ;
    wire new_AGEMA_signal_18967 ;
    wire new_AGEMA_signal_18968 ;
    wire new_AGEMA_signal_18969 ;
    wire new_AGEMA_signal_18970 ;
    wire new_AGEMA_signal_18971 ;
    wire new_AGEMA_signal_18972 ;
    wire new_AGEMA_signal_18973 ;
    wire new_AGEMA_signal_18974 ;
    wire new_AGEMA_signal_18975 ;
    wire new_AGEMA_signal_18976 ;
    wire new_AGEMA_signal_18977 ;
    wire new_AGEMA_signal_18978 ;
    wire new_AGEMA_signal_18979 ;
    wire new_AGEMA_signal_18980 ;
    wire new_AGEMA_signal_18981 ;
    wire new_AGEMA_signal_18982 ;
    wire new_AGEMA_signal_18983 ;
    wire new_AGEMA_signal_18984 ;
    wire new_AGEMA_signal_18985 ;
    wire new_AGEMA_signal_18989 ;
    wire new_AGEMA_signal_18990 ;
    wire new_AGEMA_signal_18991 ;
    wire new_AGEMA_signal_18992 ;
    wire new_AGEMA_signal_18993 ;
    wire new_AGEMA_signal_18994 ;
    wire new_AGEMA_signal_18995 ;
    wire new_AGEMA_signal_18996 ;
    wire new_AGEMA_signal_18997 ;
    wire new_AGEMA_signal_18998 ;
    wire new_AGEMA_signal_18999 ;
    wire new_AGEMA_signal_19000 ;
    wire new_AGEMA_signal_19001 ;
    wire new_AGEMA_signal_19002 ;
    wire new_AGEMA_signal_19003 ;
    wire new_AGEMA_signal_19004 ;
    wire new_AGEMA_signal_19005 ;
    wire new_AGEMA_signal_19006 ;
    wire new_AGEMA_signal_19007 ;
    wire new_AGEMA_signal_19008 ;
    wire new_AGEMA_signal_19009 ;
    wire new_AGEMA_signal_19010 ;
    wire new_AGEMA_signal_19011 ;
    wire new_AGEMA_signal_19012 ;
    wire new_AGEMA_signal_19013 ;
    wire new_AGEMA_signal_19014 ;
    wire new_AGEMA_signal_19015 ;
    wire new_AGEMA_signal_19016 ;
    wire new_AGEMA_signal_19017 ;
    wire new_AGEMA_signal_19018 ;
    wire new_AGEMA_signal_19019 ;
    wire new_AGEMA_signal_19020 ;
    wire new_AGEMA_signal_19021 ;
    wire new_AGEMA_signal_19022 ;
    wire new_AGEMA_signal_19023 ;
    wire new_AGEMA_signal_19024 ;
    wire new_AGEMA_signal_19025 ;
    wire new_AGEMA_signal_19026 ;
    wire new_AGEMA_signal_19027 ;
    wire new_AGEMA_signal_19028 ;
    wire new_AGEMA_signal_19029 ;
    wire new_AGEMA_signal_19030 ;
    wire new_AGEMA_signal_19031 ;
    wire new_AGEMA_signal_19032 ;
    wire new_AGEMA_signal_19033 ;
    wire new_AGEMA_signal_19034 ;
    wire new_AGEMA_signal_19035 ;
    wire new_AGEMA_signal_19036 ;
    wire new_AGEMA_signal_19037 ;
    wire new_AGEMA_signal_19038 ;
    wire new_AGEMA_signal_19039 ;
    wire new_AGEMA_signal_19040 ;
    wire new_AGEMA_signal_19041 ;
    wire new_AGEMA_signal_19042 ;
    wire new_AGEMA_signal_19046 ;
    wire new_AGEMA_signal_19047 ;
    wire new_AGEMA_signal_19048 ;
    wire new_AGEMA_signal_19049 ;
    wire new_AGEMA_signal_19050 ;
    wire new_AGEMA_signal_19051 ;
    wire new_AGEMA_signal_19052 ;
    wire new_AGEMA_signal_19053 ;
    wire new_AGEMA_signal_19054 ;
    wire new_AGEMA_signal_19055 ;
    wire new_AGEMA_signal_19056 ;
    wire new_AGEMA_signal_19057 ;
    wire new_AGEMA_signal_19058 ;
    wire new_AGEMA_signal_19059 ;
    wire new_AGEMA_signal_19060 ;
    wire new_AGEMA_signal_19061 ;
    wire new_AGEMA_signal_19062 ;
    wire new_AGEMA_signal_19063 ;
    wire new_AGEMA_signal_19064 ;
    wire new_AGEMA_signal_19065 ;
    wire new_AGEMA_signal_19066 ;
    wire new_AGEMA_signal_19067 ;
    wire new_AGEMA_signal_19068 ;
    wire new_AGEMA_signal_19069 ;
    wire new_AGEMA_signal_19070 ;
    wire new_AGEMA_signal_19071 ;
    wire new_AGEMA_signal_19072 ;
    wire new_AGEMA_signal_19073 ;
    wire new_AGEMA_signal_19074 ;
    wire new_AGEMA_signal_19075 ;
    wire new_AGEMA_signal_19076 ;
    wire new_AGEMA_signal_19077 ;
    wire new_AGEMA_signal_19078 ;
    wire new_AGEMA_signal_19079 ;
    wire new_AGEMA_signal_19080 ;
    wire new_AGEMA_signal_19081 ;
    wire new_AGEMA_signal_19082 ;
    wire new_AGEMA_signal_19083 ;
    wire new_AGEMA_signal_19084 ;
    wire new_AGEMA_signal_19085 ;
    wire new_AGEMA_signal_19086 ;
    wire new_AGEMA_signal_19087 ;
    wire new_AGEMA_signal_19088 ;
    wire new_AGEMA_signal_19089 ;
    wire new_AGEMA_signal_19090 ;
    wire new_AGEMA_signal_19091 ;
    wire new_AGEMA_signal_19092 ;
    wire new_AGEMA_signal_19093 ;
    wire new_AGEMA_signal_19094 ;
    wire new_AGEMA_signal_19095 ;
    wire new_AGEMA_signal_19096 ;
    wire new_AGEMA_signal_19097 ;
    wire new_AGEMA_signal_19098 ;
    wire new_AGEMA_signal_19099 ;
    wire new_AGEMA_signal_19100 ;
    wire new_AGEMA_signal_19101 ;
    wire new_AGEMA_signal_19102 ;
    wire new_AGEMA_signal_19103 ;
    wire new_AGEMA_signal_19104 ;
    wire new_AGEMA_signal_19105 ;
    wire new_AGEMA_signal_19106 ;
    wire new_AGEMA_signal_19107 ;
    wire new_AGEMA_signal_19108 ;
    wire new_AGEMA_signal_19109 ;
    wire new_AGEMA_signal_19110 ;
    wire new_AGEMA_signal_19111 ;
    wire new_AGEMA_signal_19112 ;
    wire new_AGEMA_signal_19113 ;
    wire new_AGEMA_signal_19114 ;
    wire new_AGEMA_signal_19115 ;
    wire new_AGEMA_signal_19116 ;
    wire new_AGEMA_signal_19117 ;
    wire new_AGEMA_signal_19118 ;
    wire new_AGEMA_signal_19119 ;
    wire new_AGEMA_signal_19120 ;
    wire new_AGEMA_signal_19121 ;
    wire new_AGEMA_signal_19122 ;
    wire new_AGEMA_signal_19123 ;
    wire new_AGEMA_signal_19124 ;
    wire new_AGEMA_signal_19125 ;
    wire new_AGEMA_signal_19126 ;
    wire new_AGEMA_signal_19127 ;
    wire new_AGEMA_signal_19128 ;
    wire new_AGEMA_signal_19129 ;
    wire new_AGEMA_signal_19130 ;
    wire new_AGEMA_signal_19131 ;
    wire new_AGEMA_signal_19132 ;
    wire new_AGEMA_signal_19133 ;
    wire new_AGEMA_signal_19134 ;
    wire new_AGEMA_signal_19135 ;
    wire new_AGEMA_signal_19136 ;
    wire new_AGEMA_signal_19137 ;
    wire new_AGEMA_signal_19138 ;
    wire new_AGEMA_signal_19139 ;
    wire new_AGEMA_signal_19140 ;
    wire new_AGEMA_signal_19141 ;
    wire new_AGEMA_signal_19145 ;
    wire new_AGEMA_signal_19146 ;
    wire new_AGEMA_signal_19147 ;
    wire new_AGEMA_signal_19148 ;
    wire new_AGEMA_signal_19149 ;
    wire new_AGEMA_signal_19150 ;
    wire new_AGEMA_signal_19151 ;
    wire new_AGEMA_signal_19152 ;
    wire new_AGEMA_signal_19153 ;
    wire new_AGEMA_signal_19154 ;
    wire new_AGEMA_signal_19155 ;
    wire new_AGEMA_signal_19156 ;
    wire new_AGEMA_signal_19157 ;
    wire new_AGEMA_signal_19158 ;
    wire new_AGEMA_signal_19159 ;
    wire new_AGEMA_signal_19160 ;
    wire new_AGEMA_signal_19161 ;
    wire new_AGEMA_signal_19162 ;
    wire new_AGEMA_signal_19163 ;
    wire new_AGEMA_signal_19164 ;
    wire new_AGEMA_signal_19165 ;
    wire new_AGEMA_signal_19166 ;
    wire new_AGEMA_signal_19167 ;
    wire new_AGEMA_signal_19168 ;
    wire new_AGEMA_signal_19169 ;
    wire new_AGEMA_signal_19170 ;
    wire new_AGEMA_signal_19171 ;
    wire new_AGEMA_signal_19172 ;
    wire new_AGEMA_signal_19173 ;
    wire new_AGEMA_signal_19174 ;
    wire new_AGEMA_signal_19175 ;
    wire new_AGEMA_signal_19176 ;
    wire new_AGEMA_signal_19177 ;
    wire new_AGEMA_signal_19178 ;
    wire new_AGEMA_signal_19179 ;
    wire new_AGEMA_signal_19180 ;
    wire new_AGEMA_signal_19181 ;
    wire new_AGEMA_signal_19182 ;
    wire new_AGEMA_signal_19183 ;
    wire new_AGEMA_signal_19184 ;
    wire new_AGEMA_signal_19185 ;
    wire new_AGEMA_signal_19186 ;
    wire new_AGEMA_signal_19187 ;
    wire new_AGEMA_signal_19188 ;
    wire new_AGEMA_signal_19189 ;
    wire new_AGEMA_signal_19190 ;
    wire new_AGEMA_signal_19191 ;
    wire new_AGEMA_signal_19192 ;
    wire new_AGEMA_signal_19193 ;
    wire new_AGEMA_signal_19194 ;
    wire new_AGEMA_signal_19195 ;
    wire new_AGEMA_signal_19196 ;
    wire new_AGEMA_signal_19197 ;
    wire new_AGEMA_signal_19198 ;
    wire new_AGEMA_signal_19199 ;
    wire new_AGEMA_signal_19200 ;
    wire new_AGEMA_signal_19201 ;
    wire new_AGEMA_signal_19202 ;
    wire new_AGEMA_signal_19203 ;
    wire new_AGEMA_signal_19204 ;
    wire new_AGEMA_signal_19205 ;
    wire new_AGEMA_signal_19206 ;
    wire new_AGEMA_signal_19207 ;
    wire new_AGEMA_signal_19208 ;
    wire new_AGEMA_signal_19209 ;
    wire new_AGEMA_signal_19210 ;
    wire new_AGEMA_signal_19214 ;
    wire new_AGEMA_signal_19215 ;
    wire new_AGEMA_signal_19216 ;
    wire new_AGEMA_signal_19217 ;
    wire new_AGEMA_signal_19218 ;
    wire new_AGEMA_signal_19219 ;
    wire new_AGEMA_signal_19220 ;
    wire new_AGEMA_signal_19221 ;
    wire new_AGEMA_signal_19222 ;
    wire new_AGEMA_signal_19223 ;
    wire new_AGEMA_signal_19224 ;
    wire new_AGEMA_signal_19225 ;
    wire new_AGEMA_signal_19226 ;
    wire new_AGEMA_signal_19227 ;
    wire new_AGEMA_signal_19228 ;
    wire new_AGEMA_signal_19229 ;
    wire new_AGEMA_signal_19230 ;
    wire new_AGEMA_signal_19231 ;
    wire new_AGEMA_signal_19232 ;
    wire new_AGEMA_signal_19233 ;
    wire new_AGEMA_signal_19234 ;
    wire new_AGEMA_signal_19235 ;
    wire new_AGEMA_signal_19236 ;
    wire new_AGEMA_signal_19237 ;
    wire new_AGEMA_signal_19238 ;
    wire new_AGEMA_signal_19239 ;
    wire new_AGEMA_signal_19240 ;
    wire new_AGEMA_signal_19241 ;
    wire new_AGEMA_signal_19242 ;
    wire new_AGEMA_signal_19243 ;
    wire new_AGEMA_signal_19244 ;
    wire new_AGEMA_signal_19245 ;
    wire new_AGEMA_signal_19246 ;
    wire new_AGEMA_signal_19247 ;
    wire new_AGEMA_signal_19248 ;
    wire new_AGEMA_signal_19249 ;
    wire new_AGEMA_signal_19250 ;
    wire new_AGEMA_signal_19251 ;
    wire new_AGEMA_signal_19252 ;
    wire new_AGEMA_signal_19253 ;
    wire new_AGEMA_signal_19254 ;
    wire new_AGEMA_signal_19255 ;
    wire new_AGEMA_signal_19256 ;
    wire new_AGEMA_signal_19257 ;
    wire new_AGEMA_signal_19258 ;
    wire new_AGEMA_signal_19259 ;
    wire new_AGEMA_signal_19260 ;
    wire new_AGEMA_signal_19261 ;
    wire new_AGEMA_signal_19262 ;
    wire new_AGEMA_signal_19263 ;
    wire new_AGEMA_signal_19264 ;
    wire new_AGEMA_signal_19265 ;
    wire new_AGEMA_signal_19266 ;
    wire new_AGEMA_signal_19267 ;
    wire new_AGEMA_signal_19268 ;
    wire new_AGEMA_signal_19269 ;
    wire new_AGEMA_signal_19270 ;
    wire new_AGEMA_signal_19271 ;
    wire new_AGEMA_signal_19272 ;
    wire new_AGEMA_signal_19273 ;
    wire new_AGEMA_signal_19274 ;
    wire new_AGEMA_signal_19275 ;
    wire new_AGEMA_signal_19276 ;
    wire new_AGEMA_signal_19277 ;
    wire new_AGEMA_signal_19278 ;
    wire new_AGEMA_signal_19279 ;
    wire new_AGEMA_signal_19280 ;
    wire new_AGEMA_signal_19281 ;
    wire new_AGEMA_signal_19282 ;
    wire new_AGEMA_signal_19286 ;
    wire new_AGEMA_signal_19287 ;
    wire new_AGEMA_signal_19288 ;
    wire new_AGEMA_signal_19289 ;
    wire new_AGEMA_signal_19290 ;
    wire new_AGEMA_signal_19291 ;
    wire new_AGEMA_signal_19292 ;
    wire new_AGEMA_signal_19293 ;
    wire new_AGEMA_signal_19294 ;
    wire new_AGEMA_signal_19295 ;
    wire new_AGEMA_signal_19296 ;
    wire new_AGEMA_signal_19297 ;
    wire new_AGEMA_signal_19298 ;
    wire new_AGEMA_signal_19299 ;
    wire new_AGEMA_signal_19300 ;
    wire new_AGEMA_signal_19301 ;
    wire new_AGEMA_signal_19302 ;
    wire new_AGEMA_signal_19303 ;
    wire new_AGEMA_signal_19304 ;
    wire new_AGEMA_signal_19305 ;
    wire new_AGEMA_signal_19306 ;
    wire new_AGEMA_signal_19307 ;
    wire new_AGEMA_signal_19308 ;
    wire new_AGEMA_signal_19309 ;
    wire new_AGEMA_signal_19310 ;
    wire new_AGEMA_signal_19311 ;
    wire new_AGEMA_signal_19312 ;
    wire new_AGEMA_signal_19313 ;
    wire new_AGEMA_signal_19314 ;
    wire new_AGEMA_signal_19315 ;
    wire new_AGEMA_signal_19316 ;
    wire new_AGEMA_signal_19317 ;
    wire new_AGEMA_signal_19318 ;
    wire new_AGEMA_signal_19319 ;
    wire new_AGEMA_signal_19320 ;
    wire new_AGEMA_signal_19321 ;
    wire new_AGEMA_signal_19322 ;
    wire new_AGEMA_signal_19323 ;
    wire new_AGEMA_signal_19324 ;
    wire new_AGEMA_signal_19325 ;
    wire new_AGEMA_signal_19326 ;
    wire new_AGEMA_signal_19327 ;
    wire new_AGEMA_signal_19328 ;
    wire new_AGEMA_signal_19329 ;
    wire new_AGEMA_signal_19330 ;
    wire new_AGEMA_signal_19331 ;
    wire new_AGEMA_signal_19332 ;
    wire new_AGEMA_signal_19333 ;
    wire new_AGEMA_signal_19334 ;
    wire new_AGEMA_signal_19335 ;
    wire new_AGEMA_signal_19336 ;
    wire new_AGEMA_signal_19337 ;
    wire new_AGEMA_signal_19338 ;
    wire new_AGEMA_signal_19339 ;
    wire new_AGEMA_signal_19370 ;
    wire new_AGEMA_signal_19371 ;
    wire new_AGEMA_signal_19372 ;
    wire new_AGEMA_signal_19373 ;
    wire new_AGEMA_signal_19374 ;
    wire new_AGEMA_signal_19375 ;
    wire new_AGEMA_signal_19376 ;
    wire new_AGEMA_signal_19377 ;
    wire new_AGEMA_signal_19378 ;
    wire new_AGEMA_signal_19379 ;
    wire new_AGEMA_signal_19380 ;
    wire new_AGEMA_signal_19381 ;
    wire new_AGEMA_signal_19382 ;
    wire new_AGEMA_signal_19383 ;
    wire new_AGEMA_signal_19384 ;
    wire new_AGEMA_signal_19385 ;
    wire new_AGEMA_signal_19386 ;
    wire new_AGEMA_signal_19387 ;
    wire new_AGEMA_signal_19388 ;
    wire new_AGEMA_signal_19389 ;
    wire new_AGEMA_signal_19390 ;
    wire new_AGEMA_signal_19391 ;
    wire new_AGEMA_signal_19392 ;
    wire new_AGEMA_signal_19393 ;
    wire new_AGEMA_signal_19394 ;
    wire new_AGEMA_signal_19395 ;
    wire new_AGEMA_signal_19396 ;
    wire new_AGEMA_signal_19397 ;
    wire new_AGEMA_signal_19398 ;
    wire new_AGEMA_signal_19399 ;
    wire new_AGEMA_signal_19400 ;
    wire new_AGEMA_signal_19401 ;
    wire new_AGEMA_signal_19402 ;
    wire new_AGEMA_signal_19403 ;
    wire new_AGEMA_signal_19404 ;
    wire new_AGEMA_signal_19405 ;
    wire new_AGEMA_signal_19406 ;
    wire new_AGEMA_signal_19407 ;
    wire new_AGEMA_signal_19408 ;
    wire new_AGEMA_signal_19409 ;
    wire new_AGEMA_signal_19410 ;
    wire new_AGEMA_signal_19411 ;
    wire new_AGEMA_signal_19412 ;
    wire new_AGEMA_signal_19413 ;
    wire new_AGEMA_signal_19414 ;
    wire new_AGEMA_signal_19415 ;
    wire new_AGEMA_signal_19416 ;
    wire new_AGEMA_signal_19417 ;
    wire new_AGEMA_signal_19418 ;
    wire new_AGEMA_signal_19419 ;
    wire new_AGEMA_signal_19420 ;
    wire new_AGEMA_signal_19421 ;
    wire new_AGEMA_signal_19422 ;
    wire new_AGEMA_signal_19423 ;
    wire new_AGEMA_signal_19472 ;
    wire new_AGEMA_signal_19473 ;
    wire new_AGEMA_signal_19474 ;
    wire new_AGEMA_signal_19478 ;
    wire new_AGEMA_signal_19479 ;
    wire new_AGEMA_signal_19480 ;
    wire new_AGEMA_signal_19481 ;
    wire new_AGEMA_signal_19482 ;
    wire new_AGEMA_signal_19483 ;
    wire new_AGEMA_signal_19484 ;
    wire new_AGEMA_signal_19485 ;
    wire new_AGEMA_signal_19486 ;
    wire new_AGEMA_signal_19487 ;
    wire new_AGEMA_signal_19488 ;
    wire new_AGEMA_signal_19489 ;
    wire new_AGEMA_signal_19490 ;
    wire new_AGEMA_signal_19491 ;
    wire new_AGEMA_signal_19492 ;
    wire new_AGEMA_signal_19499 ;
    wire new_AGEMA_signal_19500 ;
    wire new_AGEMA_signal_19501 ;
    wire new_AGEMA_signal_19502 ;
    wire new_AGEMA_signal_19503 ;
    wire new_AGEMA_signal_19504 ;
    wire new_AGEMA_signal_19505 ;
    wire new_AGEMA_signal_19506 ;
    wire new_AGEMA_signal_19507 ;
    wire new_AGEMA_signal_19508 ;
    wire new_AGEMA_signal_19509 ;
    wire new_AGEMA_signal_19510 ;
    wire new_AGEMA_signal_19511 ;
    wire new_AGEMA_signal_19512 ;
    wire new_AGEMA_signal_19513 ;
    wire new_AGEMA_signal_19514 ;
    wire new_AGEMA_signal_19515 ;
    wire new_AGEMA_signal_19516 ;
    wire new_AGEMA_signal_19517 ;
    wire new_AGEMA_signal_19518 ;
    wire new_AGEMA_signal_19519 ;
    wire new_AGEMA_signal_19520 ;
    wire new_AGEMA_signal_19521 ;
    wire new_AGEMA_signal_19522 ;
    wire new_AGEMA_signal_19523 ;
    wire new_AGEMA_signal_19524 ;
    wire new_AGEMA_signal_19525 ;
    wire new_AGEMA_signal_19526 ;
    wire new_AGEMA_signal_19527 ;
    wire new_AGEMA_signal_19528 ;
    wire new_AGEMA_signal_19529 ;
    wire new_AGEMA_signal_19530 ;
    wire new_AGEMA_signal_19531 ;
    wire new_AGEMA_signal_19532 ;
    wire new_AGEMA_signal_19533 ;
    wire new_AGEMA_signal_19534 ;
    wire new_AGEMA_signal_19535 ;
    wire new_AGEMA_signal_19536 ;
    wire new_AGEMA_signal_19537 ;
    wire new_AGEMA_signal_19541 ;
    wire new_AGEMA_signal_19542 ;
    wire new_AGEMA_signal_19543 ;
    wire new_AGEMA_signal_19550 ;
    wire new_AGEMA_signal_19551 ;
    wire new_AGEMA_signal_19552 ;
    wire new_AGEMA_signal_19553 ;
    wire new_AGEMA_signal_19554 ;
    wire new_AGEMA_signal_19555 ;
    wire new_AGEMA_signal_19559 ;
    wire new_AGEMA_signal_19560 ;
    wire new_AGEMA_signal_19561 ;
    wire new_AGEMA_signal_19562 ;
    wire new_AGEMA_signal_19563 ;
    wire new_AGEMA_signal_19564 ;
    wire new_AGEMA_signal_19565 ;
    wire new_AGEMA_signal_19566 ;
    wire new_AGEMA_signal_19567 ;
    wire new_AGEMA_signal_19568 ;
    wire new_AGEMA_signal_19569 ;
    wire new_AGEMA_signal_19570 ;
    wire new_AGEMA_signal_19571 ;
    wire new_AGEMA_signal_19572 ;
    wire new_AGEMA_signal_19573 ;
    wire new_AGEMA_signal_19574 ;
    wire new_AGEMA_signal_19575 ;
    wire new_AGEMA_signal_19576 ;
    wire new_AGEMA_signal_19577 ;
    wire new_AGEMA_signal_19578 ;
    wire new_AGEMA_signal_19579 ;
    wire new_AGEMA_signal_19583 ;
    wire new_AGEMA_signal_19584 ;
    wire new_AGEMA_signal_19585 ;
    wire new_AGEMA_signal_19589 ;
    wire new_AGEMA_signal_19590 ;
    wire new_AGEMA_signal_19591 ;
    wire new_AGEMA_signal_19592 ;
    wire new_AGEMA_signal_19593 ;
    wire new_AGEMA_signal_19594 ;
    wire new_AGEMA_signal_19595 ;
    wire new_AGEMA_signal_19596 ;
    wire new_AGEMA_signal_19597 ;
    wire new_AGEMA_signal_19598 ;
    wire new_AGEMA_signal_19599 ;
    wire new_AGEMA_signal_19600 ;
    wire new_AGEMA_signal_19601 ;
    wire new_AGEMA_signal_19602 ;
    wire new_AGEMA_signal_19603 ;
    wire new_AGEMA_signal_19604 ;
    wire new_AGEMA_signal_19605 ;
    wire new_AGEMA_signal_19606 ;
    wire new_AGEMA_signal_19607 ;
    wire new_AGEMA_signal_19608 ;
    wire new_AGEMA_signal_19609 ;
    wire new_AGEMA_signal_19616 ;
    wire new_AGEMA_signal_19617 ;
    wire new_AGEMA_signal_19618 ;
    wire new_AGEMA_signal_19625 ;
    wire new_AGEMA_signal_19626 ;
    wire new_AGEMA_signal_19627 ;
    wire new_AGEMA_signal_19628 ;
    wire new_AGEMA_signal_19629 ;
    wire new_AGEMA_signal_19630 ;
    wire new_AGEMA_signal_19631 ;
    wire new_AGEMA_signal_19632 ;
    wire new_AGEMA_signal_19633 ;
    wire new_AGEMA_signal_19634 ;
    wire new_AGEMA_signal_19635 ;
    wire new_AGEMA_signal_19636 ;
    wire new_AGEMA_signal_19637 ;
    wire new_AGEMA_signal_19638 ;
    wire new_AGEMA_signal_19639 ;
    wire new_AGEMA_signal_19640 ;
    wire new_AGEMA_signal_19641 ;
    wire new_AGEMA_signal_19642 ;
    wire new_AGEMA_signal_19643 ;
    wire new_AGEMA_signal_19644 ;
    wire new_AGEMA_signal_19645 ;
    wire new_AGEMA_signal_19646 ;
    wire new_AGEMA_signal_19647 ;
    wire new_AGEMA_signal_19648 ;
    wire new_AGEMA_signal_19649 ;
    wire new_AGEMA_signal_19650 ;
    wire new_AGEMA_signal_19651 ;
    wire new_AGEMA_signal_19652 ;
    wire new_AGEMA_signal_19653 ;
    wire new_AGEMA_signal_19654 ;
    wire new_AGEMA_signal_19655 ;
    wire new_AGEMA_signal_19656 ;
    wire new_AGEMA_signal_19657 ;
    wire new_AGEMA_signal_19658 ;
    wire new_AGEMA_signal_19659 ;
    wire new_AGEMA_signal_19660 ;
    wire new_AGEMA_signal_19661 ;
    wire new_AGEMA_signal_19662 ;
    wire new_AGEMA_signal_19663 ;
    wire new_AGEMA_signal_19664 ;
    wire new_AGEMA_signal_19665 ;
    wire new_AGEMA_signal_19666 ;
    wire new_AGEMA_signal_19667 ;
    wire new_AGEMA_signal_19668 ;
    wire new_AGEMA_signal_19669 ;
    wire new_AGEMA_signal_19670 ;
    wire new_AGEMA_signal_19671 ;
    wire new_AGEMA_signal_19672 ;
    wire new_AGEMA_signal_19673 ;
    wire new_AGEMA_signal_19674 ;
    wire new_AGEMA_signal_19675 ;
    wire new_AGEMA_signal_19676 ;
    wire new_AGEMA_signal_19677 ;
    wire new_AGEMA_signal_19678 ;
    wire new_AGEMA_signal_19679 ;
    wire new_AGEMA_signal_19680 ;
    wire new_AGEMA_signal_19681 ;
    wire new_AGEMA_signal_19682 ;
    wire new_AGEMA_signal_19683 ;
    wire new_AGEMA_signal_19684 ;
    wire new_AGEMA_signal_19685 ;
    wire new_AGEMA_signal_19686 ;
    wire new_AGEMA_signal_19687 ;
    wire new_AGEMA_signal_19694 ;
    wire new_AGEMA_signal_19695 ;
    wire new_AGEMA_signal_19696 ;
    wire new_AGEMA_signal_19700 ;
    wire new_AGEMA_signal_19701 ;
    wire new_AGEMA_signal_19702 ;
    wire new_AGEMA_signal_19703 ;
    wire new_AGEMA_signal_19704 ;
    wire new_AGEMA_signal_19705 ;
    wire new_AGEMA_signal_19706 ;
    wire new_AGEMA_signal_19707 ;
    wire new_AGEMA_signal_19708 ;
    wire new_AGEMA_signal_19709 ;
    wire new_AGEMA_signal_19710 ;
    wire new_AGEMA_signal_19711 ;
    wire new_AGEMA_signal_19712 ;
    wire new_AGEMA_signal_19713 ;
    wire new_AGEMA_signal_19714 ;
    wire new_AGEMA_signal_19718 ;
    wire new_AGEMA_signal_19719 ;
    wire new_AGEMA_signal_19720 ;
    wire new_AGEMA_signal_19727 ;
    wire new_AGEMA_signal_19728 ;
    wire new_AGEMA_signal_19729 ;
    wire new_AGEMA_signal_19730 ;
    wire new_AGEMA_signal_19731 ;
    wire new_AGEMA_signal_19732 ;
    wire new_AGEMA_signal_19733 ;
    wire new_AGEMA_signal_19734 ;
    wire new_AGEMA_signal_19735 ;
    wire new_AGEMA_signal_19736 ;
    wire new_AGEMA_signal_19737 ;
    wire new_AGEMA_signal_19738 ;
    wire new_AGEMA_signal_19739 ;
    wire new_AGEMA_signal_19740 ;
    wire new_AGEMA_signal_19741 ;
    wire new_AGEMA_signal_19742 ;
    wire new_AGEMA_signal_19743 ;
    wire new_AGEMA_signal_19744 ;
    wire new_AGEMA_signal_19745 ;
    wire new_AGEMA_signal_19746 ;
    wire new_AGEMA_signal_19747 ;
    wire new_AGEMA_signal_19748 ;
    wire new_AGEMA_signal_19749 ;
    wire new_AGEMA_signal_19750 ;
    wire new_AGEMA_signal_19751 ;
    wire new_AGEMA_signal_19752 ;
    wire new_AGEMA_signal_19753 ;
    wire new_AGEMA_signal_19754 ;
    wire new_AGEMA_signal_19755 ;
    wire new_AGEMA_signal_19756 ;
    wire new_AGEMA_signal_19757 ;
    wire new_AGEMA_signal_19758 ;
    wire new_AGEMA_signal_19759 ;
    wire new_AGEMA_signal_19763 ;
    wire new_AGEMA_signal_19764 ;
    wire new_AGEMA_signal_19765 ;
    wire new_AGEMA_signal_19766 ;
    wire new_AGEMA_signal_19767 ;
    wire new_AGEMA_signal_19768 ;
    wire new_AGEMA_signal_19769 ;
    wire new_AGEMA_signal_19770 ;
    wire new_AGEMA_signal_19771 ;
    wire new_AGEMA_signal_19772 ;
    wire new_AGEMA_signal_19773 ;
    wire new_AGEMA_signal_19774 ;
    wire new_AGEMA_signal_19775 ;
    wire new_AGEMA_signal_19776 ;
    wire new_AGEMA_signal_19777 ;
    wire new_AGEMA_signal_19784 ;
    wire new_AGEMA_signal_19785 ;
    wire new_AGEMA_signal_19786 ;
    wire new_AGEMA_signal_19787 ;
    wire new_AGEMA_signal_19788 ;
    wire new_AGEMA_signal_19789 ;
    wire new_AGEMA_signal_19790 ;
    wire new_AGEMA_signal_19791 ;
    wire new_AGEMA_signal_19792 ;
    wire new_AGEMA_signal_19793 ;
    wire new_AGEMA_signal_19794 ;
    wire new_AGEMA_signal_19795 ;
    wire new_AGEMA_signal_19796 ;
    wire new_AGEMA_signal_19797 ;
    wire new_AGEMA_signal_19798 ;
    wire new_AGEMA_signal_19799 ;
    wire new_AGEMA_signal_19800 ;
    wire new_AGEMA_signal_19801 ;
    wire new_AGEMA_signal_19802 ;
    wire new_AGEMA_signal_19803 ;
    wire new_AGEMA_signal_19804 ;
    wire new_AGEMA_signal_19805 ;
    wire new_AGEMA_signal_19806 ;
    wire new_AGEMA_signal_19807 ;
    wire new_AGEMA_signal_19808 ;
    wire new_AGEMA_signal_19809 ;
    wire new_AGEMA_signal_19810 ;
    wire new_AGEMA_signal_19811 ;
    wire new_AGEMA_signal_19812 ;
    wire new_AGEMA_signal_19813 ;
    wire new_AGEMA_signal_19814 ;
    wire new_AGEMA_signal_19815 ;
    wire new_AGEMA_signal_19816 ;
    wire new_AGEMA_signal_19817 ;
    wire new_AGEMA_signal_19818 ;
    wire new_AGEMA_signal_19819 ;
    wire new_AGEMA_signal_19820 ;
    wire new_AGEMA_signal_19821 ;
    wire new_AGEMA_signal_19822 ;
    wire new_AGEMA_signal_19826 ;
    wire new_AGEMA_signal_19827 ;
    wire new_AGEMA_signal_19828 ;
    wire new_AGEMA_signal_19835 ;
    wire new_AGEMA_signal_19836 ;
    wire new_AGEMA_signal_19837 ;
    wire new_AGEMA_signal_19838 ;
    wire new_AGEMA_signal_19839 ;
    wire new_AGEMA_signal_19840 ;
    wire new_AGEMA_signal_19844 ;
    wire new_AGEMA_signal_19845 ;
    wire new_AGEMA_signal_19846 ;
    wire new_AGEMA_signal_19847 ;
    wire new_AGEMA_signal_19848 ;
    wire new_AGEMA_signal_19849 ;
    wire new_AGEMA_signal_19850 ;
    wire new_AGEMA_signal_19851 ;
    wire new_AGEMA_signal_19852 ;
    wire new_AGEMA_signal_19853 ;
    wire new_AGEMA_signal_19854 ;
    wire new_AGEMA_signal_19855 ;
    wire new_AGEMA_signal_19856 ;
    wire new_AGEMA_signal_19857 ;
    wire new_AGEMA_signal_19858 ;
    wire new_AGEMA_signal_19859 ;
    wire new_AGEMA_signal_19860 ;
    wire new_AGEMA_signal_19861 ;
    wire new_AGEMA_signal_19862 ;
    wire new_AGEMA_signal_19863 ;
    wire new_AGEMA_signal_19864 ;
    wire new_AGEMA_signal_19868 ;
    wire new_AGEMA_signal_19869 ;
    wire new_AGEMA_signal_19870 ;
    wire new_AGEMA_signal_19874 ;
    wire new_AGEMA_signal_19875 ;
    wire new_AGEMA_signal_19876 ;
    wire new_AGEMA_signal_19877 ;
    wire new_AGEMA_signal_19878 ;
    wire new_AGEMA_signal_19879 ;
    wire new_AGEMA_signal_19880 ;
    wire new_AGEMA_signal_19881 ;
    wire new_AGEMA_signal_19882 ;
    wire new_AGEMA_signal_19883 ;
    wire new_AGEMA_signal_19884 ;
    wire new_AGEMA_signal_19885 ;
    wire new_AGEMA_signal_19886 ;
    wire new_AGEMA_signal_19887 ;
    wire new_AGEMA_signal_19888 ;
    wire new_AGEMA_signal_19889 ;
    wire new_AGEMA_signal_19890 ;
    wire new_AGEMA_signal_19891 ;
    wire new_AGEMA_signal_19892 ;
    wire new_AGEMA_signal_19893 ;
    wire new_AGEMA_signal_19894 ;
    wire new_AGEMA_signal_19901 ;
    wire new_AGEMA_signal_19902 ;
    wire new_AGEMA_signal_19903 ;
    wire new_AGEMA_signal_19910 ;
    wire new_AGEMA_signal_19911 ;
    wire new_AGEMA_signal_19912 ;
    wire new_AGEMA_signal_19913 ;
    wire new_AGEMA_signal_19914 ;
    wire new_AGEMA_signal_19915 ;
    wire new_AGEMA_signal_19916 ;
    wire new_AGEMA_signal_19917 ;
    wire new_AGEMA_signal_19918 ;
    wire new_AGEMA_signal_19919 ;
    wire new_AGEMA_signal_19920 ;
    wire new_AGEMA_signal_19921 ;
    wire new_AGEMA_signal_19922 ;
    wire new_AGEMA_signal_19923 ;
    wire new_AGEMA_signal_19924 ;
    wire new_AGEMA_signal_19925 ;
    wire new_AGEMA_signal_19926 ;
    wire new_AGEMA_signal_19927 ;
    wire new_AGEMA_signal_19928 ;
    wire new_AGEMA_signal_19929 ;
    wire new_AGEMA_signal_19930 ;
    wire new_AGEMA_signal_19931 ;
    wire new_AGEMA_signal_19932 ;
    wire new_AGEMA_signal_19933 ;
    wire new_AGEMA_signal_19934 ;
    wire new_AGEMA_signal_19935 ;
    wire new_AGEMA_signal_19936 ;
    wire new_AGEMA_signal_19937 ;
    wire new_AGEMA_signal_19938 ;
    wire new_AGEMA_signal_19939 ;
    wire new_AGEMA_signal_19940 ;
    wire new_AGEMA_signal_19941 ;
    wire new_AGEMA_signal_19942 ;
    wire new_AGEMA_signal_19943 ;
    wire new_AGEMA_signal_19944 ;
    wire new_AGEMA_signal_19945 ;
    wire new_AGEMA_signal_19946 ;
    wire new_AGEMA_signal_19947 ;
    wire new_AGEMA_signal_19948 ;
    wire new_AGEMA_signal_19949 ;
    wire new_AGEMA_signal_19950 ;
    wire new_AGEMA_signal_19951 ;
    wire new_AGEMA_signal_19952 ;
    wire new_AGEMA_signal_19953 ;
    wire new_AGEMA_signal_19954 ;
    wire new_AGEMA_signal_19955 ;
    wire new_AGEMA_signal_19956 ;
    wire new_AGEMA_signal_19957 ;
    wire new_AGEMA_signal_19958 ;
    wire new_AGEMA_signal_19959 ;
    wire new_AGEMA_signal_19960 ;
    wire new_AGEMA_signal_19961 ;
    wire new_AGEMA_signal_19962 ;
    wire new_AGEMA_signal_19963 ;
    wire new_AGEMA_signal_19964 ;
    wire new_AGEMA_signal_19965 ;
    wire new_AGEMA_signal_19966 ;
    wire new_AGEMA_signal_19967 ;
    wire new_AGEMA_signal_19968 ;
    wire new_AGEMA_signal_19969 ;
    wire new_AGEMA_signal_19970 ;
    wire new_AGEMA_signal_19971 ;
    wire new_AGEMA_signal_19972 ;
    wire new_AGEMA_signal_19979 ;
    wire new_AGEMA_signal_19980 ;
    wire new_AGEMA_signal_19981 ;
    wire new_AGEMA_signal_19985 ;
    wire new_AGEMA_signal_19986 ;
    wire new_AGEMA_signal_19987 ;
    wire new_AGEMA_signal_19988 ;
    wire new_AGEMA_signal_19989 ;
    wire new_AGEMA_signal_19990 ;
    wire new_AGEMA_signal_19991 ;
    wire new_AGEMA_signal_19992 ;
    wire new_AGEMA_signal_19993 ;
    wire new_AGEMA_signal_19994 ;
    wire new_AGEMA_signal_19995 ;
    wire new_AGEMA_signal_19996 ;
    wire new_AGEMA_signal_19997 ;
    wire new_AGEMA_signal_19998 ;
    wire new_AGEMA_signal_19999 ;
    wire new_AGEMA_signal_20003 ;
    wire new_AGEMA_signal_20004 ;
    wire new_AGEMA_signal_20005 ;
    wire new_AGEMA_signal_20012 ;
    wire new_AGEMA_signal_20013 ;
    wire new_AGEMA_signal_20014 ;
    wire new_AGEMA_signal_20015 ;
    wire new_AGEMA_signal_20016 ;
    wire new_AGEMA_signal_20017 ;
    wire new_AGEMA_signal_20018 ;
    wire new_AGEMA_signal_20019 ;
    wire new_AGEMA_signal_20020 ;
    wire new_AGEMA_signal_20021 ;
    wire new_AGEMA_signal_20022 ;
    wire new_AGEMA_signal_20023 ;
    wire new_AGEMA_signal_20024 ;
    wire new_AGEMA_signal_20025 ;
    wire new_AGEMA_signal_20026 ;
    wire new_AGEMA_signal_20027 ;
    wire new_AGEMA_signal_20028 ;
    wire new_AGEMA_signal_20029 ;
    wire new_AGEMA_signal_20030 ;
    wire new_AGEMA_signal_20031 ;
    wire new_AGEMA_signal_20032 ;
    wire new_AGEMA_signal_20033 ;
    wire new_AGEMA_signal_20034 ;
    wire new_AGEMA_signal_20035 ;
    wire new_AGEMA_signal_20036 ;
    wire new_AGEMA_signal_20037 ;
    wire new_AGEMA_signal_20038 ;
    wire new_AGEMA_signal_20039 ;
    wire new_AGEMA_signal_20040 ;
    wire new_AGEMA_signal_20041 ;
    wire new_AGEMA_signal_20078 ;
    wire new_AGEMA_signal_20079 ;
    wire new_AGEMA_signal_20080 ;
    wire new_AGEMA_signal_20081 ;
    wire new_AGEMA_signal_20082 ;
    wire new_AGEMA_signal_20083 ;
    wire new_AGEMA_signal_20084 ;
    wire new_AGEMA_signal_20085 ;
    wire new_AGEMA_signal_20086 ;
    wire new_AGEMA_signal_20087 ;
    wire new_AGEMA_signal_20088 ;
    wire new_AGEMA_signal_20089 ;
    wire new_AGEMA_signal_20090 ;
    wire new_AGEMA_signal_20091 ;
    wire new_AGEMA_signal_20092 ;
    wire new_AGEMA_signal_20093 ;
    wire new_AGEMA_signal_20094 ;
    wire new_AGEMA_signal_20095 ;
    wire new_AGEMA_signal_20096 ;
    wire new_AGEMA_signal_20097 ;
    wire new_AGEMA_signal_20098 ;
    wire new_AGEMA_signal_20099 ;
    wire new_AGEMA_signal_20100 ;
    wire new_AGEMA_signal_20101 ;
    wire new_AGEMA_signal_20102 ;
    wire new_AGEMA_signal_20103 ;
    wire new_AGEMA_signal_20104 ;
    wire new_AGEMA_signal_20105 ;
    wire new_AGEMA_signal_20106 ;
    wire new_AGEMA_signal_20107 ;
    wire new_AGEMA_signal_20108 ;
    wire new_AGEMA_signal_20109 ;
    wire new_AGEMA_signal_20110 ;
    wire new_AGEMA_signal_20111 ;
    wire new_AGEMA_signal_20112 ;
    wire new_AGEMA_signal_20113 ;
    wire new_AGEMA_signal_20114 ;
    wire new_AGEMA_signal_20115 ;
    wire new_AGEMA_signal_20116 ;
    wire new_AGEMA_signal_20117 ;
    wire new_AGEMA_signal_20118 ;
    wire new_AGEMA_signal_20119 ;
    wire new_AGEMA_signal_20120 ;
    wire new_AGEMA_signal_20121 ;
    wire new_AGEMA_signal_20122 ;
    wire new_AGEMA_signal_20123 ;
    wire new_AGEMA_signal_20124 ;
    wire new_AGEMA_signal_20125 ;
    wire new_AGEMA_signal_20126 ;
    wire new_AGEMA_signal_20127 ;
    wire new_AGEMA_signal_20128 ;
    wire new_AGEMA_signal_20129 ;
    wire new_AGEMA_signal_20130 ;
    wire new_AGEMA_signal_20131 ;
    wire new_AGEMA_signal_20360 ;
    wire new_AGEMA_signal_20361 ;
    wire new_AGEMA_signal_20362 ;
    wire new_AGEMA_signal_20366 ;
    wire new_AGEMA_signal_20367 ;
    wire new_AGEMA_signal_20368 ;
    wire new_AGEMA_signal_20369 ;
    wire new_AGEMA_signal_20370 ;
    wire new_AGEMA_signal_20371 ;
    wire new_AGEMA_signal_20375 ;
    wire new_AGEMA_signal_20376 ;
    wire new_AGEMA_signal_20377 ;
    wire new_AGEMA_signal_20378 ;
    wire new_AGEMA_signal_20379 ;
    wire new_AGEMA_signal_20380 ;
    wire new_AGEMA_signal_20381 ;
    wire new_AGEMA_signal_20382 ;
    wire new_AGEMA_signal_20383 ;
    wire new_AGEMA_signal_20384 ;
    wire new_AGEMA_signal_20385 ;
    wire new_AGEMA_signal_20386 ;
    wire new_AGEMA_signal_20387 ;
    wire new_AGEMA_signal_20388 ;
    wire new_AGEMA_signal_20389 ;
    wire new_AGEMA_signal_20390 ;
    wire new_AGEMA_signal_20391 ;
    wire new_AGEMA_signal_20392 ;
    wire new_AGEMA_signal_20396 ;
    wire new_AGEMA_signal_20397 ;
    wire new_AGEMA_signal_20398 ;
    wire new_AGEMA_signal_20399 ;
    wire new_AGEMA_signal_20400 ;
    wire new_AGEMA_signal_20401 ;
    wire new_AGEMA_signal_20405 ;
    wire new_AGEMA_signal_20406 ;
    wire new_AGEMA_signal_20407 ;
    wire new_AGEMA_signal_20411 ;
    wire new_AGEMA_signal_20412 ;
    wire new_AGEMA_signal_20413 ;
    wire new_AGEMA_signal_20414 ;
    wire new_AGEMA_signal_20415 ;
    wire new_AGEMA_signal_20416 ;
    wire new_AGEMA_signal_20420 ;
    wire new_AGEMA_signal_20421 ;
    wire new_AGEMA_signal_20422 ;
    wire new_AGEMA_signal_20423 ;
    wire new_AGEMA_signal_20424 ;
    wire new_AGEMA_signal_20425 ;
    wire new_AGEMA_signal_20426 ;
    wire new_AGEMA_signal_20427 ;
    wire new_AGEMA_signal_20428 ;
    wire new_AGEMA_signal_20429 ;
    wire new_AGEMA_signal_20430 ;
    wire new_AGEMA_signal_20431 ;
    wire new_AGEMA_signal_20432 ;
    wire new_AGEMA_signal_20433 ;
    wire new_AGEMA_signal_20434 ;
    wire new_AGEMA_signal_20438 ;
    wire new_AGEMA_signal_20439 ;
    wire new_AGEMA_signal_20440 ;
    wire new_AGEMA_signal_20441 ;
    wire new_AGEMA_signal_20442 ;
    wire new_AGEMA_signal_20443 ;
    wire new_AGEMA_signal_20450 ;
    wire new_AGEMA_signal_20451 ;
    wire new_AGEMA_signal_20452 ;
    wire new_AGEMA_signal_20453 ;
    wire new_AGEMA_signal_20454 ;
    wire new_AGEMA_signal_20455 ;
    wire new_AGEMA_signal_20456 ;
    wire new_AGEMA_signal_20457 ;
    wire new_AGEMA_signal_20458 ;
    wire new_AGEMA_signal_20459 ;
    wire new_AGEMA_signal_20460 ;
    wire new_AGEMA_signal_20461 ;
    wire new_AGEMA_signal_20465 ;
    wire new_AGEMA_signal_20466 ;
    wire new_AGEMA_signal_20467 ;
    wire new_AGEMA_signal_20468 ;
    wire new_AGEMA_signal_20469 ;
    wire new_AGEMA_signal_20470 ;
    wire new_AGEMA_signal_20471 ;
    wire new_AGEMA_signal_20472 ;
    wire new_AGEMA_signal_20473 ;
    wire new_AGEMA_signal_20474 ;
    wire new_AGEMA_signal_20475 ;
    wire new_AGEMA_signal_20476 ;
    wire new_AGEMA_signal_20477 ;
    wire new_AGEMA_signal_20478 ;
    wire new_AGEMA_signal_20479 ;
    wire new_AGEMA_signal_20480 ;
    wire new_AGEMA_signal_20481 ;
    wire new_AGEMA_signal_20482 ;
    wire new_AGEMA_signal_20483 ;
    wire new_AGEMA_signal_20484 ;
    wire new_AGEMA_signal_20485 ;
    wire new_AGEMA_signal_20486 ;
    wire new_AGEMA_signal_20487 ;
    wire new_AGEMA_signal_20488 ;
    wire new_AGEMA_signal_20489 ;
    wire new_AGEMA_signal_20490 ;
    wire new_AGEMA_signal_20491 ;
    wire new_AGEMA_signal_20492 ;
    wire new_AGEMA_signal_20493 ;
    wire new_AGEMA_signal_20494 ;
    wire new_AGEMA_signal_20495 ;
    wire new_AGEMA_signal_20496 ;
    wire new_AGEMA_signal_20497 ;
    wire new_AGEMA_signal_20501 ;
    wire new_AGEMA_signal_20502 ;
    wire new_AGEMA_signal_20503 ;
    wire new_AGEMA_signal_20504 ;
    wire new_AGEMA_signal_20505 ;
    wire new_AGEMA_signal_20506 ;
    wire new_AGEMA_signal_20510 ;
    wire new_AGEMA_signal_20511 ;
    wire new_AGEMA_signal_20512 ;
    wire new_AGEMA_signal_20513 ;
    wire new_AGEMA_signal_20514 ;
    wire new_AGEMA_signal_20515 ;
    wire new_AGEMA_signal_20522 ;
    wire new_AGEMA_signal_20523 ;
    wire new_AGEMA_signal_20524 ;
    wire new_AGEMA_signal_20525 ;
    wire new_AGEMA_signal_20526 ;
    wire new_AGEMA_signal_20527 ;
    wire new_AGEMA_signal_20531 ;
    wire new_AGEMA_signal_20532 ;
    wire new_AGEMA_signal_20533 ;
    wire new_AGEMA_signal_20534 ;
    wire new_AGEMA_signal_20535 ;
    wire new_AGEMA_signal_20536 ;
    wire new_AGEMA_signal_20537 ;
    wire new_AGEMA_signal_20538 ;
    wire new_AGEMA_signal_20539 ;
    wire new_AGEMA_signal_20540 ;
    wire new_AGEMA_signal_20541 ;
    wire new_AGEMA_signal_20542 ;
    wire new_AGEMA_signal_20543 ;
    wire new_AGEMA_signal_20544 ;
    wire new_AGEMA_signal_20545 ;
    wire new_AGEMA_signal_20546 ;
    wire new_AGEMA_signal_20547 ;
    wire new_AGEMA_signal_20548 ;
    wire new_AGEMA_signal_20549 ;
    wire new_AGEMA_signal_20550 ;
    wire new_AGEMA_signal_20551 ;
    wire new_AGEMA_signal_20552 ;
    wire new_AGEMA_signal_20553 ;
    wire new_AGEMA_signal_20554 ;
    wire new_AGEMA_signal_20564 ;
    wire new_AGEMA_signal_20565 ;
    wire new_AGEMA_signal_20566 ;
    wire new_AGEMA_signal_20567 ;
    wire new_AGEMA_signal_20568 ;
    wire new_AGEMA_signal_20569 ;
    wire new_AGEMA_signal_20573 ;
    wire new_AGEMA_signal_20574 ;
    wire new_AGEMA_signal_20575 ;
    wire new_AGEMA_signal_20576 ;
    wire new_AGEMA_signal_20577 ;
    wire new_AGEMA_signal_20578 ;
    wire new_AGEMA_signal_20582 ;
    wire new_AGEMA_signal_20583 ;
    wire new_AGEMA_signal_20584 ;
    wire new_AGEMA_signal_20585 ;
    wire new_AGEMA_signal_20586 ;
    wire new_AGEMA_signal_20587 ;
    wire new_AGEMA_signal_20588 ;
    wire new_AGEMA_signal_20589 ;
    wire new_AGEMA_signal_20590 ;
    wire new_AGEMA_signal_20591 ;
    wire new_AGEMA_signal_20592 ;
    wire new_AGEMA_signal_20593 ;
    wire new_AGEMA_signal_20594 ;
    wire new_AGEMA_signal_20595 ;
    wire new_AGEMA_signal_20596 ;
    wire new_AGEMA_signal_20597 ;
    wire new_AGEMA_signal_20598 ;
    wire new_AGEMA_signal_20599 ;
    wire new_AGEMA_signal_20603 ;
    wire new_AGEMA_signal_20604 ;
    wire new_AGEMA_signal_20605 ;
    wire new_AGEMA_signal_20606 ;
    wire new_AGEMA_signal_20607 ;
    wire new_AGEMA_signal_20608 ;
    wire new_AGEMA_signal_20612 ;
    wire new_AGEMA_signal_20613 ;
    wire new_AGEMA_signal_20614 ;
    wire new_AGEMA_signal_20618 ;
    wire new_AGEMA_signal_20619 ;
    wire new_AGEMA_signal_20620 ;
    wire new_AGEMA_signal_20621 ;
    wire new_AGEMA_signal_20622 ;
    wire new_AGEMA_signal_20623 ;
    wire new_AGEMA_signal_20627 ;
    wire new_AGEMA_signal_20628 ;
    wire new_AGEMA_signal_20629 ;
    wire new_AGEMA_signal_20630 ;
    wire new_AGEMA_signal_20631 ;
    wire new_AGEMA_signal_20632 ;
    wire new_AGEMA_signal_20633 ;
    wire new_AGEMA_signal_20634 ;
    wire new_AGEMA_signal_20635 ;
    wire new_AGEMA_signal_20636 ;
    wire new_AGEMA_signal_20637 ;
    wire new_AGEMA_signal_20638 ;
    wire new_AGEMA_signal_20639 ;
    wire new_AGEMA_signal_20640 ;
    wire new_AGEMA_signal_20641 ;
    wire new_AGEMA_signal_20645 ;
    wire new_AGEMA_signal_20646 ;
    wire new_AGEMA_signal_20647 ;
    wire new_AGEMA_signal_20648 ;
    wire new_AGEMA_signal_20649 ;
    wire new_AGEMA_signal_20650 ;
    wire new_AGEMA_signal_20657 ;
    wire new_AGEMA_signal_20658 ;
    wire new_AGEMA_signal_20659 ;
    wire new_AGEMA_signal_20660 ;
    wire new_AGEMA_signal_20661 ;
    wire new_AGEMA_signal_20662 ;
    wire new_AGEMA_signal_20663 ;
    wire new_AGEMA_signal_20664 ;
    wire new_AGEMA_signal_20665 ;
    wire new_AGEMA_signal_20666 ;
    wire new_AGEMA_signal_20667 ;
    wire new_AGEMA_signal_20668 ;
    wire new_AGEMA_signal_20672 ;
    wire new_AGEMA_signal_20673 ;
    wire new_AGEMA_signal_20674 ;
    wire new_AGEMA_signal_20675 ;
    wire new_AGEMA_signal_20676 ;
    wire new_AGEMA_signal_20677 ;
    wire new_AGEMA_signal_20678 ;
    wire new_AGEMA_signal_20679 ;
    wire new_AGEMA_signal_20680 ;
    wire new_AGEMA_signal_20681 ;
    wire new_AGEMA_signal_20682 ;
    wire new_AGEMA_signal_20683 ;
    wire new_AGEMA_signal_20684 ;
    wire new_AGEMA_signal_20685 ;
    wire new_AGEMA_signal_20686 ;
    wire new_AGEMA_signal_20687 ;
    wire new_AGEMA_signal_20688 ;
    wire new_AGEMA_signal_20689 ;
    wire new_AGEMA_signal_20690 ;
    wire new_AGEMA_signal_20691 ;
    wire new_AGEMA_signal_20692 ;
    wire new_AGEMA_signal_20693 ;
    wire new_AGEMA_signal_20694 ;
    wire new_AGEMA_signal_20695 ;
    wire new_AGEMA_signal_20696 ;
    wire new_AGEMA_signal_20697 ;
    wire new_AGEMA_signal_20698 ;
    wire new_AGEMA_signal_20699 ;
    wire new_AGEMA_signal_20700 ;
    wire new_AGEMA_signal_20701 ;
    wire new_AGEMA_signal_20702 ;
    wire new_AGEMA_signal_20703 ;
    wire new_AGEMA_signal_20704 ;
    wire new_AGEMA_signal_20708 ;
    wire new_AGEMA_signal_20709 ;
    wire new_AGEMA_signal_20710 ;
    wire new_AGEMA_signal_20711 ;
    wire new_AGEMA_signal_20712 ;
    wire new_AGEMA_signal_20713 ;
    wire new_AGEMA_signal_20717 ;
    wire new_AGEMA_signal_20718 ;
    wire new_AGEMA_signal_20719 ;
    wire new_AGEMA_signal_20720 ;
    wire new_AGEMA_signal_20721 ;
    wire new_AGEMA_signal_20722 ;
    wire new_AGEMA_signal_20729 ;
    wire new_AGEMA_signal_20730 ;
    wire new_AGEMA_signal_20731 ;
    wire new_AGEMA_signal_20732 ;
    wire new_AGEMA_signal_20733 ;
    wire new_AGEMA_signal_20734 ;
    wire new_AGEMA_signal_20738 ;
    wire new_AGEMA_signal_20739 ;
    wire new_AGEMA_signal_20740 ;
    wire new_AGEMA_signal_20741 ;
    wire new_AGEMA_signal_20742 ;
    wire new_AGEMA_signal_20743 ;
    wire new_AGEMA_signal_20744 ;
    wire new_AGEMA_signal_20745 ;
    wire new_AGEMA_signal_20746 ;
    wire new_AGEMA_signal_20747 ;
    wire new_AGEMA_signal_20748 ;
    wire new_AGEMA_signal_20749 ;
    wire new_AGEMA_signal_20750 ;
    wire new_AGEMA_signal_20751 ;
    wire new_AGEMA_signal_20752 ;
    wire new_AGEMA_signal_20753 ;
    wire new_AGEMA_signal_20754 ;
    wire new_AGEMA_signal_20755 ;
    wire new_AGEMA_signal_20756 ;
    wire new_AGEMA_signal_20757 ;
    wire new_AGEMA_signal_20758 ;
    wire new_AGEMA_signal_20759 ;
    wire new_AGEMA_signal_20760 ;
    wire new_AGEMA_signal_20761 ;
    wire new_AGEMA_signal_20771 ;
    wire new_AGEMA_signal_20772 ;
    wire new_AGEMA_signal_20773 ;
    wire new_AGEMA_signal_20828 ;
    wire new_AGEMA_signal_20829 ;
    wire new_AGEMA_signal_20830 ;
    wire new_AGEMA_signal_20831 ;
    wire new_AGEMA_signal_20832 ;
    wire new_AGEMA_signal_20833 ;
    wire new_AGEMA_signal_20834 ;
    wire new_AGEMA_signal_20835 ;
    wire new_AGEMA_signal_20836 ;
    wire new_AGEMA_signal_20837 ;
    wire new_AGEMA_signal_20838 ;
    wire new_AGEMA_signal_20839 ;
    wire new_AGEMA_signal_20840 ;
    wire new_AGEMA_signal_20841 ;
    wire new_AGEMA_signal_20842 ;
    wire new_AGEMA_signal_20843 ;
    wire new_AGEMA_signal_20844 ;
    wire new_AGEMA_signal_20845 ;
    wire new_AGEMA_signal_20846 ;
    wire new_AGEMA_signal_20847 ;
    wire new_AGEMA_signal_20848 ;
    wire new_AGEMA_signal_20849 ;
    wire new_AGEMA_signal_20850 ;
    wire new_AGEMA_signal_20851 ;
    wire new_AGEMA_signal_20852 ;
    wire new_AGEMA_signal_20853 ;
    wire new_AGEMA_signal_20854 ;
    wire new_AGEMA_signal_20855 ;
    wire new_AGEMA_signal_20856 ;
    wire new_AGEMA_signal_20857 ;
    wire new_AGEMA_signal_20858 ;
    wire new_AGEMA_signal_20859 ;
    wire new_AGEMA_signal_20860 ;
    wire new_AGEMA_signal_20861 ;
    wire new_AGEMA_signal_20862 ;
    wire new_AGEMA_signal_20863 ;
    wire new_AGEMA_signal_20864 ;
    wire new_AGEMA_signal_20865 ;
    wire new_AGEMA_signal_20866 ;
    wire new_AGEMA_signal_20867 ;
    wire new_AGEMA_signal_20868 ;
    wire new_AGEMA_signal_20869 ;
    wire new_AGEMA_signal_20870 ;
    wire new_AGEMA_signal_20871 ;
    wire new_AGEMA_signal_20872 ;
    wire new_AGEMA_signal_20873 ;
    wire new_AGEMA_signal_20874 ;
    wire new_AGEMA_signal_20875 ;
    wire new_AGEMA_signal_20876 ;
    wire new_AGEMA_signal_20877 ;
    wire new_AGEMA_signal_20878 ;
    wire new_AGEMA_signal_20879 ;
    wire new_AGEMA_signal_20880 ;
    wire new_AGEMA_signal_20881 ;
    wire new_AGEMA_signal_20882 ;
    wire new_AGEMA_signal_20883 ;
    wire new_AGEMA_signal_20884 ;
    wire new_AGEMA_signal_20885 ;
    wire new_AGEMA_signal_20886 ;
    wire new_AGEMA_signal_20887 ;
    wire new_AGEMA_signal_20888 ;
    wire new_AGEMA_signal_20889 ;
    wire new_AGEMA_signal_20890 ;
    wire new_AGEMA_signal_20891 ;
    wire new_AGEMA_signal_20892 ;
    wire new_AGEMA_signal_20893 ;
    wire new_AGEMA_signal_20894 ;
    wire new_AGEMA_signal_20895 ;
    wire new_AGEMA_signal_20896 ;
    wire new_AGEMA_signal_20897 ;
    wire new_AGEMA_signal_20898 ;
    wire new_AGEMA_signal_20899 ;
    wire new_AGEMA_signal_20900 ;
    wire new_AGEMA_signal_20901 ;
    wire new_AGEMA_signal_20902 ;
    wire new_AGEMA_signal_20903 ;
    wire new_AGEMA_signal_20904 ;
    wire new_AGEMA_signal_20905 ;
    wire new_AGEMA_signal_20906 ;
    wire new_AGEMA_signal_20907 ;
    wire new_AGEMA_signal_20908 ;
    wire new_AGEMA_signal_20909 ;
    wire new_AGEMA_signal_20910 ;
    wire new_AGEMA_signal_20911 ;
    wire new_AGEMA_signal_21128 ;
    wire new_AGEMA_signal_21129 ;
    wire new_AGEMA_signal_21130 ;
    wire new_AGEMA_signal_21140 ;
    wire new_AGEMA_signal_21141 ;
    wire new_AGEMA_signal_21142 ;
    wire new_AGEMA_signal_21143 ;
    wire new_AGEMA_signal_21144 ;
    wire new_AGEMA_signal_21145 ;
    wire new_AGEMA_signal_21146 ;
    wire new_AGEMA_signal_21147 ;
    wire new_AGEMA_signal_21148 ;
    wire new_AGEMA_signal_21149 ;
    wire new_AGEMA_signal_21150 ;
    wire new_AGEMA_signal_21151 ;
    wire new_AGEMA_signal_21152 ;
    wire new_AGEMA_signal_21153 ;
    wire new_AGEMA_signal_21154 ;
    wire new_AGEMA_signal_21155 ;
    wire new_AGEMA_signal_21156 ;
    wire new_AGEMA_signal_21157 ;
    wire new_AGEMA_signal_21161 ;
    wire new_AGEMA_signal_21162 ;
    wire new_AGEMA_signal_21163 ;
    wire new_AGEMA_signal_21164 ;
    wire new_AGEMA_signal_21165 ;
    wire new_AGEMA_signal_21166 ;
    wire new_AGEMA_signal_21170 ;
    wire new_AGEMA_signal_21171 ;
    wire new_AGEMA_signal_21172 ;
    wire new_AGEMA_signal_21173 ;
    wire new_AGEMA_signal_21174 ;
    wire new_AGEMA_signal_21175 ;
    wire new_AGEMA_signal_21176 ;
    wire new_AGEMA_signal_21177 ;
    wire new_AGEMA_signal_21178 ;
    wire new_AGEMA_signal_21179 ;
    wire new_AGEMA_signal_21180 ;
    wire new_AGEMA_signal_21181 ;
    wire new_AGEMA_signal_21182 ;
    wire new_AGEMA_signal_21183 ;
    wire new_AGEMA_signal_21184 ;
    wire new_AGEMA_signal_21194 ;
    wire new_AGEMA_signal_21195 ;
    wire new_AGEMA_signal_21196 ;
    wire new_AGEMA_signal_21197 ;
    wire new_AGEMA_signal_21198 ;
    wire new_AGEMA_signal_21199 ;
    wire new_AGEMA_signal_21200 ;
    wire new_AGEMA_signal_21201 ;
    wire new_AGEMA_signal_21202 ;
    wire new_AGEMA_signal_21203 ;
    wire new_AGEMA_signal_21204 ;
    wire new_AGEMA_signal_21205 ;
    wire new_AGEMA_signal_21215 ;
    wire new_AGEMA_signal_21216 ;
    wire new_AGEMA_signal_21217 ;
    wire new_AGEMA_signal_21221 ;
    wire new_AGEMA_signal_21222 ;
    wire new_AGEMA_signal_21223 ;
    wire new_AGEMA_signal_21224 ;
    wire new_AGEMA_signal_21225 ;
    wire new_AGEMA_signal_21226 ;
    wire new_AGEMA_signal_21227 ;
    wire new_AGEMA_signal_21228 ;
    wire new_AGEMA_signal_21229 ;
    wire new_AGEMA_signal_21230 ;
    wire new_AGEMA_signal_21231 ;
    wire new_AGEMA_signal_21232 ;
    wire new_AGEMA_signal_21233 ;
    wire new_AGEMA_signal_21234 ;
    wire new_AGEMA_signal_21235 ;
    wire new_AGEMA_signal_21239 ;
    wire new_AGEMA_signal_21240 ;
    wire new_AGEMA_signal_21241 ;
    wire new_AGEMA_signal_21251 ;
    wire new_AGEMA_signal_21252 ;
    wire new_AGEMA_signal_21253 ;
    wire new_AGEMA_signal_21254 ;
    wire new_AGEMA_signal_21255 ;
    wire new_AGEMA_signal_21256 ;
    wire new_AGEMA_signal_21257 ;
    wire new_AGEMA_signal_21258 ;
    wire new_AGEMA_signal_21259 ;
    wire new_AGEMA_signal_21260 ;
    wire new_AGEMA_signal_21261 ;
    wire new_AGEMA_signal_21262 ;
    wire new_AGEMA_signal_21263 ;
    wire new_AGEMA_signal_21264 ;
    wire new_AGEMA_signal_21265 ;
    wire new_AGEMA_signal_21266 ;
    wire new_AGEMA_signal_21267 ;
    wire new_AGEMA_signal_21268 ;
    wire new_AGEMA_signal_21272 ;
    wire new_AGEMA_signal_21273 ;
    wire new_AGEMA_signal_21274 ;
    wire new_AGEMA_signal_21275 ;
    wire new_AGEMA_signal_21276 ;
    wire new_AGEMA_signal_21277 ;
    wire new_AGEMA_signal_21281 ;
    wire new_AGEMA_signal_21282 ;
    wire new_AGEMA_signal_21283 ;
    wire new_AGEMA_signal_21284 ;
    wire new_AGEMA_signal_21285 ;
    wire new_AGEMA_signal_21286 ;
    wire new_AGEMA_signal_21287 ;
    wire new_AGEMA_signal_21288 ;
    wire new_AGEMA_signal_21289 ;
    wire new_AGEMA_signal_21290 ;
    wire new_AGEMA_signal_21291 ;
    wire new_AGEMA_signal_21292 ;
    wire new_AGEMA_signal_21293 ;
    wire new_AGEMA_signal_21294 ;
    wire new_AGEMA_signal_21295 ;
    wire new_AGEMA_signal_21305 ;
    wire new_AGEMA_signal_21306 ;
    wire new_AGEMA_signal_21307 ;
    wire new_AGEMA_signal_21308 ;
    wire new_AGEMA_signal_21309 ;
    wire new_AGEMA_signal_21310 ;
    wire new_AGEMA_signal_21311 ;
    wire new_AGEMA_signal_21312 ;
    wire new_AGEMA_signal_21313 ;
    wire new_AGEMA_signal_21314 ;
    wire new_AGEMA_signal_21315 ;
    wire new_AGEMA_signal_21316 ;
    wire new_AGEMA_signal_21326 ;
    wire new_AGEMA_signal_21327 ;
    wire new_AGEMA_signal_21328 ;
    wire new_AGEMA_signal_21332 ;
    wire new_AGEMA_signal_21333 ;
    wire new_AGEMA_signal_21334 ;
    wire new_AGEMA_signal_21335 ;
    wire new_AGEMA_signal_21336 ;
    wire new_AGEMA_signal_21337 ;
    wire new_AGEMA_signal_21338 ;
    wire new_AGEMA_signal_21339 ;
    wire new_AGEMA_signal_21340 ;
    wire new_AGEMA_signal_21341 ;
    wire new_AGEMA_signal_21342 ;
    wire new_AGEMA_signal_21343 ;
    wire new_AGEMA_signal_21344 ;
    wire new_AGEMA_signal_21345 ;
    wire new_AGEMA_signal_21346 ;
    wire new_AGEMA_signal_21404 ;
    wire new_AGEMA_signal_21405 ;
    wire new_AGEMA_signal_21406 ;
    wire new_AGEMA_signal_21407 ;
    wire new_AGEMA_signal_21408 ;
    wire new_AGEMA_signal_21409 ;
    wire new_AGEMA_signal_21410 ;
    wire new_AGEMA_signal_21411 ;
    wire new_AGEMA_signal_21412 ;
    wire new_AGEMA_signal_21413 ;
    wire new_AGEMA_signal_21414 ;
    wire new_AGEMA_signal_21415 ;
    wire new_AGEMA_signal_21416 ;
    wire new_AGEMA_signal_21417 ;
    wire new_AGEMA_signal_21418 ;
    wire new_AGEMA_signal_21419 ;
    wire new_AGEMA_signal_21420 ;
    wire new_AGEMA_signal_21421 ;
    wire new_AGEMA_signal_21422 ;
    wire new_AGEMA_signal_21423 ;
    wire new_AGEMA_signal_21424 ;
    wire new_AGEMA_signal_21425 ;
    wire new_AGEMA_signal_21426 ;
    wire new_AGEMA_signal_21427 ;
    wire new_AGEMA_signal_21428 ;
    wire new_AGEMA_signal_21429 ;
    wire new_AGEMA_signal_21430 ;
    wire new_AGEMA_signal_21431 ;
    wire new_AGEMA_signal_21432 ;
    wire new_AGEMA_signal_21433 ;
    wire new_AGEMA_signal_21434 ;
    wire new_AGEMA_signal_21435 ;
    wire new_AGEMA_signal_21436 ;
    wire new_AGEMA_signal_21437 ;
    wire new_AGEMA_signal_21438 ;
    wire new_AGEMA_signal_21439 ;
    wire new_AGEMA_signal_21440 ;
    wire new_AGEMA_signal_21441 ;
    wire new_AGEMA_signal_21442 ;
    wire new_AGEMA_signal_21443 ;
    wire new_AGEMA_signal_21444 ;
    wire new_AGEMA_signal_21445 ;
    wire new_AGEMA_signal_21446 ;
    wire new_AGEMA_signal_21447 ;
    wire new_AGEMA_signal_21448 ;
    wire new_AGEMA_signal_21449 ;
    wire new_AGEMA_signal_21450 ;
    wire new_AGEMA_signal_21451 ;
    wire new_AGEMA_signal_21452 ;
    wire new_AGEMA_signal_21453 ;
    wire new_AGEMA_signal_21454 ;
    wire new_AGEMA_signal_21455 ;
    wire new_AGEMA_signal_21456 ;
    wire new_AGEMA_signal_21457 ;
    wire new_AGEMA_signal_21458 ;
    wire new_AGEMA_signal_21459 ;
    wire new_AGEMA_signal_21460 ;
    wire new_AGEMA_signal_21461 ;
    wire new_AGEMA_signal_21462 ;
    wire new_AGEMA_signal_21463 ;
    wire new_AGEMA_signal_21464 ;
    wire new_AGEMA_signal_21465 ;
    wire new_AGEMA_signal_21466 ;
    wire new_AGEMA_signal_21467 ;
    wire new_AGEMA_signal_21468 ;
    wire new_AGEMA_signal_21469 ;
    wire new_AGEMA_signal_21470 ;
    wire new_AGEMA_signal_21471 ;
    wire new_AGEMA_signal_21472 ;
    wire new_AGEMA_signal_21473 ;
    wire new_AGEMA_signal_21474 ;
    wire new_AGEMA_signal_21475 ;
    wire new_AGEMA_signal_21476 ;
    wire new_AGEMA_signal_21477 ;
    wire new_AGEMA_signal_21478 ;
    wire new_AGEMA_signal_21479 ;
    wire new_AGEMA_signal_21480 ;
    wire new_AGEMA_signal_21481 ;
    wire new_AGEMA_signal_21482 ;
    wire new_AGEMA_signal_21483 ;
    wire new_AGEMA_signal_21484 ;
    wire new_AGEMA_signal_21485 ;
    wire new_AGEMA_signal_21486 ;
    wire new_AGEMA_signal_21487 ;
    wire new_AGEMA_signal_21488 ;
    wire new_AGEMA_signal_21489 ;
    wire new_AGEMA_signal_21490 ;
    wire new_AGEMA_signal_21491 ;
    wire new_AGEMA_signal_21492 ;
    wire new_AGEMA_signal_21493 ;
    wire new_AGEMA_signal_21494 ;
    wire new_AGEMA_signal_21495 ;
    wire new_AGEMA_signal_21496 ;
    wire new_AGEMA_signal_21497 ;
    wire new_AGEMA_signal_21498 ;
    wire new_AGEMA_signal_21499 ;
    wire new_AGEMA_signal_21500 ;
    wire new_AGEMA_signal_21501 ;
    wire new_AGEMA_signal_21502 ;
    wire new_AGEMA_signal_21503 ;
    wire new_AGEMA_signal_21504 ;
    wire new_AGEMA_signal_21505 ;
    wire new_AGEMA_signal_21506 ;
    wire new_AGEMA_signal_21507 ;
    wire new_AGEMA_signal_21508 ;
    wire new_AGEMA_signal_21509 ;
    wire new_AGEMA_signal_21510 ;
    wire new_AGEMA_signal_21511 ;
    wire new_AGEMA_signal_21677 ;
    wire new_AGEMA_signal_21678 ;
    wire new_AGEMA_signal_21679 ;
    wire new_AGEMA_signal_21680 ;
    wire new_AGEMA_signal_21681 ;
    wire new_AGEMA_signal_21682 ;
    wire new_AGEMA_signal_21683 ;
    wire new_AGEMA_signal_21684 ;
    wire new_AGEMA_signal_21685 ;
    wire new_AGEMA_signal_21695 ;
    wire new_AGEMA_signal_21696 ;
    wire new_AGEMA_signal_21697 ;
    wire new_AGEMA_signal_21698 ;
    wire new_AGEMA_signal_21699 ;
    wire new_AGEMA_signal_21700 ;
    wire new_AGEMA_signal_21701 ;
    wire new_AGEMA_signal_21702 ;
    wire new_AGEMA_signal_21703 ;
    wire new_AGEMA_signal_21788 ;
    wire new_AGEMA_signal_21789 ;
    wire new_AGEMA_signal_21790 ;
    wire new_AGEMA_signal_21791 ;
    wire new_AGEMA_signal_21792 ;
    wire new_AGEMA_signal_21793 ;
    wire new_AGEMA_signal_21830 ;
    wire new_AGEMA_signal_21831 ;
    wire new_AGEMA_signal_21832 ;
    wire new_AGEMA_signal_21836 ;
    wire new_AGEMA_signal_21837 ;
    wire new_AGEMA_signal_21838 ;
    wire new_AGEMA_signal_21950 ;
    wire new_AGEMA_signal_21951 ;
    wire new_AGEMA_signal_21952 ;
    wire new_AGEMA_signal_21953 ;
    wire new_AGEMA_signal_21954 ;
    wire new_AGEMA_signal_21955 ;
    wire clk_gated ;

    /* cells in depth 0 */
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_0_U1 ( .s (p256_sel), .b ({w0_s3[0], w0_s2[0], w0_s1[0], w0_s0[0]}), .a ({w1_s3[0], w1_s2[0], w1_s1[0], w1_s0[0]}), .c ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, new_AGEMA_signal_5738, addc_in[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_1_U1 ( .s (p256_sel), .b ({w0_s3[1], w0_s2[1], w0_s1[1], w0_s0[1]}), .a ({w1_s3[1], w1_s2[1], w1_s1[1], w1_s0[1]}), .c ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, new_AGEMA_signal_5747, addc_in[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_2_U1 ( .s (p256_sel), .b ({w0_s3[2], w0_s2[2], w0_s1[2], w0_s0[2]}), .a ({w1_s3[2], w1_s2[2], w1_s1[2], w1_s0[2]}), .c ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, new_AGEMA_signal_5756, addc_in[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_3_U1 ( .s (p256_sel), .b ({w0_s3[3], w0_s2[3], w0_s1[3], w0_s0[3]}), .a ({w1_s3[3], w1_s2[3], w1_s1[3], w1_s0[3]}), .c ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, new_AGEMA_signal_5765, addc_in[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_4_U1 ( .s (p256_sel), .b ({w0_s3[4], w0_s2[4], w0_s1[4], w0_s0[4]}), .a ({w1_s3[4], w1_s2[4], w1_s1[4], w1_s0[4]}), .c ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, new_AGEMA_signal_5774, addc_in[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_5_U1 ( .s (p256_sel), .b ({w0_s3[5], w0_s2[5], w0_s1[5], w0_s0[5]}), .a ({w1_s3[5], w1_s2[5], w1_s1[5], w1_s0[5]}), .c ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, new_AGEMA_signal_5783, addc_in[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_6_U1 ( .s (p256_sel), .b ({w0_s3[6], w0_s2[6], w0_s1[6], w0_s0[6]}), .a ({w1_s3[6], w1_s2[6], w1_s1[6], w1_s0[6]}), .c ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, new_AGEMA_signal_5792, addc_in[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_7_U1 ( .s (p256_sel), .b ({w0_s3[7], w0_s2[7], w0_s1[7], w0_s0[7]}), .a ({w1_s3[7], w1_s2[7], w1_s1[7], w1_s0[7]}), .c ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, new_AGEMA_signal_5801, addc_in[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_8_U1 ( .s (p256_sel), .b ({w0_s3[8], w0_s2[8], w0_s1[8], w0_s0[8]}), .a ({w1_s3[8], w1_s2[8], w1_s1[8], w1_s0[8]}), .c ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, new_AGEMA_signal_5810, addc_in[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_9_U1 ( .s (p256_sel), .b ({w0_s3[9], w0_s2[9], w0_s1[9], w0_s0[9]}), .a ({w1_s3[9], w1_s2[9], w1_s1[9], w1_s0[9]}), .c ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, new_AGEMA_signal_5819, addc_in[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_10_U1 ( .s (p256_sel), .b ({w0_s3[10], w0_s2[10], w0_s1[10], w0_s0[10]}), .a ({w1_s3[10], w1_s2[10], w1_s1[10], w1_s0[10]}), .c ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, new_AGEMA_signal_5828, addc_in[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_11_U1 ( .s (p256_sel), .b ({w0_s3[11], w0_s2[11], w0_s1[11], w0_s0[11]}), .a ({w1_s3[11], w1_s2[11], w1_s1[11], w1_s0[11]}), .c ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, new_AGEMA_signal_5837, addc_in[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_12_U1 ( .s (p256_sel), .b ({w0_s3[12], w0_s2[12], w0_s1[12], w0_s0[12]}), .a ({w1_s3[12], w1_s2[12], w1_s1[12], w1_s0[12]}), .c ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, new_AGEMA_signal_5846, addc_in[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_13_U1 ( .s (p256_sel), .b ({w0_s3[13], w0_s2[13], w0_s1[13], w0_s0[13]}), .a ({w1_s3[13], w1_s2[13], w1_s1[13], w1_s0[13]}), .c ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, new_AGEMA_signal_5855, addc_in[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_14_U1 ( .s (p256_sel), .b ({w0_s3[14], w0_s2[14], w0_s1[14], w0_s0[14]}), .a ({w1_s3[14], w1_s2[14], w1_s1[14], w1_s0[14]}), .c ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, new_AGEMA_signal_5864, addc_in[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_15_U1 ( .s (p256_sel), .b ({w0_s3[15], w0_s2[15], w0_s1[15], w0_s0[15]}), .a ({w1_s3[15], w1_s2[15], w1_s1[15], w1_s0[15]}), .c ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, new_AGEMA_signal_5873, addc_in[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_16_U1 ( .s (p256_sel), .b ({w0_s3[16], w0_s2[16], w0_s1[16], w0_s0[16]}), .a ({w1_s3[16], w1_s2[16], w1_s1[16], w1_s0[16]}), .c ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, new_AGEMA_signal_5882, addc_in[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_17_U1 ( .s (p256_sel), .b ({w0_s3[17], w0_s2[17], w0_s1[17], w0_s0[17]}), .a ({w1_s3[17], w1_s2[17], w1_s1[17], w1_s0[17]}), .c ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, new_AGEMA_signal_5891, addc_in[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_18_U1 ( .s (p256_sel), .b ({w0_s3[18], w0_s2[18], w0_s1[18], w0_s0[18]}), .a ({w1_s3[18], w1_s2[18], w1_s1[18], w1_s0[18]}), .c ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, new_AGEMA_signal_5900, addc_in[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_19_U1 ( .s (p256_sel), .b ({w0_s3[19], w0_s2[19], w0_s1[19], w0_s0[19]}), .a ({w1_s3[19], w1_s2[19], w1_s1[19], w1_s0[19]}), .c ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, new_AGEMA_signal_5909, addc_in[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_20_U1 ( .s (p256_sel), .b ({w0_s3[20], w0_s2[20], w0_s1[20], w0_s0[20]}), .a ({w1_s3[20], w1_s2[20], w1_s1[20], w1_s0[20]}), .c ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, new_AGEMA_signal_5918, addc_in[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_21_U1 ( .s (p256_sel), .b ({w0_s3[21], w0_s2[21], w0_s1[21], w0_s0[21]}), .a ({w1_s3[21], w1_s2[21], w1_s1[21], w1_s0[21]}), .c ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, new_AGEMA_signal_5927, addc_in[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_22_U1 ( .s (p256_sel), .b ({w0_s3[22], w0_s2[22], w0_s1[22], w0_s0[22]}), .a ({w1_s3[22], w1_s2[22], w1_s1[22], w1_s0[22]}), .c ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, new_AGEMA_signal_5936, addc_in[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_23_U1 ( .s (p256_sel), .b ({w0_s3[23], w0_s2[23], w0_s1[23], w0_s0[23]}), .a ({w1_s3[23], w1_s2[23], w1_s1[23], w1_s0[23]}), .c ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, new_AGEMA_signal_5945, addc_in[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_24_U1 ( .s (p256_sel), .b ({w0_s3[24], w0_s2[24], w0_s1[24], w0_s0[24]}), .a ({w1_s3[24], w1_s2[24], w1_s1[24], w1_s0[24]}), .c ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, new_AGEMA_signal_5954, addc_in[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_25_U1 ( .s (p256_sel), .b ({w0_s3[25], w0_s2[25], w0_s1[25], w0_s0[25]}), .a ({w1_s3[25], w1_s2[25], w1_s1[25], w1_s0[25]}), .c ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, new_AGEMA_signal_5963, addc_in[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_26_U1 ( .s (p256_sel), .b ({w0_s3[26], w0_s2[26], w0_s1[26], w0_s0[26]}), .a ({w1_s3[26], w1_s2[26], w1_s1[26], w1_s0[26]}), .c ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, new_AGEMA_signal_5972, addc_in[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_27_U1 ( .s (p256_sel), .b ({w0_s3[27], w0_s2[27], w0_s1[27], w0_s0[27]}), .a ({w1_s3[27], w1_s2[27], w1_s1[27], w1_s0[27]}), .c ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, new_AGEMA_signal_5981, addc_in[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_28_U1 ( .s (p256_sel), .b ({w0_s3[28], w0_s2[28], w0_s1[28], w0_s0[28]}), .a ({w1_s3[28], w1_s2[28], w1_s1[28], w1_s0[28]}), .c ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, new_AGEMA_signal_5990, addc_in[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_29_U1 ( .s (p256_sel), .b ({w0_s3[29], w0_s2[29], w0_s1[29], w0_s0[29]}), .a ({w1_s3[29], w1_s2[29], w1_s1[29], w1_s0[29]}), .c ({new_AGEMA_signal_6001, new_AGEMA_signal_6000, new_AGEMA_signal_5999, addc_in[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_30_U1 ( .s (p256_sel), .b ({w0_s3[30], w0_s2[30], w0_s1[30], w0_s0[30]}), .a ({w1_s3[30], w1_s2[30], w1_s1[30], w1_s0[30]}), .c ({new_AGEMA_signal_6010, new_AGEMA_signal_6009, new_AGEMA_signal_6008, addc_in[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_31_U1 ( .s (p256_sel), .b ({w0_s3[31], w0_s2[31], w0_s1[31], w0_s0[31]}), .a ({w1_s3[31], w1_s2[31], w1_s1[31], w1_s0[31]}), .c ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, new_AGEMA_signal_6017, addc_in[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_32_U1 ( .s (p256_sel), .b ({w0_s3[32], w0_s2[32], w0_s1[32], w0_s0[32]}), .a ({w1_s3[32], w1_s2[32], w1_s1[32], w1_s0[32]}), .c ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, new_AGEMA_signal_6026, addc_in[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_33_U1 ( .s (p256_sel), .b ({w0_s3[33], w0_s2[33], w0_s1[33], w0_s0[33]}), .a ({w1_s3[33], w1_s2[33], w1_s1[33], w1_s0[33]}), .c ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, new_AGEMA_signal_6035, addc_in[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_34_U1 ( .s (p256_sel), .b ({w0_s3[34], w0_s2[34], w0_s1[34], w0_s0[34]}), .a ({w1_s3[34], w1_s2[34], w1_s1[34], w1_s0[34]}), .c ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, new_AGEMA_signal_6044, addc_in[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_35_U1 ( .s (p256_sel), .b ({w0_s3[35], w0_s2[35], w0_s1[35], w0_s0[35]}), .a ({w1_s3[35], w1_s2[35], w1_s1[35], w1_s0[35]}), .c ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, new_AGEMA_signal_6053, addc_in[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_36_U1 ( .s (p256_sel), .b ({w0_s3[36], w0_s2[36], w0_s1[36], w0_s0[36]}), .a ({w1_s3[36], w1_s2[36], w1_s1[36], w1_s0[36]}), .c ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, new_AGEMA_signal_6062, addc_in[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_37_U1 ( .s (p256_sel), .b ({w0_s3[37], w0_s2[37], w0_s1[37], w0_s0[37]}), .a ({w1_s3[37], w1_s2[37], w1_s1[37], w1_s0[37]}), .c ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, new_AGEMA_signal_6071, addc_in[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_38_U1 ( .s (p256_sel), .b ({w0_s3[38], w0_s2[38], w0_s1[38], w0_s0[38]}), .a ({w1_s3[38], w1_s2[38], w1_s1[38], w1_s0[38]}), .c ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, new_AGEMA_signal_6080, addc_in[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_39_U1 ( .s (p256_sel), .b ({w0_s3[39], w0_s2[39], w0_s1[39], w0_s0[39]}), .a ({w1_s3[39], w1_s2[39], w1_s1[39], w1_s0[39]}), .c ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, new_AGEMA_signal_6089, addc_in[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_40_U1 ( .s (p256_sel), .b ({w0_s3[40], w0_s2[40], w0_s1[40], w0_s0[40]}), .a ({w1_s3[40], w1_s2[40], w1_s1[40], w1_s0[40]}), .c ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, new_AGEMA_signal_6098, addc_in[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_41_U1 ( .s (p256_sel), .b ({w0_s3[41], w0_s2[41], w0_s1[41], w0_s0[41]}), .a ({w1_s3[41], w1_s2[41], w1_s1[41], w1_s0[41]}), .c ({new_AGEMA_signal_6109, new_AGEMA_signal_6108, new_AGEMA_signal_6107, addc_in[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_42_U1 ( .s (p256_sel), .b ({w0_s3[42], w0_s2[42], w0_s1[42], w0_s0[42]}), .a ({w1_s3[42], w1_s2[42], w1_s1[42], w1_s0[42]}), .c ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, new_AGEMA_signal_6116, addc_in[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_43_U1 ( .s (p256_sel), .b ({w0_s3[43], w0_s2[43], w0_s1[43], w0_s0[43]}), .a ({w1_s3[43], w1_s2[43], w1_s1[43], w1_s0[43]}), .c ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, new_AGEMA_signal_6125, addc_in[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_44_U1 ( .s (p256_sel), .b ({w0_s3[44], w0_s2[44], w0_s1[44], w0_s0[44]}), .a ({w1_s3[44], w1_s2[44], w1_s1[44], w1_s0[44]}), .c ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, new_AGEMA_signal_6134, addc_in[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_45_U1 ( .s (p256_sel), .b ({w0_s3[45], w0_s2[45], w0_s1[45], w0_s0[45]}), .a ({w1_s3[45], w1_s2[45], w1_s1[45], w1_s0[45]}), .c ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, new_AGEMA_signal_6143, addc_in[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_46_U1 ( .s (p256_sel), .b ({w0_s3[46], w0_s2[46], w0_s1[46], w0_s0[46]}), .a ({w1_s3[46], w1_s2[46], w1_s1[46], w1_s0[46]}), .c ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, new_AGEMA_signal_6152, addc_in[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_47_U1 ( .s (p256_sel), .b ({w0_s3[47], w0_s2[47], w0_s1[47], w0_s0[47]}), .a ({w1_s3[47], w1_s2[47], w1_s1[47], w1_s0[47]}), .c ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, new_AGEMA_signal_6161, addc_in[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_48_U1 ( .s (p256_sel), .b ({w0_s3[48], w0_s2[48], w0_s1[48], w0_s0[48]}), .a ({w1_s3[48], w1_s2[48], w1_s1[48], w1_s0[48]}), .c ({new_AGEMA_signal_6172, new_AGEMA_signal_6171, new_AGEMA_signal_6170, addc_in[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_49_U1 ( .s (p256_sel), .b ({w0_s3[49], w0_s2[49], w0_s1[49], w0_s0[49]}), .a ({w1_s3[49], w1_s2[49], w1_s1[49], w1_s0[49]}), .c ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, new_AGEMA_signal_6179, addc_in[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_50_U1 ( .s (p256_sel), .b ({w0_s3[50], w0_s2[50], w0_s1[50], w0_s0[50]}), .a ({w1_s3[50], w1_s2[50], w1_s1[50], w1_s0[50]}), .c ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, addc_in[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_51_U1 ( .s (p256_sel), .b ({w0_s3[51], w0_s2[51], w0_s1[51], w0_s0[51]}), .a ({w1_s3[51], w1_s2[51], w1_s1[51], w1_s0[51]}), .c ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, new_AGEMA_signal_6197, addc_in[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_52_U1 ( .s (p256_sel), .b ({w0_s3[52], w0_s2[52], w0_s1[52], w0_s0[52]}), .a ({w1_s3[52], w1_s2[52], w1_s1[52], w1_s0[52]}), .c ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, new_AGEMA_signal_6206, addc_in[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_53_U1 ( .s (p256_sel), .b ({w0_s3[53], w0_s2[53], w0_s1[53], w0_s0[53]}), .a ({w1_s3[53], w1_s2[53], w1_s1[53], w1_s0[53]}), .c ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, new_AGEMA_signal_6215, addc_in[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_54_U1 ( .s (p256_sel), .b ({w0_s3[54], w0_s2[54], w0_s1[54], w0_s0[54]}), .a ({w1_s3[54], w1_s2[54], w1_s1[54], w1_s0[54]}), .c ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, new_AGEMA_signal_6224, addc_in[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_55_U1 ( .s (p256_sel), .b ({w0_s3[55], w0_s2[55], w0_s1[55], w0_s0[55]}), .a ({w1_s3[55], w1_s2[55], w1_s1[55], w1_s0[55]}), .c ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, addc_in[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_56_U1 ( .s (p256_sel), .b ({w0_s3[56], w0_s2[56], w0_s1[56], w0_s0[56]}), .a ({w1_s3[56], w1_s2[56], w1_s1[56], w1_s0[56]}), .c ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, new_AGEMA_signal_6242, addc_in[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_57_U1 ( .s (p256_sel), .b ({w0_s3[57], w0_s2[57], w0_s1[57], w0_s0[57]}), .a ({w1_s3[57], w1_s2[57], w1_s1[57], w1_s0[57]}), .c ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, new_AGEMA_signal_6251, addc_in[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_58_U1 ( .s (p256_sel), .b ({w0_s3[58], w0_s2[58], w0_s1[58], w0_s0[58]}), .a ({w1_s3[58], w1_s2[58], w1_s1[58], w1_s0[58]}), .c ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, new_AGEMA_signal_6260, addc_in[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_59_U1 ( .s (p256_sel), .b ({w0_s3[59], w0_s2[59], w0_s1[59], w0_s0[59]}), .a ({w1_s3[59], w1_s2[59], w1_s1[59], w1_s0[59]}), .c ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, new_AGEMA_signal_6269, addc_in[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_60_U1 ( .s (p256_sel), .b ({w0_s3[60], w0_s2[60], w0_s1[60], w0_s0[60]}), .a ({w1_s3[60], w1_s2[60], w1_s1[60], w1_s0[60]}), .c ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, new_AGEMA_signal_6278, addc_in[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_61_U1 ( .s (p256_sel), .b ({w0_s3[61], w0_s2[61], w0_s1[61], w0_s0[61]}), .a ({w1_s3[61], w1_s2[61], w1_s1[61], w1_s0[61]}), .c ({new_AGEMA_signal_6289, new_AGEMA_signal_6288, new_AGEMA_signal_6287, addc_in[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_62_U1 ( .s (p256_sel), .b ({w0_s3[62], w0_s2[62], w0_s1[62], w0_s0[62]}), .a ({w1_s3[62], w1_s2[62], w1_s1[62], w1_s0[62]}), .c ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, new_AGEMA_signal_6296, addc_in[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_63_U1 ( .s (p256_sel), .b ({w0_s3[63], w0_s2[63], w0_s1[63], w0_s0[63]}), .a ({w1_s3[63], w1_s2[63], w1_s1[63], w1_s0[63]}), .c ({new_AGEMA_signal_6307, new_AGEMA_signal_6306, new_AGEMA_signal_6305, addc_in[63]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_64_U1 ( .s (p256_sel), .b ({w0_s3[64], w0_s2[64], w0_s1[64], w0_s0[64]}), .a ({w1_s3[64], w1_s2[64], w1_s1[64], w1_s0[64]}), .c ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, new_AGEMA_signal_6314, addc_in[64]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_65_U1 ( .s (p256_sel), .b ({w0_s3[65], w0_s2[65], w0_s1[65], w0_s0[65]}), .a ({w1_s3[65], w1_s2[65], w1_s1[65], w1_s0[65]}), .c ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, new_AGEMA_signal_6323, addc_in[65]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_66_U1 ( .s (p256_sel), .b ({w0_s3[66], w0_s2[66], w0_s1[66], w0_s0[66]}), .a ({w1_s3[66], w1_s2[66], w1_s1[66], w1_s0[66]}), .c ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, new_AGEMA_signal_6332, addc_in[66]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_67_U1 ( .s (p256_sel), .b ({w0_s3[67], w0_s2[67], w0_s1[67], w0_s0[67]}), .a ({w1_s3[67], w1_s2[67], w1_s1[67], w1_s0[67]}), .c ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, new_AGEMA_signal_6341, addc_in[67]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_68_U1 ( .s (p256_sel), .b ({w0_s3[68], w0_s2[68], w0_s1[68], w0_s0[68]}), .a ({w1_s3[68], w1_s2[68], w1_s1[68], w1_s0[68]}), .c ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, new_AGEMA_signal_6350, addc_in[68]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_69_U1 ( .s (p256_sel), .b ({w0_s3[69], w0_s2[69], w0_s1[69], w0_s0[69]}), .a ({w1_s3[69], w1_s2[69], w1_s1[69], w1_s0[69]}), .c ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, new_AGEMA_signal_6359, addc_in[69]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_70_U1 ( .s (p256_sel), .b ({w0_s3[70], w0_s2[70], w0_s1[70], w0_s0[70]}), .a ({w1_s3[70], w1_s2[70], w1_s1[70], w1_s0[70]}), .c ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, new_AGEMA_signal_6368, addc_in[70]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_71_U1 ( .s (p256_sel), .b ({w0_s3[71], w0_s2[71], w0_s1[71], w0_s0[71]}), .a ({w1_s3[71], w1_s2[71], w1_s1[71], w1_s0[71]}), .c ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, new_AGEMA_signal_6377, addc_in[71]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_72_U1 ( .s (p256_sel), .b ({w0_s3[72], w0_s2[72], w0_s1[72], w0_s0[72]}), .a ({w1_s3[72], w1_s2[72], w1_s1[72], w1_s0[72]}), .c ({new_AGEMA_signal_6388, new_AGEMA_signal_6387, new_AGEMA_signal_6386, addc_in[72]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_73_U1 ( .s (p256_sel), .b ({w0_s3[73], w0_s2[73], w0_s1[73], w0_s0[73]}), .a ({w1_s3[73], w1_s2[73], w1_s1[73], w1_s0[73]}), .c ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, new_AGEMA_signal_6395, addc_in[73]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_74_U1 ( .s (p256_sel), .b ({w0_s3[74], w0_s2[74], w0_s1[74], w0_s0[74]}), .a ({w1_s3[74], w1_s2[74], w1_s1[74], w1_s0[74]}), .c ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, new_AGEMA_signal_6404, addc_in[74]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_75_U1 ( .s (p256_sel), .b ({w0_s3[75], w0_s2[75], w0_s1[75], w0_s0[75]}), .a ({w1_s3[75], w1_s2[75], w1_s1[75], w1_s0[75]}), .c ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, new_AGEMA_signal_6413, addc_in[75]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_76_U1 ( .s (p256_sel), .b ({w0_s3[76], w0_s2[76], w0_s1[76], w0_s0[76]}), .a ({w1_s3[76], w1_s2[76], w1_s1[76], w1_s0[76]}), .c ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, new_AGEMA_signal_6422, addc_in[76]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_77_U1 ( .s (p256_sel), .b ({w0_s3[77], w0_s2[77], w0_s1[77], w0_s0[77]}), .a ({w1_s3[77], w1_s2[77], w1_s1[77], w1_s0[77]}), .c ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, new_AGEMA_signal_6431, addc_in[77]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_78_U1 ( .s (p256_sel), .b ({w0_s3[78], w0_s2[78], w0_s1[78], w0_s0[78]}), .a ({w1_s3[78], w1_s2[78], w1_s1[78], w1_s0[78]}), .c ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, new_AGEMA_signal_6440, addc_in[78]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_79_U1 ( .s (p256_sel), .b ({w0_s3[79], w0_s2[79], w0_s1[79], w0_s0[79]}), .a ({w1_s3[79], w1_s2[79], w1_s1[79], w1_s0[79]}), .c ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, new_AGEMA_signal_6449, addc_in[79]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_80_U1 ( .s (p256_sel), .b ({w0_s3[80], w0_s2[80], w0_s1[80], w0_s0[80]}), .a ({w1_s3[80], w1_s2[80], w1_s1[80], w1_s0[80]}), .c ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, new_AGEMA_signal_6458, addc_in[80]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_81_U1 ( .s (p256_sel), .b ({w0_s3[81], w0_s2[81], w0_s1[81], w0_s0[81]}), .a ({w1_s3[81], w1_s2[81], w1_s1[81], w1_s0[81]}), .c ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, new_AGEMA_signal_6467, addc_in[81]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_82_U1 ( .s (p256_sel), .b ({w0_s3[82], w0_s2[82], w0_s1[82], w0_s0[82]}), .a ({w1_s3[82], w1_s2[82], w1_s1[82], w1_s0[82]}), .c ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, new_AGEMA_signal_6476, addc_in[82]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_83_U1 ( .s (p256_sel), .b ({w0_s3[83], w0_s2[83], w0_s1[83], w0_s0[83]}), .a ({w1_s3[83], w1_s2[83], w1_s1[83], w1_s0[83]}), .c ({new_AGEMA_signal_6487, new_AGEMA_signal_6486, new_AGEMA_signal_6485, addc_in[83]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_84_U1 ( .s (p256_sel), .b ({w0_s3[84], w0_s2[84], w0_s1[84], w0_s0[84]}), .a ({w1_s3[84], w1_s2[84], w1_s1[84], w1_s0[84]}), .c ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, new_AGEMA_signal_6494, addc_in[84]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_85_U1 ( .s (p256_sel), .b ({w0_s3[85], w0_s2[85], w0_s1[85], w0_s0[85]}), .a ({w1_s3[85], w1_s2[85], w1_s1[85], w1_s0[85]}), .c ({new_AGEMA_signal_6505, new_AGEMA_signal_6504, new_AGEMA_signal_6503, addc_in[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_86_U1 ( .s (p256_sel), .b ({w0_s3[86], w0_s2[86], w0_s1[86], w0_s0[86]}), .a ({w1_s3[86], w1_s2[86], w1_s1[86], w1_s0[86]}), .c ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, new_AGEMA_signal_6512, addc_in[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_87_U1 ( .s (p256_sel), .b ({w0_s3[87], w0_s2[87], w0_s1[87], w0_s0[87]}), .a ({w1_s3[87], w1_s2[87], w1_s1[87], w1_s0[87]}), .c ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, new_AGEMA_signal_6521, addc_in[87]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_88_U1 ( .s (p256_sel), .b ({w0_s3[88], w0_s2[88], w0_s1[88], w0_s0[88]}), .a ({w1_s3[88], w1_s2[88], w1_s1[88], w1_s0[88]}), .c ({new_AGEMA_signal_6532, new_AGEMA_signal_6531, new_AGEMA_signal_6530, addc_in[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_89_U1 ( .s (p256_sel), .b ({w0_s3[89], w0_s2[89], w0_s1[89], w0_s0[89]}), .a ({w1_s3[89], w1_s2[89], w1_s1[89], w1_s0[89]}), .c ({new_AGEMA_signal_6541, new_AGEMA_signal_6540, new_AGEMA_signal_6539, addc_in[89]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_90_U1 ( .s (p256_sel), .b ({w0_s3[90], w0_s2[90], w0_s1[90], w0_s0[90]}), .a ({w1_s3[90], w1_s2[90], w1_s1[90], w1_s0[90]}), .c ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, new_AGEMA_signal_6548, addc_in[90]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_91_U1 ( .s (p256_sel), .b ({w0_s3[91], w0_s2[91], w0_s1[91], w0_s0[91]}), .a ({w1_s3[91], w1_s2[91], w1_s1[91], w1_s0[91]}), .c ({new_AGEMA_signal_6559, new_AGEMA_signal_6558, new_AGEMA_signal_6557, addc_in[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_92_U1 ( .s (p256_sel), .b ({w0_s3[92], w0_s2[92], w0_s1[92], w0_s0[92]}), .a ({w1_s3[92], w1_s2[92], w1_s1[92], w1_s0[92]}), .c ({new_AGEMA_signal_6568, new_AGEMA_signal_6567, new_AGEMA_signal_6566, addc_in[92]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_93_U1 ( .s (p256_sel), .b ({w0_s3[93], w0_s2[93], w0_s1[93], w0_s0[93]}), .a ({w1_s3[93], w1_s2[93], w1_s1[93], w1_s0[93]}), .c ({new_AGEMA_signal_6577, new_AGEMA_signal_6576, new_AGEMA_signal_6575, addc_in[93]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_94_U1 ( .s (p256_sel), .b ({w0_s3[94], w0_s2[94], w0_s1[94], w0_s0[94]}), .a ({w1_s3[94], w1_s2[94], w1_s1[94], w1_s0[94]}), .c ({new_AGEMA_signal_6586, new_AGEMA_signal_6585, new_AGEMA_signal_6584, addc_in[94]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_95_U1 ( .s (p256_sel), .b ({w0_s3[95], w0_s2[95], w0_s1[95], w0_s0[95]}), .a ({w1_s3[95], w1_s2[95], w1_s1[95], w1_s0[95]}), .c ({new_AGEMA_signal_6595, new_AGEMA_signal_6594, new_AGEMA_signal_6593, addc_in[95]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_96_U1 ( .s (p256_sel), .b ({w0_s3[96], w0_s2[96], w0_s1[96], w0_s0[96]}), .a ({w1_s3[96], w1_s2[96], w1_s1[96], w1_s0[96]}), .c ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, new_AGEMA_signal_6602, addc_in[96]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_97_U1 ( .s (p256_sel), .b ({w0_s3[97], w0_s2[97], w0_s1[97], w0_s0[97]}), .a ({w1_s3[97], w1_s2[97], w1_s1[97], w1_s0[97]}), .c ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, new_AGEMA_signal_6611, addc_in[97]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_98_U1 ( .s (p256_sel), .b ({w0_s3[98], w0_s2[98], w0_s1[98], w0_s0[98]}), .a ({w1_s3[98], w1_s2[98], w1_s1[98], w1_s0[98]}), .c ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, new_AGEMA_signal_6620, addc_in[98]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_99_U1 ( .s (p256_sel), .b ({w0_s3[99], w0_s2[99], w0_s1[99], w0_s0[99]}), .a ({w1_s3[99], w1_s2[99], w1_s1[99], w1_s0[99]}), .c ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, new_AGEMA_signal_6629, addc_in[99]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_100_U1 ( .s (p256_sel), .b ({w0_s3[100], w0_s2[100], w0_s1[100], w0_s0[100]}), .a ({w1_s3[100], w1_s2[100], w1_s1[100], w1_s0[100]}), .c ({new_AGEMA_signal_6640, new_AGEMA_signal_6639, new_AGEMA_signal_6638, addc_in[100]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_101_U1 ( .s (p256_sel), .b ({w0_s3[101], w0_s2[101], w0_s1[101], w0_s0[101]}), .a ({w1_s3[101], w1_s2[101], w1_s1[101], w1_s0[101]}), .c ({new_AGEMA_signal_6649, new_AGEMA_signal_6648, new_AGEMA_signal_6647, addc_in[101]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_102_U1 ( .s (p256_sel), .b ({w0_s3[102], w0_s2[102], w0_s1[102], w0_s0[102]}), .a ({w1_s3[102], w1_s2[102], w1_s1[102], w1_s0[102]}), .c ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, new_AGEMA_signal_6656, addc_in[102]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_103_U1 ( .s (p256_sel), .b ({w0_s3[103], w0_s2[103], w0_s1[103], w0_s0[103]}), .a ({w1_s3[103], w1_s2[103], w1_s1[103], w1_s0[103]}), .c ({new_AGEMA_signal_6667, new_AGEMA_signal_6666, new_AGEMA_signal_6665, addc_in[103]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_104_U1 ( .s (p256_sel), .b ({w0_s3[104], w0_s2[104], w0_s1[104], w0_s0[104]}), .a ({w1_s3[104], w1_s2[104], w1_s1[104], w1_s0[104]}), .c ({new_AGEMA_signal_6676, new_AGEMA_signal_6675, new_AGEMA_signal_6674, addc_in[104]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_105_U1 ( .s (p256_sel), .b ({w0_s3[105], w0_s2[105], w0_s1[105], w0_s0[105]}), .a ({w1_s3[105], w1_s2[105], w1_s1[105], w1_s0[105]}), .c ({new_AGEMA_signal_6685, new_AGEMA_signal_6684, new_AGEMA_signal_6683, addc_in[105]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_106_U1 ( .s (p256_sel), .b ({w0_s3[106], w0_s2[106], w0_s1[106], w0_s0[106]}), .a ({w1_s3[106], w1_s2[106], w1_s1[106], w1_s0[106]}), .c ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, new_AGEMA_signal_6692, addc_in[106]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_107_U1 ( .s (p256_sel), .b ({w0_s3[107], w0_s2[107], w0_s1[107], w0_s0[107]}), .a ({w1_s3[107], w1_s2[107], w1_s1[107], w1_s0[107]}), .c ({new_AGEMA_signal_6703, new_AGEMA_signal_6702, new_AGEMA_signal_6701, addc_in[107]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_108_U1 ( .s (p256_sel), .b ({w0_s3[108], w0_s2[108], w0_s1[108], w0_s0[108]}), .a ({w1_s3[108], w1_s2[108], w1_s1[108], w1_s0[108]}), .c ({new_AGEMA_signal_6712, new_AGEMA_signal_6711, new_AGEMA_signal_6710, addc_in[108]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_109_U1 ( .s (p256_sel), .b ({w0_s3[109], w0_s2[109], w0_s1[109], w0_s0[109]}), .a ({w1_s3[109], w1_s2[109], w1_s1[109], w1_s0[109]}), .c ({new_AGEMA_signal_6721, new_AGEMA_signal_6720, new_AGEMA_signal_6719, addc_in[109]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_110_U1 ( .s (p256_sel), .b ({w0_s3[110], w0_s2[110], w0_s1[110], w0_s0[110]}), .a ({w1_s3[110], w1_s2[110], w1_s1[110], w1_s0[110]}), .c ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, new_AGEMA_signal_6728, addc_in[110]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_111_U1 ( .s (p256_sel), .b ({w0_s3[111], w0_s2[111], w0_s1[111], w0_s0[111]}), .a ({w1_s3[111], w1_s2[111], w1_s1[111], w1_s0[111]}), .c ({new_AGEMA_signal_6739, new_AGEMA_signal_6738, new_AGEMA_signal_6737, addc_in[111]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_112_U1 ( .s (p256_sel), .b ({w0_s3[112], w0_s2[112], w0_s1[112], w0_s0[112]}), .a ({w1_s3[112], w1_s2[112], w1_s1[112], w1_s0[112]}), .c ({new_AGEMA_signal_6748, new_AGEMA_signal_6747, new_AGEMA_signal_6746, addc_in[112]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_113_U1 ( .s (p256_sel), .b ({w0_s3[113], w0_s2[113], w0_s1[113], w0_s0[113]}), .a ({w1_s3[113], w1_s2[113], w1_s1[113], w1_s0[113]}), .c ({new_AGEMA_signal_6757, new_AGEMA_signal_6756, new_AGEMA_signal_6755, addc_in[113]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_114_U1 ( .s (p256_sel), .b ({w0_s3[114], w0_s2[114], w0_s1[114], w0_s0[114]}), .a ({w1_s3[114], w1_s2[114], w1_s1[114], w1_s0[114]}), .c ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, new_AGEMA_signal_6764, addc_in[114]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_115_U1 ( .s (p256_sel), .b ({w0_s3[115], w0_s2[115], w0_s1[115], w0_s0[115]}), .a ({w1_s3[115], w1_s2[115], w1_s1[115], w1_s0[115]}), .c ({new_AGEMA_signal_6775, new_AGEMA_signal_6774, new_AGEMA_signal_6773, addc_in[115]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_116_U1 ( .s (p256_sel), .b ({w0_s3[116], w0_s2[116], w0_s1[116], w0_s0[116]}), .a ({w1_s3[116], w1_s2[116], w1_s1[116], w1_s0[116]}), .c ({new_AGEMA_signal_6784, new_AGEMA_signal_6783, new_AGEMA_signal_6782, addc_in[116]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_117_U1 ( .s (p256_sel), .b ({w0_s3[117], w0_s2[117], w0_s1[117], w0_s0[117]}), .a ({w1_s3[117], w1_s2[117], w1_s1[117], w1_s0[117]}), .c ({new_AGEMA_signal_6793, new_AGEMA_signal_6792, new_AGEMA_signal_6791, addc_in[117]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_118_U1 ( .s (p256_sel), .b ({w0_s3[118], w0_s2[118], w0_s1[118], w0_s0[118]}), .a ({w1_s3[118], w1_s2[118], w1_s1[118], w1_s0[118]}), .c ({new_AGEMA_signal_6802, new_AGEMA_signal_6801, new_AGEMA_signal_6800, addc_in[118]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_119_U1 ( .s (p256_sel), .b ({w0_s3[119], w0_s2[119], w0_s1[119], w0_s0[119]}), .a ({w1_s3[119], w1_s2[119], w1_s1[119], w1_s0[119]}), .c ({new_AGEMA_signal_6811, new_AGEMA_signal_6810, new_AGEMA_signal_6809, addc_in[119]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_120_U1 ( .s (p256_sel), .b ({w0_s3[120], w0_s2[120], w0_s1[120], w0_s0[120]}), .a ({w1_s3[120], w1_s2[120], w1_s1[120], w1_s0[120]}), .c ({new_AGEMA_signal_6820, new_AGEMA_signal_6819, new_AGEMA_signal_6818, addc_in[120]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_121_U1 ( .s (p256_sel), .b ({w0_s3[121], w0_s2[121], w0_s1[121], w0_s0[121]}), .a ({w1_s3[121], w1_s2[121], w1_s1[121], w1_s0[121]}), .c ({new_AGEMA_signal_6829, new_AGEMA_signal_6828, new_AGEMA_signal_6827, addc_in[121]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_122_U1 ( .s (p256_sel), .b ({w0_s3[122], w0_s2[122], w0_s1[122], w0_s0[122]}), .a ({w1_s3[122], w1_s2[122], w1_s1[122], w1_s0[122]}), .c ({new_AGEMA_signal_6838, new_AGEMA_signal_6837, new_AGEMA_signal_6836, addc_in[122]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_123_U1 ( .s (p256_sel), .b ({w0_s3[123], w0_s2[123], w0_s1[123], w0_s0[123]}), .a ({w1_s3[123], w1_s2[123], w1_s1[123], w1_s0[123]}), .c ({new_AGEMA_signal_6847, new_AGEMA_signal_6846, new_AGEMA_signal_6845, addc_in[123]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_124_U1 ( .s (p256_sel), .b ({w0_s3[124], w0_s2[124], w0_s1[124], w0_s0[124]}), .a ({w1_s3[124], w1_s2[124], w1_s1[124], w1_s0[124]}), .c ({new_AGEMA_signal_6856, new_AGEMA_signal_6855, new_AGEMA_signal_6854, addc_in[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_125_U1 ( .s (p256_sel), .b ({w0_s3[125], w0_s2[125], w0_s1[125], w0_s0[125]}), .a ({w1_s3[125], w1_s2[125], w1_s1[125], w1_s0[125]}), .c ({new_AGEMA_signal_6865, new_AGEMA_signal_6864, new_AGEMA_signal_6863, addc_in[125]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_126_U1 ( .s (p256_sel), .b ({w0_s3[126], w0_s2[126], w0_s1[126], w0_s0[126]}), .a ({w1_s3[126], w1_s2[126], w1_s1[126], w1_s0[126]}), .c ({new_AGEMA_signal_6874, new_AGEMA_signal_6873, new_AGEMA_signal_6872, addc_in[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst1_MUXInst_127_U1 ( .s (p256_sel), .b ({w0_s3[127], w0_s2[127], w0_s1[127], w0_s0[127]}), .a ({w1_s3[127], w1_s2[127], w1_s1[127], w1_s0[127]}), .c ({new_AGEMA_signal_6883, new_AGEMA_signal_6882, new_AGEMA_signal_6881, addc_in[127]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_U8 ( .a ({new_AGEMA_signal_6886, new_AGEMA_signal_6885, new_AGEMA_signal_6884, add_sub1_0_n8}), .b ({1'b0, 1'b0, 1'b0, add_sub1_0_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, new_AGEMA_signal_8432, add_sub1_0_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_U7 ( .a ({new_AGEMA_signal_6883, new_AGEMA_signal_6882, new_AGEMA_signal_6881, addc_in[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .c ({new_AGEMA_signal_6886, new_AGEMA_signal_6885, new_AGEMA_signal_6884, add_sub1_0_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_U6 ( .a ({new_AGEMA_signal_7498, new_AGEMA_signal_7497, new_AGEMA_signal_7496, add_sub1_0_n7}), .b ({1'b0, 1'b0, 1'b0, add_sub1_0_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_8437, new_AGEMA_signal_8436, new_AGEMA_signal_8435, add_sub1_0_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_U5 ( .a ({new_AGEMA_signal_6874, new_AGEMA_signal_6873, new_AGEMA_signal_6872, addc_in[126]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_0_addc_rom_ic_out[2]}), .c ({new_AGEMA_signal_7498, new_AGEMA_signal_7497, new_AGEMA_signal_7496, add_sub1_0_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_U4 ( .a ({new_AGEMA_signal_6889, new_AGEMA_signal_6888, new_AGEMA_signal_6887, add_sub1_0_n6}), .b ({1'b0, 1'b0, 1'b0, add_sub1_0_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, new_AGEMA_signal_8438, add_sub1_0_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_U3 ( .a ({new_AGEMA_signal_6865, new_AGEMA_signal_6864, new_AGEMA_signal_6863, addc_in[125]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_0_addc_rom_ic_out[1]}), .c ({new_AGEMA_signal_6889, new_AGEMA_signal_6888, new_AGEMA_signal_6887, add_sub1_0_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_U2 ( .a ({new_AGEMA_signal_8182, new_AGEMA_signal_8181, new_AGEMA_signal_8180, add_sub1_0_n5}), .b ({1'b0, 1'b0, 1'b0, add_sub1_0_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_8443, new_AGEMA_signal_8442, new_AGEMA_signal_8441, add_sub1_0_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_U1 ( .a ({new_AGEMA_signal_6856, new_AGEMA_signal_6855, new_AGEMA_signal_6854, addc_in[124]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_0_addc_rom_ic_out[0]}), .c ({new_AGEMA_signal_8182, new_AGEMA_signal_8181, new_AGEMA_signal_8180, add_sub1_0_n5}) ) ;
    XOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U4 ( .A (1'b0), .B (p256_sel), .Z (add_sub1_0_addc_rom_ic_out[1]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_0_addc_rom_ic1_ANF_0_n2), .B (1'b0), .ZN (add_sub1_0_addc_rom_ic_out[0]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U2 ( .A (1'b0), .B (add_sub1_0_addc_rom_ic_out[2]), .ZN (add_sub1_0_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_0_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_0_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_0_addc_rom_ic_out[2]) ) ;
    AND2_X1 add_sub1_0_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b0), .A2 (1'b0), .ZN (add_sub1_0_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n21), .B (add_sub1_0_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_0_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n19), .B (add_sub1_0_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t5), .B (add_sub1_0_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t7), .B (add_sub1_0_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n17), .B (add_sub1_0_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_0_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t6), .B (add_sub1_0_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n14), .B (add_sub1_0_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_0_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t5), .B (add_sub1_0_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_0_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_0_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_0_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_n12), .B (add_sub1_0_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_0_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t0), .B (add_sub1_0_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_0_addc_rom_rc1_ANF_1_t4), .B (add_sub1_0_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_0_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_0_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_0_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_0_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_0_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_0_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_0_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, new_AGEMA_signal_8432, add_sub1_0_addc_out[3]}), .b ({new_AGEMA_signal_8437, new_AGEMA_signal_8436, new_AGEMA_signal_8435, add_sub1_0_addc_out[2]}), .c ({new_AGEMA_signal_9142, new_AGEMA_signal_9141, new_AGEMA_signal_9140, add_sub1_0_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, new_AGEMA_signal_8438, add_sub1_0_addc_out[1]}), .b ({new_AGEMA_signal_8437, new_AGEMA_signal_8436, new_AGEMA_signal_8435, add_sub1_0_addc_out[2]}), .c ({new_AGEMA_signal_9145, new_AGEMA_signal_9144, new_AGEMA_signal_9143, add_sub1_0_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_6847, new_AGEMA_signal_6846, new_AGEMA_signal_6845, addc_in[123]}), .b ({new_AGEMA_signal_6838, new_AGEMA_signal_6837, new_AGEMA_signal_6836, addc_in[122]}), .c ({new_AGEMA_signal_6892, new_AGEMA_signal_6891, new_AGEMA_signal_6890, add_sub1_0_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_6829, new_AGEMA_signal_6828, new_AGEMA_signal_6827, addc_in[121]}), .b ({new_AGEMA_signal_6838, new_AGEMA_signal_6837, new_AGEMA_signal_6836, addc_in[122]}), .c ({new_AGEMA_signal_6895, new_AGEMA_signal_6894, new_AGEMA_signal_6893, add_sub1_0_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_6811, new_AGEMA_signal_6810, new_AGEMA_signal_6809, addc_in[119]}), .b ({new_AGEMA_signal_6802, new_AGEMA_signal_6801, new_AGEMA_signal_6800, addc_in[118]}), .c ({new_AGEMA_signal_6913, new_AGEMA_signal_6912, new_AGEMA_signal_6911, add_sub1_0_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_6793, new_AGEMA_signal_6792, new_AGEMA_signal_6791, addc_in[117]}), .b ({new_AGEMA_signal_6802, new_AGEMA_signal_6801, new_AGEMA_signal_6800, addc_in[118]}), .c ({new_AGEMA_signal_6916, new_AGEMA_signal_6915, new_AGEMA_signal_6914, add_sub1_0_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_6775, new_AGEMA_signal_6774, new_AGEMA_signal_6773, addc_in[115]}), .b ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, new_AGEMA_signal_6764, addc_in[114]}), .c ({new_AGEMA_signal_6934, new_AGEMA_signal_6933, new_AGEMA_signal_6932, add_sub1_0_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_6757, new_AGEMA_signal_6756, new_AGEMA_signal_6755, addc_in[113]}), .b ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, new_AGEMA_signal_6764, addc_in[114]}), .c ({new_AGEMA_signal_6937, new_AGEMA_signal_6936, new_AGEMA_signal_6935, add_sub1_0_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_6739, new_AGEMA_signal_6738, new_AGEMA_signal_6737, addc_in[111]}), .b ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, new_AGEMA_signal_6728, addc_in[110]}), .c ({new_AGEMA_signal_6955, new_AGEMA_signal_6954, new_AGEMA_signal_6953, add_sub1_0_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_6721, new_AGEMA_signal_6720, new_AGEMA_signal_6719, addc_in[109]}), .b ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, new_AGEMA_signal_6728, addc_in[110]}), .c ({new_AGEMA_signal_6958, new_AGEMA_signal_6957, new_AGEMA_signal_6956, add_sub1_0_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_6703, new_AGEMA_signal_6702, new_AGEMA_signal_6701, addc_in[107]}), .b ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, new_AGEMA_signal_6692, addc_in[106]}), .c ({new_AGEMA_signal_6976, new_AGEMA_signal_6975, new_AGEMA_signal_6974, add_sub1_0_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_6685, new_AGEMA_signal_6684, new_AGEMA_signal_6683, addc_in[105]}), .b ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, new_AGEMA_signal_6692, addc_in[106]}), .c ({new_AGEMA_signal_6979, new_AGEMA_signal_6978, new_AGEMA_signal_6977, add_sub1_0_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_6667, new_AGEMA_signal_6666, new_AGEMA_signal_6665, addc_in[103]}), .b ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, new_AGEMA_signal_6656, addc_in[102]}), .c ({new_AGEMA_signal_6997, new_AGEMA_signal_6996, new_AGEMA_signal_6995, add_sub1_0_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_6649, new_AGEMA_signal_6648, new_AGEMA_signal_6647, addc_in[101]}), .b ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, new_AGEMA_signal_6656, addc_in[102]}), .c ({new_AGEMA_signal_7000, new_AGEMA_signal_6999, new_AGEMA_signal_6998, add_sub1_0_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, new_AGEMA_signal_6629, addc_in[99]}), .b ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, new_AGEMA_signal_6620, addc_in[98]}), .c ({new_AGEMA_signal_7018, new_AGEMA_signal_7017, new_AGEMA_signal_7016, add_sub1_0_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, new_AGEMA_signal_6611, addc_in[97]}), .b ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, new_AGEMA_signal_6620, addc_in[98]}), .c ({new_AGEMA_signal_7021, new_AGEMA_signal_7020, new_AGEMA_signal_7019, add_sub1_0_subc_rom_sbox_0_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_U8 ( .a ({new_AGEMA_signal_7039, new_AGEMA_signal_7038, new_AGEMA_signal_7037, add_sub1_1_n8}), .b ({1'b0, 1'b0, 1'b0, add_sub1_1_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_8467, new_AGEMA_signal_8466, new_AGEMA_signal_8465, add_sub1_1_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_U7 ( .a ({new_AGEMA_signal_6595, new_AGEMA_signal_6594, new_AGEMA_signal_6593, addc_in[95]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .c ({new_AGEMA_signal_7039, new_AGEMA_signal_7038, new_AGEMA_signal_7037, add_sub1_1_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_U6 ( .a ({new_AGEMA_signal_7606, new_AGEMA_signal_7605, new_AGEMA_signal_7604, add_sub1_1_n7}), .b ({1'b0, 1'b0, 1'b0, add_sub1_1_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, new_AGEMA_signal_8468, add_sub1_1_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_U5 ( .a ({new_AGEMA_signal_6586, new_AGEMA_signal_6585, new_AGEMA_signal_6584, addc_in[94]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_1_addc_rom_ic_out[2]}), .c ({new_AGEMA_signal_7606, new_AGEMA_signal_7605, new_AGEMA_signal_7604, add_sub1_1_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_U4 ( .a ({new_AGEMA_signal_7042, new_AGEMA_signal_7041, new_AGEMA_signal_7040, add_sub1_1_n6}), .b ({1'b0, 1'b0, 1'b0, add_sub1_1_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_8473, new_AGEMA_signal_8472, new_AGEMA_signal_8471, add_sub1_1_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_U3 ( .a ({new_AGEMA_signal_6577, new_AGEMA_signal_6576, new_AGEMA_signal_6575, addc_in[93]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_1_addc_rom_ic_out[1]}), .c ({new_AGEMA_signal_7042, new_AGEMA_signal_7041, new_AGEMA_signal_7040, add_sub1_1_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_U2 ( .a ({new_AGEMA_signal_8227, new_AGEMA_signal_8226, new_AGEMA_signal_8225, add_sub1_1_n5}), .b ({1'b0, 1'b0, 1'b0, add_sub1_1_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_8476, new_AGEMA_signal_8475, new_AGEMA_signal_8474, add_sub1_1_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_U1 ( .a ({new_AGEMA_signal_6568, new_AGEMA_signal_6567, new_AGEMA_signal_6566, addc_in[92]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_1_addc_rom_ic_out[0]}), .c ({new_AGEMA_signal_8227, new_AGEMA_signal_8226, new_AGEMA_signal_8225, add_sub1_1_n5}) ) ;
    XOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U4 ( .A (1'b0), .B (p256_sel), .Z (add_sub1_1_addc_rom_ic_out[1]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_1_addc_rom_ic1_ANF_0_n2), .B (1'b1), .ZN (add_sub1_1_addc_rom_ic_out[0]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U2 ( .A (1'b0), .B (add_sub1_1_addc_rom_ic_out[2]), .ZN (add_sub1_1_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_1_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_1_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_1_addc_rom_ic_out[2]) ) ;
    AND2_X1 add_sub1_1_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b1), .A2 (1'b0), .ZN (add_sub1_1_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n21), .B (add_sub1_1_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_1_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n19), .B (add_sub1_1_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t5), .B (add_sub1_1_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t7), .B (add_sub1_1_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n17), .B (add_sub1_1_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_1_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t6), .B (add_sub1_1_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n14), .B (add_sub1_1_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_1_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t5), .B (add_sub1_1_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_1_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_1_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_1_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_n12), .B (add_sub1_1_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_1_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t0), .B (add_sub1_1_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_1_addc_rom_rc1_ANF_1_t4), .B (add_sub1_1_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_1_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_1_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_1_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_1_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_1_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_1_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_1_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_8467, new_AGEMA_signal_8466, new_AGEMA_signal_8465, add_sub1_1_addc_out[3]}), .b ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, new_AGEMA_signal_8468, add_sub1_1_addc_out[2]}), .c ({new_AGEMA_signal_9205, new_AGEMA_signal_9204, new_AGEMA_signal_9203, add_sub1_1_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_8473, new_AGEMA_signal_8472, new_AGEMA_signal_8471, add_sub1_1_addc_out[1]}), .b ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, new_AGEMA_signal_8468, add_sub1_1_addc_out[2]}), .c ({new_AGEMA_signal_9208, new_AGEMA_signal_9207, new_AGEMA_signal_9206, add_sub1_1_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_6559, new_AGEMA_signal_6558, new_AGEMA_signal_6557, addc_in[91]}), .b ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, new_AGEMA_signal_6548, addc_in[90]}), .c ({new_AGEMA_signal_7045, new_AGEMA_signal_7044, new_AGEMA_signal_7043, add_sub1_1_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_6541, new_AGEMA_signal_6540, new_AGEMA_signal_6539, addc_in[89]}), .b ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, new_AGEMA_signal_6548, addc_in[90]}), .c ({new_AGEMA_signal_7048, new_AGEMA_signal_7047, new_AGEMA_signal_7046, add_sub1_1_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, new_AGEMA_signal_6521, addc_in[87]}), .b ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, new_AGEMA_signal_6512, addc_in[86]}), .c ({new_AGEMA_signal_7066, new_AGEMA_signal_7065, new_AGEMA_signal_7064, add_sub1_1_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_6505, new_AGEMA_signal_6504, new_AGEMA_signal_6503, addc_in[85]}), .b ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, new_AGEMA_signal_6512, addc_in[86]}), .c ({new_AGEMA_signal_7069, new_AGEMA_signal_7068, new_AGEMA_signal_7067, add_sub1_1_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_6487, new_AGEMA_signal_6486, new_AGEMA_signal_6485, addc_in[83]}), .b ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, new_AGEMA_signal_6476, addc_in[82]}), .c ({new_AGEMA_signal_7087, new_AGEMA_signal_7086, new_AGEMA_signal_7085, add_sub1_1_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, new_AGEMA_signal_6467, addc_in[81]}), .b ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, new_AGEMA_signal_6476, addc_in[82]}), .c ({new_AGEMA_signal_7090, new_AGEMA_signal_7089, new_AGEMA_signal_7088, add_sub1_1_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, new_AGEMA_signal_6449, addc_in[79]}), .b ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, new_AGEMA_signal_6440, addc_in[78]}), .c ({new_AGEMA_signal_7108, new_AGEMA_signal_7107, new_AGEMA_signal_7106, add_sub1_1_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, new_AGEMA_signal_6431, addc_in[77]}), .b ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, new_AGEMA_signal_6440, addc_in[78]}), .c ({new_AGEMA_signal_7111, new_AGEMA_signal_7110, new_AGEMA_signal_7109, add_sub1_1_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, new_AGEMA_signal_6413, addc_in[75]}), .b ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, new_AGEMA_signal_6404, addc_in[74]}), .c ({new_AGEMA_signal_7129, new_AGEMA_signal_7128, new_AGEMA_signal_7127, add_sub1_1_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, new_AGEMA_signal_6395, addc_in[73]}), .b ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, new_AGEMA_signal_6404, addc_in[74]}), .c ({new_AGEMA_signal_7132, new_AGEMA_signal_7131, new_AGEMA_signal_7130, add_sub1_1_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, new_AGEMA_signal_6377, addc_in[71]}), .b ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, new_AGEMA_signal_6368, addc_in[70]}), .c ({new_AGEMA_signal_7150, new_AGEMA_signal_7149, new_AGEMA_signal_7148, add_sub1_1_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, new_AGEMA_signal_6359, addc_in[69]}), .b ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, new_AGEMA_signal_6368, addc_in[70]}), .c ({new_AGEMA_signal_7153, new_AGEMA_signal_7152, new_AGEMA_signal_7151, add_sub1_1_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, new_AGEMA_signal_6341, addc_in[67]}), .b ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, new_AGEMA_signal_6332, addc_in[66]}), .c ({new_AGEMA_signal_7171, new_AGEMA_signal_7170, new_AGEMA_signal_7169, add_sub1_1_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, new_AGEMA_signal_6323, addc_in[65]}), .b ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, new_AGEMA_signal_6332, addc_in[66]}), .c ({new_AGEMA_signal_7174, new_AGEMA_signal_7173, new_AGEMA_signal_7172, add_sub1_1_subc_rom_sbox_0_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_U8 ( .a ({new_AGEMA_signal_7192, new_AGEMA_signal_7191, new_AGEMA_signal_7190, add_sub1_2_n8}), .b ({1'b0, 1'b0, 1'b0, add_sub1_2_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_8500, new_AGEMA_signal_8499, new_AGEMA_signal_8498, add_sub1_2_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_U7 ( .a ({new_AGEMA_signal_6307, new_AGEMA_signal_6306, new_AGEMA_signal_6305, addc_in[63]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .c ({new_AGEMA_signal_7192, new_AGEMA_signal_7191, new_AGEMA_signal_7190, add_sub1_2_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_U6 ( .a ({new_AGEMA_signal_7714, new_AGEMA_signal_7713, new_AGEMA_signal_7712, add_sub1_2_n7}), .b ({1'b0, 1'b0, 1'b0, add_sub1_2_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_8503, new_AGEMA_signal_8502, new_AGEMA_signal_8501, add_sub1_2_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_U5 ( .a ({new_AGEMA_signal_6298, new_AGEMA_signal_6297, new_AGEMA_signal_6296, addc_in[62]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_2_addc_rom_ic_out[2]}), .c ({new_AGEMA_signal_7714, new_AGEMA_signal_7713, new_AGEMA_signal_7712, add_sub1_2_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_U4 ( .a ({new_AGEMA_signal_7195, new_AGEMA_signal_7194, new_AGEMA_signal_7193, add_sub1_2_n6}), .b ({1'b0, 1'b0, 1'b0, add_sub1_2_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_8506, new_AGEMA_signal_8505, new_AGEMA_signal_8504, add_sub1_2_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_U3 ( .a ({new_AGEMA_signal_6289, new_AGEMA_signal_6288, new_AGEMA_signal_6287, addc_in[61]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_2_addc_rom_ic_out[1]}), .c ({new_AGEMA_signal_7195, new_AGEMA_signal_7194, new_AGEMA_signal_7193, add_sub1_2_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_U2 ( .a ({new_AGEMA_signal_8272, new_AGEMA_signal_8271, new_AGEMA_signal_8270, add_sub1_2_n5}), .b ({1'b0, 1'b0, 1'b0, add_sub1_2_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_8509, new_AGEMA_signal_8508, new_AGEMA_signal_8507, add_sub1_2_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_U1 ( .a ({new_AGEMA_signal_6280, new_AGEMA_signal_6279, new_AGEMA_signal_6278, addc_in[60]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_2_addc_rom_ic_out[0]}), .c ({new_AGEMA_signal_8272, new_AGEMA_signal_8271, new_AGEMA_signal_8270, add_sub1_2_n5}) ) ;
    XOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U4 ( .A (1'b1), .B (p256_sel), .Z (add_sub1_2_addc_rom_ic_out[1]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_2_addc_rom_ic1_ANF_0_n2), .B (1'b0), .ZN (add_sub1_2_addc_rom_ic_out[0]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U2 ( .A (1'b1), .B (add_sub1_2_addc_rom_ic_out[2]), .ZN (add_sub1_2_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_2_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_2_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_2_addc_rom_ic_out[2]) ) ;
    AND2_X1 add_sub1_2_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b0), .A2 (1'b1), .ZN (add_sub1_2_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n21), .B (add_sub1_2_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_2_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n19), .B (add_sub1_2_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t5), .B (add_sub1_2_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t7), .B (add_sub1_2_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n17), .B (add_sub1_2_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_2_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t6), .B (add_sub1_2_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n14), .B (add_sub1_2_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_2_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t5), .B (add_sub1_2_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_2_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_2_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_2_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_n12), .B (add_sub1_2_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_2_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t0), .B (add_sub1_2_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_2_addc_rom_rc1_ANF_1_t4), .B (add_sub1_2_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_2_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_2_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_2_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_2_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_2_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_2_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_2_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_8500, new_AGEMA_signal_8499, new_AGEMA_signal_8498, add_sub1_2_addc_out[3]}), .b ({new_AGEMA_signal_8503, new_AGEMA_signal_8502, new_AGEMA_signal_8501, add_sub1_2_addc_out[2]}), .c ({new_AGEMA_signal_9268, new_AGEMA_signal_9267, new_AGEMA_signal_9266, add_sub1_2_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_8506, new_AGEMA_signal_8505, new_AGEMA_signal_8504, add_sub1_2_addc_out[1]}), .b ({new_AGEMA_signal_8503, new_AGEMA_signal_8502, new_AGEMA_signal_8501, add_sub1_2_addc_out[2]}), .c ({new_AGEMA_signal_9271, new_AGEMA_signal_9270, new_AGEMA_signal_9269, add_sub1_2_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, new_AGEMA_signal_6269, addc_in[59]}), .b ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, new_AGEMA_signal_6260, addc_in[58]}), .c ({new_AGEMA_signal_7198, new_AGEMA_signal_7197, new_AGEMA_signal_7196, add_sub1_2_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, new_AGEMA_signal_6251, addc_in[57]}), .b ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, new_AGEMA_signal_6260, addc_in[58]}), .c ({new_AGEMA_signal_7201, new_AGEMA_signal_7200, new_AGEMA_signal_7199, add_sub1_2_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, addc_in[55]}), .b ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, new_AGEMA_signal_6224, addc_in[54]}), .c ({new_AGEMA_signal_7219, new_AGEMA_signal_7218, new_AGEMA_signal_7217, add_sub1_2_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, new_AGEMA_signal_6215, addc_in[53]}), .b ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, new_AGEMA_signal_6224, addc_in[54]}), .c ({new_AGEMA_signal_7222, new_AGEMA_signal_7221, new_AGEMA_signal_7220, add_sub1_2_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, new_AGEMA_signal_6197, addc_in[51]}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, addc_in[50]}), .c ({new_AGEMA_signal_7240, new_AGEMA_signal_7239, new_AGEMA_signal_7238, add_sub1_2_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, new_AGEMA_signal_6179, addc_in[49]}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, addc_in[50]}), .c ({new_AGEMA_signal_7243, new_AGEMA_signal_7242, new_AGEMA_signal_7241, add_sub1_2_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, new_AGEMA_signal_6161, addc_in[47]}), .b ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, new_AGEMA_signal_6152, addc_in[46]}), .c ({new_AGEMA_signal_7261, new_AGEMA_signal_7260, new_AGEMA_signal_7259, add_sub1_2_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, new_AGEMA_signal_6143, addc_in[45]}), .b ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, new_AGEMA_signal_6152, addc_in[46]}), .c ({new_AGEMA_signal_7264, new_AGEMA_signal_7263, new_AGEMA_signal_7262, add_sub1_2_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, new_AGEMA_signal_6125, addc_in[43]}), .b ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, new_AGEMA_signal_6116, addc_in[42]}), .c ({new_AGEMA_signal_7282, new_AGEMA_signal_7281, new_AGEMA_signal_7280, add_sub1_2_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_6109, new_AGEMA_signal_6108, new_AGEMA_signal_6107, addc_in[41]}), .b ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, new_AGEMA_signal_6116, addc_in[42]}), .c ({new_AGEMA_signal_7285, new_AGEMA_signal_7284, new_AGEMA_signal_7283, add_sub1_2_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, new_AGEMA_signal_6089, addc_in[39]}), .b ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, new_AGEMA_signal_6080, addc_in[38]}), .c ({new_AGEMA_signal_7303, new_AGEMA_signal_7302, new_AGEMA_signal_7301, add_sub1_2_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, new_AGEMA_signal_6071, addc_in[37]}), .b ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, new_AGEMA_signal_6080, addc_in[38]}), .c ({new_AGEMA_signal_7306, new_AGEMA_signal_7305, new_AGEMA_signal_7304, add_sub1_2_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, new_AGEMA_signal_6053, addc_in[35]}), .b ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, new_AGEMA_signal_6044, addc_in[34]}), .c ({new_AGEMA_signal_7324, new_AGEMA_signal_7323, new_AGEMA_signal_7322, add_sub1_2_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, new_AGEMA_signal_6035, addc_in[33]}), .b ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, new_AGEMA_signal_6044, addc_in[34]}), .c ({new_AGEMA_signal_7327, new_AGEMA_signal_7326, new_AGEMA_signal_7325, add_sub1_2_subc_rom_sbox_0_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_U8 ( .a ({new_AGEMA_signal_7345, new_AGEMA_signal_7344, new_AGEMA_signal_7343, add_sub1_3_n8}), .b ({1'b0, 1'b0, 1'b0, add_sub1_3_addc_rom_rc_out[3]}), .c ({new_AGEMA_signal_8533, new_AGEMA_signal_8532, new_AGEMA_signal_8531, add_sub1_3_addc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_U7 ( .a ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, new_AGEMA_signal_6017, addc_in[31]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .c ({new_AGEMA_signal_7345, new_AGEMA_signal_7344, new_AGEMA_signal_7343, add_sub1_3_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_U6 ( .a ({new_AGEMA_signal_7822, new_AGEMA_signal_7821, new_AGEMA_signal_7820, add_sub1_3_n7}), .b ({1'b0, 1'b0, 1'b0, add_sub1_3_addc_rom_rc_out[2]}), .c ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, new_AGEMA_signal_8534, add_sub1_3_addc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_U5 ( .a ({new_AGEMA_signal_6010, new_AGEMA_signal_6009, new_AGEMA_signal_6008, addc_in[30]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_3_addc_rom_ic_out_2_}), .c ({new_AGEMA_signal_7822, new_AGEMA_signal_7821, new_AGEMA_signal_7820, add_sub1_3_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_U4 ( .a ({new_AGEMA_signal_7348, new_AGEMA_signal_7347, new_AGEMA_signal_7346, add_sub1_3_n6}), .b ({1'b0, 1'b0, 1'b0, add_sub1_3_addc_rom_rc_out[1]}), .c ({new_AGEMA_signal_8539, new_AGEMA_signal_8538, new_AGEMA_signal_8537, add_sub1_3_addc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_U3 ( .a ({new_AGEMA_signal_6001, new_AGEMA_signal_6000, new_AGEMA_signal_5999, addc_in[29]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_3_addc_rom_ic_out_1_}), .c ({new_AGEMA_signal_7348, new_AGEMA_signal_7347, new_AGEMA_signal_7346, add_sub1_3_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_U2 ( .a ({new_AGEMA_signal_8317, new_AGEMA_signal_8316, new_AGEMA_signal_8315, add_sub1_3_n5}), .b ({1'b0, 1'b0, 1'b0, add_sub1_3_addc_rom_rc_out[0]}), .c ({new_AGEMA_signal_8542, new_AGEMA_signal_8541, new_AGEMA_signal_8540, add_sub1_3_addc_out[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_U1 ( .a ({new_AGEMA_signal_5992, new_AGEMA_signal_5991, new_AGEMA_signal_5990, addc_in[28]}), .b ({1'b0, 1'b0, 1'b0, add_sub1_3_addc_rom_ic_out_0_}), .c ({new_AGEMA_signal_8317, new_AGEMA_signal_8316, new_AGEMA_signal_8315, add_sub1_3_n5}) ) ;
    XOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U4 ( .A (1'b1), .B (p256_sel), .Z (add_sub1_3_addc_rom_ic_out_1_) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U3 ( .A (add_sub1_3_addc_rom_ic1_ANF_0_n2), .B (1'b1), .ZN (add_sub1_3_addc_rom_ic_out_0_) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U2 ( .A (1'b1), .B (add_sub1_3_addc_rom_ic_out_2_), .ZN (add_sub1_3_addc_rom_ic1_ANF_0_n2) ) ;
    XOR2_X1 add_sub1_3_addc_rom_ic1_ANF_0_U1 ( .A (p256_sel), .B (add_sub1_3_addc_rom_ic1_ANF_0_t0), .Z (add_sub1_3_addc_rom_ic_out_2_) ) ;
    AND2_X1 add_sub1_3_addc_rom_ic1_ANF_0_t0_AND_U1 ( .A1 (1'b1), .A2 (1'b1), .ZN (add_sub1_3_addc_rom_ic1_ANF_0_t0) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U15 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n21), .B (add_sub1_3_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_3_addc_rom_rc_out[3]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U14 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n19), .B (add_sub1_3_addc_rom_rc1_ANF_1_n18), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n21) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U13 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t5), .B (add_sub1_3_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n18) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U12 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t7), .B (add_sub1_3_addc_rom_rc1_ANF_1_t2), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n19) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U11 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n17), .B (add_sub1_3_addc_rom_rc1_ANF_1_n16), .ZN (add_sub1_3_addc_rom_rc_out[2]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U10 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n15), .B (k[2]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n16) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U9 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t6), .B (add_sub1_3_addc_rom_rc1_ANF_1_t1), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n17) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U8 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n14), .B (add_sub1_3_addc_rom_rc1_ANF_1_n13), .ZN (add_sub1_3_addc_rom_rc_out[1]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U7 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t5), .B (add_sub1_3_addc_rom_rc1_ANF_1_t0), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n13) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U6 ( .A (k[0]), .B (add_sub1_3_addc_rom_rc1_ANF_1_n15), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n14) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U5 ( .A (k[1]), .B (add_sub1_3_addc_rom_rc1_ANF_1_t4), .Z (add_sub1_3_addc_rom_rc1_ANF_1_n15) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U4 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_n12), .B (add_sub1_3_addc_rom_rc1_ANF_1_n20), .ZN (add_sub1_3_addc_rom_rc_out[0]) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U3 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t0), .B (add_sub1_3_addc_rom_rc1_ANF_1_t1), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n20) ) ;
    XNOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U2 ( .A (add_sub1_3_addc_rom_rc1_ANF_1_t4), .B (add_sub1_3_addc_rom_rc1_ANF_1_t2), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_n12) ) ;
    XOR2_X1 add_sub1_3_addc_rom_rc1_ANF_1_U1 ( .A (k[2]), .B (k[3]), .Z (add_sub1_3_addc_rom_rc1_ANF_1_t3) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t0_AND_U1 ( .A1 (k[0]), .A2 (k[1]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t0) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t1_AND_U1 ( .A1 (k[1]), .A2 (k[2]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t1) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t2_AND_U1 ( .A1 (k[0]), .A2 (k[3]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t2) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t4_AND_U1 ( .A1 (add_sub1_3_addc_rom_rc1_ANF_1_t0), .A2 (add_sub1_3_addc_rom_rc1_ANF_1_t3), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t4) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t5_AND_U1 ( .A1 (k[1]), .A2 (k[3]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t5) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t6_AND_U1 ( .A1 (k[0]), .A2 (k[2]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t6) ) ;
    AND2_X1 add_sub1_3_addc_rom_rc1_ANF_1_t7_AND_U1 ( .A1 (add_sub1_3_addc_rom_rc1_ANF_1_t0), .A2 (k[3]), .ZN (add_sub1_3_addc_rom_rc1_ANF_1_t7) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U2 ( .a ({new_AGEMA_signal_8533, new_AGEMA_signal_8532, new_AGEMA_signal_8531, add_sub1_3_addc_out[3]}), .b ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, new_AGEMA_signal_8534, add_sub1_3_addc_out[2]}), .c ({new_AGEMA_signal_9331, new_AGEMA_signal_9330, new_AGEMA_signal_9329, add_sub1_3_subc_rom_sbox_7_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U1 ( .a ({new_AGEMA_signal_8539, new_AGEMA_signal_8538, new_AGEMA_signal_8537, add_sub1_3_addc_out[1]}), .b ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, new_AGEMA_signal_8534, add_sub1_3_addc_out[2]}), .c ({new_AGEMA_signal_9334, new_AGEMA_signal_9333, new_AGEMA_signal_9332, add_sub1_3_subc_rom_sbox_7_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U2 ( .a ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, new_AGEMA_signal_5981, addc_in[27]}), .b ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, new_AGEMA_signal_5972, addc_in[26]}), .c ({new_AGEMA_signal_7351, new_AGEMA_signal_7350, new_AGEMA_signal_7349, add_sub1_3_subc_rom_sbox_6_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U1 ( .a ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, new_AGEMA_signal_5963, addc_in[25]}), .b ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, new_AGEMA_signal_5972, addc_in[26]}), .c ({new_AGEMA_signal_7354, new_AGEMA_signal_7353, new_AGEMA_signal_7352, add_sub1_3_subc_rom_sbox_6_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U2 ( .a ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, new_AGEMA_signal_5945, addc_in[23]}), .b ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, new_AGEMA_signal_5936, addc_in[22]}), .c ({new_AGEMA_signal_7372, new_AGEMA_signal_7371, new_AGEMA_signal_7370, add_sub1_3_subc_rom_sbox_5_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U1 ( .a ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, new_AGEMA_signal_5927, addc_in[21]}), .b ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, new_AGEMA_signal_5936, addc_in[22]}), .c ({new_AGEMA_signal_7375, new_AGEMA_signal_7374, new_AGEMA_signal_7373, add_sub1_3_subc_rom_sbox_5_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U2 ( .a ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, new_AGEMA_signal_5909, addc_in[19]}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, new_AGEMA_signal_5900, addc_in[18]}), .c ({new_AGEMA_signal_7393, new_AGEMA_signal_7392, new_AGEMA_signal_7391, add_sub1_3_subc_rom_sbox_4_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U1 ( .a ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, new_AGEMA_signal_5891, addc_in[17]}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, new_AGEMA_signal_5900, addc_in[18]}), .c ({new_AGEMA_signal_7396, new_AGEMA_signal_7395, new_AGEMA_signal_7394, add_sub1_3_subc_rom_sbox_4_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U2 ( .a ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, new_AGEMA_signal_5873, addc_in[15]}), .b ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, new_AGEMA_signal_5864, addc_in[14]}), .c ({new_AGEMA_signal_7414, new_AGEMA_signal_7413, new_AGEMA_signal_7412, add_sub1_3_subc_rom_sbox_3_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U1 ( .a ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, new_AGEMA_signal_5855, addc_in[13]}), .b ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, new_AGEMA_signal_5864, addc_in[14]}), .c ({new_AGEMA_signal_7417, new_AGEMA_signal_7416, new_AGEMA_signal_7415, add_sub1_3_subc_rom_sbox_3_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U2 ( .a ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, new_AGEMA_signal_5837, addc_in[11]}), .b ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, new_AGEMA_signal_5828, addc_in[10]}), .c ({new_AGEMA_signal_7435, new_AGEMA_signal_7434, new_AGEMA_signal_7433, add_sub1_3_subc_rom_sbox_2_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U1 ( .a ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, new_AGEMA_signal_5819, addc_in[9]}), .b ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, new_AGEMA_signal_5828, addc_in[10]}), .c ({new_AGEMA_signal_7438, new_AGEMA_signal_7437, new_AGEMA_signal_7436, add_sub1_3_subc_rom_sbox_2_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U2 ( .a ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, new_AGEMA_signal_5801, addc_in[7]}), .b ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, new_AGEMA_signal_5792, addc_in[6]}), .c ({new_AGEMA_signal_7456, new_AGEMA_signal_7455, new_AGEMA_signal_7454, add_sub1_3_subc_rom_sbox_1_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U1 ( .a ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, new_AGEMA_signal_5783, addc_in[5]}), .b ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, new_AGEMA_signal_5792, addc_in[6]}), .c ({new_AGEMA_signal_7459, new_AGEMA_signal_7458, new_AGEMA_signal_7457, add_sub1_3_subc_rom_sbox_1_ANF_2_t5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U2 ( .a ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, new_AGEMA_signal_5765, addc_in[3]}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, new_AGEMA_signal_5756, addc_in[2]}), .c ({new_AGEMA_signal_7477, new_AGEMA_signal_7476, new_AGEMA_signal_7475, add_sub1_3_subc_rom_sbox_0_ANF_2_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U1 ( .a ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, new_AGEMA_signal_5747, addc_in[1]}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, new_AGEMA_signal_5756, addc_in[2]}), .c ({new_AGEMA_signal_7480, new_AGEMA_signal_7479, new_AGEMA_signal_7478, add_sub1_3_subc_rom_sbox_0_ANF_2_t5}) ) ;
    //ClockGatingController #(6) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_10063, new_AGEMA_signal_10062, new_AGEMA_signal_10061, add_sub1_0_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_10060, new_AGEMA_signal_10059, new_AGEMA_signal_10058, add_sub1_0_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, new_AGEMA_signal_10364, add_sub1_0_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_9151, new_AGEMA_signal_9150, new_AGEMA_signal_9149, add_sub1_0_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_9157, new_AGEMA_signal_9156, new_AGEMA_signal_9155, add_sub1_0_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_10060, new_AGEMA_signal_10059, new_AGEMA_signal_10058, add_sub1_0_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_9160, new_AGEMA_signal_9159, new_AGEMA_signal_9158, add_sub1_0_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_8437, new_AGEMA_signal_8436, new_AGEMA_signal_8435, add_sub1_0_addc_out[2]}), .c ({new_AGEMA_signal_10063, new_AGEMA_signal_10062, new_AGEMA_signal_10061, add_sub1_0_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_9142, new_AGEMA_signal_9141, new_AGEMA_signal_9140, add_sub1_0_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_10066, new_AGEMA_signal_10065, new_AGEMA_signal_10064, add_sub1_0_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, new_AGEMA_signal_10370, subc_out[124]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_9148, new_AGEMA_signal_9147, new_AGEMA_signal_9146, add_sub1_0_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_8443, new_AGEMA_signal_8442, new_AGEMA_signal_8441, add_sub1_0_addc_out[0]}), .c ({new_AGEMA_signal_10066, new_AGEMA_signal_10065, new_AGEMA_signal_10064, add_sub1_0_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, new_AGEMA_signal_8438, add_sub1_0_addc_out[1]}), .b ({new_AGEMA_signal_8437, new_AGEMA_signal_8436, new_AGEMA_signal_8435, add_sub1_0_addc_out[2]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_9148, new_AGEMA_signal_9147, new_AGEMA_signal_9146, add_sub1_0_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, new_AGEMA_signal_8438, add_sub1_0_addc_out[1]}), .b ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, new_AGEMA_signal_8432, add_sub1_0_addc_out[3]}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_9151, new_AGEMA_signal_9150, new_AGEMA_signal_9149, add_sub1_0_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_8437, new_AGEMA_signal_8436, new_AGEMA_signal_8435, add_sub1_0_addc_out[2]}), .b ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, new_AGEMA_signal_8432, add_sub1_0_addc_out[3]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_9154, new_AGEMA_signal_9153, new_AGEMA_signal_9152, add_sub1_0_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_8443, new_AGEMA_signal_8442, new_AGEMA_signal_8441, add_sub1_0_addc_out[0]}), .b ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, new_AGEMA_signal_8432, add_sub1_0_addc_out[3]}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_9157, new_AGEMA_signal_9156, new_AGEMA_signal_9155, add_sub1_0_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_8443, new_AGEMA_signal_8442, new_AGEMA_signal_8441, add_sub1_0_addc_out[0]}), .b ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, new_AGEMA_signal_8438, add_sub1_0_addc_out[1]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_9160, new_AGEMA_signal_9159, new_AGEMA_signal_9158, add_sub1_0_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_7504, new_AGEMA_signal_7503, new_AGEMA_signal_7502, add_sub1_0_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, new_AGEMA_signal_7499, add_sub1_0_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, new_AGEMA_signal_7928, add_sub1_0_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_6901, new_AGEMA_signal_6900, new_AGEMA_signal_6899, add_sub1_0_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_6907, new_AGEMA_signal_6906, new_AGEMA_signal_6905, add_sub1_0_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_7501, new_AGEMA_signal_7500, new_AGEMA_signal_7499, add_sub1_0_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_6910, new_AGEMA_signal_6909, new_AGEMA_signal_6908, add_sub1_0_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_6838, new_AGEMA_signal_6837, new_AGEMA_signal_6836, addc_in[122]}), .c ({new_AGEMA_signal_7504, new_AGEMA_signal_7503, new_AGEMA_signal_7502, add_sub1_0_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_6892, new_AGEMA_signal_6891, new_AGEMA_signal_6890, add_sub1_0_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, new_AGEMA_signal_7505, add_sub1_0_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, new_AGEMA_signal_7934, subc_out[120]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_6898, new_AGEMA_signal_6897, new_AGEMA_signal_6896, add_sub1_0_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_6820, new_AGEMA_signal_6819, new_AGEMA_signal_6818, addc_in[120]}), .c ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, new_AGEMA_signal_7505, add_sub1_0_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6829, new_AGEMA_signal_6828, new_AGEMA_signal_6827, addc_in[121]}), .b ({new_AGEMA_signal_6838, new_AGEMA_signal_6837, new_AGEMA_signal_6836, addc_in[122]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_6898, new_AGEMA_signal_6897, new_AGEMA_signal_6896, add_sub1_0_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6829, new_AGEMA_signal_6828, new_AGEMA_signal_6827, addc_in[121]}), .b ({new_AGEMA_signal_6847, new_AGEMA_signal_6846, new_AGEMA_signal_6845, addc_in[123]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_6901, new_AGEMA_signal_6900, new_AGEMA_signal_6899, add_sub1_0_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6838, new_AGEMA_signal_6837, new_AGEMA_signal_6836, addc_in[122]}), .b ({new_AGEMA_signal_6847, new_AGEMA_signal_6846, new_AGEMA_signal_6845, addc_in[123]}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_6904, new_AGEMA_signal_6903, new_AGEMA_signal_6902, add_sub1_0_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6820, new_AGEMA_signal_6819, new_AGEMA_signal_6818, addc_in[120]}), .b ({new_AGEMA_signal_6847, new_AGEMA_signal_6846, new_AGEMA_signal_6845, addc_in[123]}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_6907, new_AGEMA_signal_6906, new_AGEMA_signal_6905, add_sub1_0_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6820, new_AGEMA_signal_6819, new_AGEMA_signal_6818, addc_in[120]}), .b ({new_AGEMA_signal_6829, new_AGEMA_signal_6828, new_AGEMA_signal_6827, addc_in[121]}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_6910, new_AGEMA_signal_6909, new_AGEMA_signal_6908, add_sub1_0_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, new_AGEMA_signal_7517, add_sub1_0_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_7516, new_AGEMA_signal_7515, new_AGEMA_signal_7514, add_sub1_0_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_7939, new_AGEMA_signal_7938, new_AGEMA_signal_7937, add_sub1_0_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_6922, new_AGEMA_signal_6921, new_AGEMA_signal_6920, add_sub1_0_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_6928, new_AGEMA_signal_6927, new_AGEMA_signal_6926, add_sub1_0_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_7516, new_AGEMA_signal_7515, new_AGEMA_signal_7514, add_sub1_0_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_6931, new_AGEMA_signal_6930, new_AGEMA_signal_6929, add_sub1_0_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_6802, new_AGEMA_signal_6801, new_AGEMA_signal_6800, addc_in[118]}), .c ({new_AGEMA_signal_7519, new_AGEMA_signal_7518, new_AGEMA_signal_7517, add_sub1_0_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_6913, new_AGEMA_signal_6912, new_AGEMA_signal_6911, add_sub1_0_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_7522, new_AGEMA_signal_7521, new_AGEMA_signal_7520, add_sub1_0_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_7945, new_AGEMA_signal_7944, new_AGEMA_signal_7943, subc_out[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_6919, new_AGEMA_signal_6918, new_AGEMA_signal_6917, add_sub1_0_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_6784, new_AGEMA_signal_6783, new_AGEMA_signal_6782, addc_in[116]}), .c ({new_AGEMA_signal_7522, new_AGEMA_signal_7521, new_AGEMA_signal_7520, add_sub1_0_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6793, new_AGEMA_signal_6792, new_AGEMA_signal_6791, addc_in[117]}), .b ({new_AGEMA_signal_6802, new_AGEMA_signal_6801, new_AGEMA_signal_6800, addc_in[118]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_6919, new_AGEMA_signal_6918, new_AGEMA_signal_6917, add_sub1_0_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6793, new_AGEMA_signal_6792, new_AGEMA_signal_6791, addc_in[117]}), .b ({new_AGEMA_signal_6811, new_AGEMA_signal_6810, new_AGEMA_signal_6809, addc_in[119]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_6922, new_AGEMA_signal_6921, new_AGEMA_signal_6920, add_sub1_0_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6802, new_AGEMA_signal_6801, new_AGEMA_signal_6800, addc_in[118]}), .b ({new_AGEMA_signal_6811, new_AGEMA_signal_6810, new_AGEMA_signal_6809, addc_in[119]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_6925, new_AGEMA_signal_6924, new_AGEMA_signal_6923, add_sub1_0_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6784, new_AGEMA_signal_6783, new_AGEMA_signal_6782, addc_in[116]}), .b ({new_AGEMA_signal_6811, new_AGEMA_signal_6810, new_AGEMA_signal_6809, addc_in[119]}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_6928, new_AGEMA_signal_6927, new_AGEMA_signal_6926, add_sub1_0_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6784, new_AGEMA_signal_6783, new_AGEMA_signal_6782, addc_in[116]}), .b ({new_AGEMA_signal_6793, new_AGEMA_signal_6792, new_AGEMA_signal_6791, addc_in[117]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_6931, new_AGEMA_signal_6930, new_AGEMA_signal_6929, add_sub1_0_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_7534, new_AGEMA_signal_7533, new_AGEMA_signal_7532, add_sub1_0_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, new_AGEMA_signal_7529, add_sub1_0_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, new_AGEMA_signal_7946, add_sub1_0_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_6943, new_AGEMA_signal_6942, new_AGEMA_signal_6941, add_sub1_0_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_6949, new_AGEMA_signal_6948, new_AGEMA_signal_6947, add_sub1_0_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_7531, new_AGEMA_signal_7530, new_AGEMA_signal_7529, add_sub1_0_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_6952, new_AGEMA_signal_6951, new_AGEMA_signal_6950, add_sub1_0_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, new_AGEMA_signal_6764, addc_in[114]}), .c ({new_AGEMA_signal_7534, new_AGEMA_signal_7533, new_AGEMA_signal_7532, add_sub1_0_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_6934, new_AGEMA_signal_6933, new_AGEMA_signal_6932, add_sub1_0_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_7537, new_AGEMA_signal_7536, new_AGEMA_signal_7535, add_sub1_0_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, new_AGEMA_signal_7952, subc_out[112]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_6940, new_AGEMA_signal_6939, new_AGEMA_signal_6938, add_sub1_0_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_6748, new_AGEMA_signal_6747, new_AGEMA_signal_6746, addc_in[112]}), .c ({new_AGEMA_signal_7537, new_AGEMA_signal_7536, new_AGEMA_signal_7535, add_sub1_0_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6757, new_AGEMA_signal_6756, new_AGEMA_signal_6755, addc_in[113]}), .b ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, new_AGEMA_signal_6764, addc_in[114]}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_6940, new_AGEMA_signal_6939, new_AGEMA_signal_6938, add_sub1_0_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6757, new_AGEMA_signal_6756, new_AGEMA_signal_6755, addc_in[113]}), .b ({new_AGEMA_signal_6775, new_AGEMA_signal_6774, new_AGEMA_signal_6773, addc_in[115]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_6943, new_AGEMA_signal_6942, new_AGEMA_signal_6941, add_sub1_0_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, new_AGEMA_signal_6764, addc_in[114]}), .b ({new_AGEMA_signal_6775, new_AGEMA_signal_6774, new_AGEMA_signal_6773, addc_in[115]}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_6946, new_AGEMA_signal_6945, new_AGEMA_signal_6944, add_sub1_0_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6748, new_AGEMA_signal_6747, new_AGEMA_signal_6746, addc_in[112]}), .b ({new_AGEMA_signal_6775, new_AGEMA_signal_6774, new_AGEMA_signal_6773, addc_in[115]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_6949, new_AGEMA_signal_6948, new_AGEMA_signal_6947, add_sub1_0_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6748, new_AGEMA_signal_6747, new_AGEMA_signal_6746, addc_in[112]}), .b ({new_AGEMA_signal_6757, new_AGEMA_signal_6756, new_AGEMA_signal_6755, addc_in[113]}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_6952, new_AGEMA_signal_6951, new_AGEMA_signal_6950, add_sub1_0_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_7549, new_AGEMA_signal_7548, new_AGEMA_signal_7547, add_sub1_0_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_7546, new_AGEMA_signal_7545, new_AGEMA_signal_7544, add_sub1_0_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_7957, new_AGEMA_signal_7956, new_AGEMA_signal_7955, add_sub1_0_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_6964, new_AGEMA_signal_6963, new_AGEMA_signal_6962, add_sub1_0_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_6970, new_AGEMA_signal_6969, new_AGEMA_signal_6968, add_sub1_0_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_7546, new_AGEMA_signal_7545, new_AGEMA_signal_7544, add_sub1_0_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_6973, new_AGEMA_signal_6972, new_AGEMA_signal_6971, add_sub1_0_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, new_AGEMA_signal_6728, addc_in[110]}), .c ({new_AGEMA_signal_7549, new_AGEMA_signal_7548, new_AGEMA_signal_7547, add_sub1_0_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_6955, new_AGEMA_signal_6954, new_AGEMA_signal_6953, add_sub1_0_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_7552, new_AGEMA_signal_7551, new_AGEMA_signal_7550, add_sub1_0_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_7963, new_AGEMA_signal_7962, new_AGEMA_signal_7961, subc_out[108]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_6961, new_AGEMA_signal_6960, new_AGEMA_signal_6959, add_sub1_0_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_6712, new_AGEMA_signal_6711, new_AGEMA_signal_6710, addc_in[108]}), .c ({new_AGEMA_signal_7552, new_AGEMA_signal_7551, new_AGEMA_signal_7550, add_sub1_0_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6721, new_AGEMA_signal_6720, new_AGEMA_signal_6719, addc_in[109]}), .b ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, new_AGEMA_signal_6728, addc_in[110]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_6961, new_AGEMA_signal_6960, new_AGEMA_signal_6959, add_sub1_0_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6721, new_AGEMA_signal_6720, new_AGEMA_signal_6719, addc_in[109]}), .b ({new_AGEMA_signal_6739, new_AGEMA_signal_6738, new_AGEMA_signal_6737, addc_in[111]}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_6964, new_AGEMA_signal_6963, new_AGEMA_signal_6962, add_sub1_0_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, new_AGEMA_signal_6728, addc_in[110]}), .b ({new_AGEMA_signal_6739, new_AGEMA_signal_6738, new_AGEMA_signal_6737, addc_in[111]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_6967, new_AGEMA_signal_6966, new_AGEMA_signal_6965, add_sub1_0_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6712, new_AGEMA_signal_6711, new_AGEMA_signal_6710, addc_in[108]}), .b ({new_AGEMA_signal_6739, new_AGEMA_signal_6738, new_AGEMA_signal_6737, addc_in[111]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_6970, new_AGEMA_signal_6969, new_AGEMA_signal_6968, add_sub1_0_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6712, new_AGEMA_signal_6711, new_AGEMA_signal_6710, addc_in[108]}), .b ({new_AGEMA_signal_6721, new_AGEMA_signal_6720, new_AGEMA_signal_6719, addc_in[109]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_6973, new_AGEMA_signal_6972, new_AGEMA_signal_6971, add_sub1_0_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_7564, new_AGEMA_signal_7563, new_AGEMA_signal_7562, add_sub1_0_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_7561, new_AGEMA_signal_7560, new_AGEMA_signal_7559, add_sub1_0_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, new_AGEMA_signal_7964, add_sub1_0_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_6985, new_AGEMA_signal_6984, new_AGEMA_signal_6983, add_sub1_0_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_6991, new_AGEMA_signal_6990, new_AGEMA_signal_6989, add_sub1_0_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_7561, new_AGEMA_signal_7560, new_AGEMA_signal_7559, add_sub1_0_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_6994, new_AGEMA_signal_6993, new_AGEMA_signal_6992, add_sub1_0_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, new_AGEMA_signal_6692, addc_in[106]}), .c ({new_AGEMA_signal_7564, new_AGEMA_signal_7563, new_AGEMA_signal_7562, add_sub1_0_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_6976, new_AGEMA_signal_6975, new_AGEMA_signal_6974, add_sub1_0_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_7567, new_AGEMA_signal_7566, new_AGEMA_signal_7565, add_sub1_0_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, new_AGEMA_signal_7970, subc_out[104]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_6982, new_AGEMA_signal_6981, new_AGEMA_signal_6980, add_sub1_0_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_6676, new_AGEMA_signal_6675, new_AGEMA_signal_6674, addc_in[104]}), .c ({new_AGEMA_signal_7567, new_AGEMA_signal_7566, new_AGEMA_signal_7565, add_sub1_0_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6685, new_AGEMA_signal_6684, new_AGEMA_signal_6683, addc_in[105]}), .b ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, new_AGEMA_signal_6692, addc_in[106]}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_6982, new_AGEMA_signal_6981, new_AGEMA_signal_6980, add_sub1_0_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6685, new_AGEMA_signal_6684, new_AGEMA_signal_6683, addc_in[105]}), .b ({new_AGEMA_signal_6703, new_AGEMA_signal_6702, new_AGEMA_signal_6701, addc_in[107]}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_6985, new_AGEMA_signal_6984, new_AGEMA_signal_6983, add_sub1_0_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, new_AGEMA_signal_6692, addc_in[106]}), .b ({new_AGEMA_signal_6703, new_AGEMA_signal_6702, new_AGEMA_signal_6701, addc_in[107]}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_6988, new_AGEMA_signal_6987, new_AGEMA_signal_6986, add_sub1_0_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6676, new_AGEMA_signal_6675, new_AGEMA_signal_6674, addc_in[104]}), .b ({new_AGEMA_signal_6703, new_AGEMA_signal_6702, new_AGEMA_signal_6701, addc_in[107]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_6991, new_AGEMA_signal_6990, new_AGEMA_signal_6989, add_sub1_0_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6676, new_AGEMA_signal_6675, new_AGEMA_signal_6674, addc_in[104]}), .b ({new_AGEMA_signal_6685, new_AGEMA_signal_6684, new_AGEMA_signal_6683, addc_in[105]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_6994, new_AGEMA_signal_6993, new_AGEMA_signal_6992, add_sub1_0_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_7579, new_AGEMA_signal_7578, new_AGEMA_signal_7577, add_sub1_0_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_7576, new_AGEMA_signal_7575, new_AGEMA_signal_7574, add_sub1_0_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_7975, new_AGEMA_signal_7974, new_AGEMA_signal_7973, add_sub1_0_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_7006, new_AGEMA_signal_7005, new_AGEMA_signal_7004, add_sub1_0_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_7012, new_AGEMA_signal_7011, new_AGEMA_signal_7010, add_sub1_0_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_7576, new_AGEMA_signal_7575, new_AGEMA_signal_7574, add_sub1_0_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_7015, new_AGEMA_signal_7014, new_AGEMA_signal_7013, add_sub1_0_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, new_AGEMA_signal_6656, addc_in[102]}), .c ({new_AGEMA_signal_7579, new_AGEMA_signal_7578, new_AGEMA_signal_7577, add_sub1_0_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_6997, new_AGEMA_signal_6996, new_AGEMA_signal_6995, add_sub1_0_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_7582, new_AGEMA_signal_7581, new_AGEMA_signal_7580, add_sub1_0_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_7981, new_AGEMA_signal_7980, new_AGEMA_signal_7979, subc_out[100]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_7003, new_AGEMA_signal_7002, new_AGEMA_signal_7001, add_sub1_0_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_6640, new_AGEMA_signal_6639, new_AGEMA_signal_6638, addc_in[100]}), .c ({new_AGEMA_signal_7582, new_AGEMA_signal_7581, new_AGEMA_signal_7580, add_sub1_0_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6649, new_AGEMA_signal_6648, new_AGEMA_signal_6647, addc_in[101]}), .b ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, new_AGEMA_signal_6656, addc_in[102]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_7003, new_AGEMA_signal_7002, new_AGEMA_signal_7001, add_sub1_0_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6649, new_AGEMA_signal_6648, new_AGEMA_signal_6647, addc_in[101]}), .b ({new_AGEMA_signal_6667, new_AGEMA_signal_6666, new_AGEMA_signal_6665, addc_in[103]}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_7006, new_AGEMA_signal_7005, new_AGEMA_signal_7004, add_sub1_0_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, new_AGEMA_signal_6656, addc_in[102]}), .b ({new_AGEMA_signal_6667, new_AGEMA_signal_6666, new_AGEMA_signal_6665, addc_in[103]}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_7009, new_AGEMA_signal_7008, new_AGEMA_signal_7007, add_sub1_0_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6640, new_AGEMA_signal_6639, new_AGEMA_signal_6638, addc_in[100]}), .b ({new_AGEMA_signal_6667, new_AGEMA_signal_6666, new_AGEMA_signal_6665, addc_in[103]}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_7012, new_AGEMA_signal_7011, new_AGEMA_signal_7010, add_sub1_0_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6640, new_AGEMA_signal_6639, new_AGEMA_signal_6638, addc_in[100]}), .b ({new_AGEMA_signal_6649, new_AGEMA_signal_6648, new_AGEMA_signal_6647, addc_in[101]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_7015, new_AGEMA_signal_7014, new_AGEMA_signal_7013, add_sub1_0_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_7594, new_AGEMA_signal_7593, new_AGEMA_signal_7592, add_sub1_0_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_7591, new_AGEMA_signal_7590, new_AGEMA_signal_7589, add_sub1_0_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, new_AGEMA_signal_7982, add_sub1_0_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_7027, new_AGEMA_signal_7026, new_AGEMA_signal_7025, add_sub1_0_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_7033, new_AGEMA_signal_7032, new_AGEMA_signal_7031, add_sub1_0_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_7591, new_AGEMA_signal_7590, new_AGEMA_signal_7589, add_sub1_0_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_7036, new_AGEMA_signal_7035, new_AGEMA_signal_7034, add_sub1_0_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, new_AGEMA_signal_6620, addc_in[98]}), .c ({new_AGEMA_signal_7594, new_AGEMA_signal_7593, new_AGEMA_signal_7592, add_sub1_0_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_7018, new_AGEMA_signal_7017, new_AGEMA_signal_7016, add_sub1_0_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_7597, new_AGEMA_signal_7596, new_AGEMA_signal_7595, add_sub1_0_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, new_AGEMA_signal_7988, subc_out[96]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_7024, new_AGEMA_signal_7023, new_AGEMA_signal_7022, add_sub1_0_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, new_AGEMA_signal_6602, addc_in[96]}), .c ({new_AGEMA_signal_7597, new_AGEMA_signal_7596, new_AGEMA_signal_7595, add_sub1_0_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, new_AGEMA_signal_6611, addc_in[97]}), .b ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, new_AGEMA_signal_6620, addc_in[98]}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_7024, new_AGEMA_signal_7023, new_AGEMA_signal_7022, add_sub1_0_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, new_AGEMA_signal_6611, addc_in[97]}), .b ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, new_AGEMA_signal_6629, addc_in[99]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_7027, new_AGEMA_signal_7026, new_AGEMA_signal_7025, add_sub1_0_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6622, new_AGEMA_signal_6621, new_AGEMA_signal_6620, addc_in[98]}), .b ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, new_AGEMA_signal_6629, addc_in[99]}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_7030, new_AGEMA_signal_7029, new_AGEMA_signal_7028, add_sub1_0_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, new_AGEMA_signal_6602, addc_in[96]}), .b ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, new_AGEMA_signal_6629, addc_in[99]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_7033, new_AGEMA_signal_7032, new_AGEMA_signal_7031, add_sub1_0_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, new_AGEMA_signal_6602, addc_in[96]}), .b ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, new_AGEMA_signal_6611, addc_in[97]}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_7036, new_AGEMA_signal_7035, new_AGEMA_signal_7034, add_sub1_0_subc_rom_sbox_0_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_10099, new_AGEMA_signal_10098, new_AGEMA_signal_10097, add_sub1_1_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_10096, new_AGEMA_signal_10095, new_AGEMA_signal_10094, add_sub1_1_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_10375, new_AGEMA_signal_10374, new_AGEMA_signal_10373, add_sub1_1_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_9214, new_AGEMA_signal_9213, new_AGEMA_signal_9212, add_sub1_1_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_9220, new_AGEMA_signal_9219, new_AGEMA_signal_9218, add_sub1_1_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_10096, new_AGEMA_signal_10095, new_AGEMA_signal_10094, add_sub1_1_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_9223, new_AGEMA_signal_9222, new_AGEMA_signal_9221, add_sub1_1_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, new_AGEMA_signal_8468, add_sub1_1_addc_out[2]}), .c ({new_AGEMA_signal_10099, new_AGEMA_signal_10098, new_AGEMA_signal_10097, add_sub1_1_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_9205, new_AGEMA_signal_9204, new_AGEMA_signal_9203, add_sub1_1_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_10102, new_AGEMA_signal_10101, new_AGEMA_signal_10100, add_sub1_1_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_10381, new_AGEMA_signal_10380, new_AGEMA_signal_10379, subc_out[92]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_9211, new_AGEMA_signal_9210, new_AGEMA_signal_9209, add_sub1_1_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_8476, new_AGEMA_signal_8475, new_AGEMA_signal_8474, add_sub1_1_addc_out[0]}), .c ({new_AGEMA_signal_10102, new_AGEMA_signal_10101, new_AGEMA_signal_10100, add_sub1_1_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_8473, new_AGEMA_signal_8472, new_AGEMA_signal_8471, add_sub1_1_addc_out[1]}), .b ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, new_AGEMA_signal_8468, add_sub1_1_addc_out[2]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_9211, new_AGEMA_signal_9210, new_AGEMA_signal_9209, add_sub1_1_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_8473, new_AGEMA_signal_8472, new_AGEMA_signal_8471, add_sub1_1_addc_out[1]}), .b ({new_AGEMA_signal_8467, new_AGEMA_signal_8466, new_AGEMA_signal_8465, add_sub1_1_addc_out[3]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_9214, new_AGEMA_signal_9213, new_AGEMA_signal_9212, add_sub1_1_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_8470, new_AGEMA_signal_8469, new_AGEMA_signal_8468, add_sub1_1_addc_out[2]}), .b ({new_AGEMA_signal_8467, new_AGEMA_signal_8466, new_AGEMA_signal_8465, add_sub1_1_addc_out[3]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_9217, new_AGEMA_signal_9216, new_AGEMA_signal_9215, add_sub1_1_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_8476, new_AGEMA_signal_8475, new_AGEMA_signal_8474, add_sub1_1_addc_out[0]}), .b ({new_AGEMA_signal_8467, new_AGEMA_signal_8466, new_AGEMA_signal_8465, add_sub1_1_addc_out[3]}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_9220, new_AGEMA_signal_9219, new_AGEMA_signal_9218, add_sub1_1_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_8476, new_AGEMA_signal_8475, new_AGEMA_signal_8474, add_sub1_1_addc_out[0]}), .b ({new_AGEMA_signal_8473, new_AGEMA_signal_8472, new_AGEMA_signal_8471, add_sub1_1_addc_out[1]}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_9223, new_AGEMA_signal_9222, new_AGEMA_signal_9221, add_sub1_1_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_7612, new_AGEMA_signal_7611, new_AGEMA_signal_7610, add_sub1_1_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_7609, new_AGEMA_signal_7608, new_AGEMA_signal_7607, add_sub1_1_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_7993, new_AGEMA_signal_7992, new_AGEMA_signal_7991, add_sub1_1_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_7054, new_AGEMA_signal_7053, new_AGEMA_signal_7052, add_sub1_1_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_7060, new_AGEMA_signal_7059, new_AGEMA_signal_7058, add_sub1_1_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_7609, new_AGEMA_signal_7608, new_AGEMA_signal_7607, add_sub1_1_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_7063, new_AGEMA_signal_7062, new_AGEMA_signal_7061, add_sub1_1_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, new_AGEMA_signal_6548, addc_in[90]}), .c ({new_AGEMA_signal_7612, new_AGEMA_signal_7611, new_AGEMA_signal_7610, add_sub1_1_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_7045, new_AGEMA_signal_7044, new_AGEMA_signal_7043, add_sub1_1_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_7615, new_AGEMA_signal_7614, new_AGEMA_signal_7613, add_sub1_1_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_7999, new_AGEMA_signal_7998, new_AGEMA_signal_7997, subc_out[88]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_7051, new_AGEMA_signal_7050, new_AGEMA_signal_7049, add_sub1_1_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_6532, new_AGEMA_signal_6531, new_AGEMA_signal_6530, addc_in[88]}), .c ({new_AGEMA_signal_7615, new_AGEMA_signal_7614, new_AGEMA_signal_7613, add_sub1_1_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6541, new_AGEMA_signal_6540, new_AGEMA_signal_6539, addc_in[89]}), .b ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, new_AGEMA_signal_6548, addc_in[90]}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_7051, new_AGEMA_signal_7050, new_AGEMA_signal_7049, add_sub1_1_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6541, new_AGEMA_signal_6540, new_AGEMA_signal_6539, addc_in[89]}), .b ({new_AGEMA_signal_6559, new_AGEMA_signal_6558, new_AGEMA_signal_6557, addc_in[91]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_7054, new_AGEMA_signal_7053, new_AGEMA_signal_7052, add_sub1_1_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6550, new_AGEMA_signal_6549, new_AGEMA_signal_6548, addc_in[90]}), .b ({new_AGEMA_signal_6559, new_AGEMA_signal_6558, new_AGEMA_signal_6557, addc_in[91]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_7057, new_AGEMA_signal_7056, new_AGEMA_signal_7055, add_sub1_1_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6532, new_AGEMA_signal_6531, new_AGEMA_signal_6530, addc_in[88]}), .b ({new_AGEMA_signal_6559, new_AGEMA_signal_6558, new_AGEMA_signal_6557, addc_in[91]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_7060, new_AGEMA_signal_7059, new_AGEMA_signal_7058, add_sub1_1_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6532, new_AGEMA_signal_6531, new_AGEMA_signal_6530, addc_in[88]}), .b ({new_AGEMA_signal_6541, new_AGEMA_signal_6540, new_AGEMA_signal_6539, addc_in[89]}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_7063, new_AGEMA_signal_7062, new_AGEMA_signal_7061, add_sub1_1_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, new_AGEMA_signal_7625, add_sub1_1_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_7624, new_AGEMA_signal_7623, new_AGEMA_signal_7622, add_sub1_1_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_8002, new_AGEMA_signal_8001, new_AGEMA_signal_8000, add_sub1_1_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_7075, new_AGEMA_signal_7074, new_AGEMA_signal_7073, add_sub1_1_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_7081, new_AGEMA_signal_7080, new_AGEMA_signal_7079, add_sub1_1_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_7624, new_AGEMA_signal_7623, new_AGEMA_signal_7622, add_sub1_1_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_7084, new_AGEMA_signal_7083, new_AGEMA_signal_7082, add_sub1_1_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, new_AGEMA_signal_6512, addc_in[86]}), .c ({new_AGEMA_signal_7627, new_AGEMA_signal_7626, new_AGEMA_signal_7625, add_sub1_1_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_7066, new_AGEMA_signal_7065, new_AGEMA_signal_7064, add_sub1_1_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_7630, new_AGEMA_signal_7629, new_AGEMA_signal_7628, add_sub1_1_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_8008, new_AGEMA_signal_8007, new_AGEMA_signal_8006, subc_out[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_7072, new_AGEMA_signal_7071, new_AGEMA_signal_7070, add_sub1_1_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, new_AGEMA_signal_6494, addc_in[84]}), .c ({new_AGEMA_signal_7630, new_AGEMA_signal_7629, new_AGEMA_signal_7628, add_sub1_1_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6505, new_AGEMA_signal_6504, new_AGEMA_signal_6503, addc_in[85]}), .b ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, new_AGEMA_signal_6512, addc_in[86]}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_7072, new_AGEMA_signal_7071, new_AGEMA_signal_7070, add_sub1_1_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6505, new_AGEMA_signal_6504, new_AGEMA_signal_6503, addc_in[85]}), .b ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, new_AGEMA_signal_6521, addc_in[87]}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_7075, new_AGEMA_signal_7074, new_AGEMA_signal_7073, add_sub1_1_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6514, new_AGEMA_signal_6513, new_AGEMA_signal_6512, addc_in[86]}), .b ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, new_AGEMA_signal_6521, addc_in[87]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_7078, new_AGEMA_signal_7077, new_AGEMA_signal_7076, add_sub1_1_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, new_AGEMA_signal_6494, addc_in[84]}), .b ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, new_AGEMA_signal_6521, addc_in[87]}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_7081, new_AGEMA_signal_7080, new_AGEMA_signal_7079, add_sub1_1_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, new_AGEMA_signal_6494, addc_in[84]}), .b ({new_AGEMA_signal_6505, new_AGEMA_signal_6504, new_AGEMA_signal_6503, addc_in[85]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_7084, new_AGEMA_signal_7083, new_AGEMA_signal_7082, add_sub1_1_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_7642, new_AGEMA_signal_7641, new_AGEMA_signal_7640, add_sub1_1_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, new_AGEMA_signal_7637, add_sub1_1_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_8011, new_AGEMA_signal_8010, new_AGEMA_signal_8009, add_sub1_1_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_7096, new_AGEMA_signal_7095, new_AGEMA_signal_7094, add_sub1_1_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_7102, new_AGEMA_signal_7101, new_AGEMA_signal_7100, add_sub1_1_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_7639, new_AGEMA_signal_7638, new_AGEMA_signal_7637, add_sub1_1_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_7105, new_AGEMA_signal_7104, new_AGEMA_signal_7103, add_sub1_1_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, new_AGEMA_signal_6476, addc_in[82]}), .c ({new_AGEMA_signal_7642, new_AGEMA_signal_7641, new_AGEMA_signal_7640, add_sub1_1_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_7087, new_AGEMA_signal_7086, new_AGEMA_signal_7085, add_sub1_1_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, new_AGEMA_signal_7643, add_sub1_1_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_8017, new_AGEMA_signal_8016, new_AGEMA_signal_8015, subc_out[80]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_7093, new_AGEMA_signal_7092, new_AGEMA_signal_7091, add_sub1_1_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, new_AGEMA_signal_6458, addc_in[80]}), .c ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, new_AGEMA_signal_7643, add_sub1_1_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, new_AGEMA_signal_6467, addc_in[81]}), .b ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, new_AGEMA_signal_6476, addc_in[82]}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_7093, new_AGEMA_signal_7092, new_AGEMA_signal_7091, add_sub1_1_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, new_AGEMA_signal_6467, addc_in[81]}), .b ({new_AGEMA_signal_6487, new_AGEMA_signal_6486, new_AGEMA_signal_6485, addc_in[83]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_7096, new_AGEMA_signal_7095, new_AGEMA_signal_7094, add_sub1_1_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6478, new_AGEMA_signal_6477, new_AGEMA_signal_6476, addc_in[82]}), .b ({new_AGEMA_signal_6487, new_AGEMA_signal_6486, new_AGEMA_signal_6485, addc_in[83]}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_7099, new_AGEMA_signal_7098, new_AGEMA_signal_7097, add_sub1_1_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, new_AGEMA_signal_6458, addc_in[80]}), .b ({new_AGEMA_signal_6487, new_AGEMA_signal_6486, new_AGEMA_signal_6485, addc_in[83]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_7102, new_AGEMA_signal_7101, new_AGEMA_signal_7100, add_sub1_1_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, new_AGEMA_signal_6458, addc_in[80]}), .b ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, new_AGEMA_signal_6467, addc_in[81]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_7105, new_AGEMA_signal_7104, new_AGEMA_signal_7103, add_sub1_1_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, new_AGEMA_signal_7655, add_sub1_1_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_7654, new_AGEMA_signal_7653, new_AGEMA_signal_7652, add_sub1_1_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_8020, new_AGEMA_signal_8019, new_AGEMA_signal_8018, add_sub1_1_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_7117, new_AGEMA_signal_7116, new_AGEMA_signal_7115, add_sub1_1_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_7123, new_AGEMA_signal_7122, new_AGEMA_signal_7121, add_sub1_1_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_7654, new_AGEMA_signal_7653, new_AGEMA_signal_7652, add_sub1_1_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_7126, new_AGEMA_signal_7125, new_AGEMA_signal_7124, add_sub1_1_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, new_AGEMA_signal_6440, addc_in[78]}), .c ({new_AGEMA_signal_7657, new_AGEMA_signal_7656, new_AGEMA_signal_7655, add_sub1_1_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_7108, new_AGEMA_signal_7107, new_AGEMA_signal_7106, add_sub1_1_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_7660, new_AGEMA_signal_7659, new_AGEMA_signal_7658, add_sub1_1_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_8026, new_AGEMA_signal_8025, new_AGEMA_signal_8024, subc_out[76]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_7114, new_AGEMA_signal_7113, new_AGEMA_signal_7112, add_sub1_1_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, new_AGEMA_signal_6422, addc_in[76]}), .c ({new_AGEMA_signal_7660, new_AGEMA_signal_7659, new_AGEMA_signal_7658, add_sub1_1_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, new_AGEMA_signal_6431, addc_in[77]}), .b ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, new_AGEMA_signal_6440, addc_in[78]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_7114, new_AGEMA_signal_7113, new_AGEMA_signal_7112, add_sub1_1_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, new_AGEMA_signal_6431, addc_in[77]}), .b ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, new_AGEMA_signal_6449, addc_in[79]}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_7117, new_AGEMA_signal_7116, new_AGEMA_signal_7115, add_sub1_1_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6442, new_AGEMA_signal_6441, new_AGEMA_signal_6440, addc_in[78]}), .b ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, new_AGEMA_signal_6449, addc_in[79]}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_7120, new_AGEMA_signal_7119, new_AGEMA_signal_7118, add_sub1_1_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, new_AGEMA_signal_6422, addc_in[76]}), .b ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, new_AGEMA_signal_6449, addc_in[79]}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_7123, new_AGEMA_signal_7122, new_AGEMA_signal_7121, add_sub1_1_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, new_AGEMA_signal_6422, addc_in[76]}), .b ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, new_AGEMA_signal_6431, addc_in[77]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_7126, new_AGEMA_signal_7125, new_AGEMA_signal_7124, add_sub1_1_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_7672, new_AGEMA_signal_7671, new_AGEMA_signal_7670, add_sub1_1_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_7669, new_AGEMA_signal_7668, new_AGEMA_signal_7667, add_sub1_1_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_8029, new_AGEMA_signal_8028, new_AGEMA_signal_8027, add_sub1_1_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, new_AGEMA_signal_7136, add_sub1_1_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, new_AGEMA_signal_7142, add_sub1_1_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_7669, new_AGEMA_signal_7668, new_AGEMA_signal_7667, add_sub1_1_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_7147, new_AGEMA_signal_7146, new_AGEMA_signal_7145, add_sub1_1_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, new_AGEMA_signal_6404, addc_in[74]}), .c ({new_AGEMA_signal_7672, new_AGEMA_signal_7671, new_AGEMA_signal_7670, add_sub1_1_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_7129, new_AGEMA_signal_7128, new_AGEMA_signal_7127, add_sub1_1_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_7675, new_AGEMA_signal_7674, new_AGEMA_signal_7673, add_sub1_1_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_8035, new_AGEMA_signal_8034, new_AGEMA_signal_8033, subc_out[72]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_7135, new_AGEMA_signal_7134, new_AGEMA_signal_7133, add_sub1_1_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_6388, new_AGEMA_signal_6387, new_AGEMA_signal_6386, addc_in[72]}), .c ({new_AGEMA_signal_7675, new_AGEMA_signal_7674, new_AGEMA_signal_7673, add_sub1_1_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, new_AGEMA_signal_6395, addc_in[73]}), .b ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, new_AGEMA_signal_6404, addc_in[74]}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_7135, new_AGEMA_signal_7134, new_AGEMA_signal_7133, add_sub1_1_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, new_AGEMA_signal_6395, addc_in[73]}), .b ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, new_AGEMA_signal_6413, addc_in[75]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, new_AGEMA_signal_7136, add_sub1_1_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6406, new_AGEMA_signal_6405, new_AGEMA_signal_6404, addc_in[74]}), .b ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, new_AGEMA_signal_6413, addc_in[75]}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_7141, new_AGEMA_signal_7140, new_AGEMA_signal_7139, add_sub1_1_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6388, new_AGEMA_signal_6387, new_AGEMA_signal_6386, addc_in[72]}), .b ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, new_AGEMA_signal_6413, addc_in[75]}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, new_AGEMA_signal_7142, add_sub1_1_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6388, new_AGEMA_signal_6387, new_AGEMA_signal_6386, addc_in[72]}), .b ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, new_AGEMA_signal_6395, addc_in[73]}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_7147, new_AGEMA_signal_7146, new_AGEMA_signal_7145, add_sub1_1_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_7687, new_AGEMA_signal_7686, new_AGEMA_signal_7685, add_sub1_1_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_7684, new_AGEMA_signal_7683, new_AGEMA_signal_7682, add_sub1_1_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_8038, new_AGEMA_signal_8037, new_AGEMA_signal_8036, add_sub1_1_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_7159, new_AGEMA_signal_7158, new_AGEMA_signal_7157, add_sub1_1_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_7165, new_AGEMA_signal_7164, new_AGEMA_signal_7163, add_sub1_1_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_7684, new_AGEMA_signal_7683, new_AGEMA_signal_7682, add_sub1_1_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_7168, new_AGEMA_signal_7167, new_AGEMA_signal_7166, add_sub1_1_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, new_AGEMA_signal_6368, addc_in[70]}), .c ({new_AGEMA_signal_7687, new_AGEMA_signal_7686, new_AGEMA_signal_7685, add_sub1_1_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_7150, new_AGEMA_signal_7149, new_AGEMA_signal_7148, add_sub1_1_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_7690, new_AGEMA_signal_7689, new_AGEMA_signal_7688, add_sub1_1_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_8044, new_AGEMA_signal_8043, new_AGEMA_signal_8042, subc_out[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, new_AGEMA_signal_7154, add_sub1_1_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, new_AGEMA_signal_6350, addc_in[68]}), .c ({new_AGEMA_signal_7690, new_AGEMA_signal_7689, new_AGEMA_signal_7688, add_sub1_1_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, new_AGEMA_signal_6359, addc_in[69]}), .b ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, new_AGEMA_signal_6368, addc_in[70]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, new_AGEMA_signal_7154, add_sub1_1_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, new_AGEMA_signal_6359, addc_in[69]}), .b ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, new_AGEMA_signal_6377, addc_in[71]}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_7159, new_AGEMA_signal_7158, new_AGEMA_signal_7157, add_sub1_1_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6370, new_AGEMA_signal_6369, new_AGEMA_signal_6368, addc_in[70]}), .b ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, new_AGEMA_signal_6377, addc_in[71]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_7162, new_AGEMA_signal_7161, new_AGEMA_signal_7160, add_sub1_1_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, new_AGEMA_signal_6350, addc_in[68]}), .b ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, new_AGEMA_signal_6377, addc_in[71]}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_7165, new_AGEMA_signal_7164, new_AGEMA_signal_7163, add_sub1_1_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, new_AGEMA_signal_6350, addc_in[68]}), .b ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, new_AGEMA_signal_6359, addc_in[69]}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_7168, new_AGEMA_signal_7167, new_AGEMA_signal_7166, add_sub1_1_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_7702, new_AGEMA_signal_7701, new_AGEMA_signal_7700, add_sub1_1_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_7699, new_AGEMA_signal_7698, new_AGEMA_signal_7697, add_sub1_1_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_8047, new_AGEMA_signal_8046, new_AGEMA_signal_8045, add_sub1_1_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, new_AGEMA_signal_7178, add_sub1_1_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, new_AGEMA_signal_7184, add_sub1_1_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_7699, new_AGEMA_signal_7698, new_AGEMA_signal_7697, add_sub1_1_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_7189, new_AGEMA_signal_7188, new_AGEMA_signal_7187, add_sub1_1_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, new_AGEMA_signal_6332, addc_in[66]}), .c ({new_AGEMA_signal_7702, new_AGEMA_signal_7701, new_AGEMA_signal_7700, add_sub1_1_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_7171, new_AGEMA_signal_7170, new_AGEMA_signal_7169, add_sub1_1_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_7705, new_AGEMA_signal_7704, new_AGEMA_signal_7703, add_sub1_1_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_8053, new_AGEMA_signal_8052, new_AGEMA_signal_8051, subc_out[64]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_7177, new_AGEMA_signal_7176, new_AGEMA_signal_7175, add_sub1_1_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, new_AGEMA_signal_6314, addc_in[64]}), .c ({new_AGEMA_signal_7705, new_AGEMA_signal_7704, new_AGEMA_signal_7703, add_sub1_1_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, new_AGEMA_signal_6323, addc_in[65]}), .b ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, new_AGEMA_signal_6332, addc_in[66]}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_7177, new_AGEMA_signal_7176, new_AGEMA_signal_7175, add_sub1_1_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, new_AGEMA_signal_6323, addc_in[65]}), .b ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, new_AGEMA_signal_6341, addc_in[67]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, new_AGEMA_signal_7178, add_sub1_1_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6334, new_AGEMA_signal_6333, new_AGEMA_signal_6332, addc_in[66]}), .b ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, new_AGEMA_signal_6341, addc_in[67]}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_7183, new_AGEMA_signal_7182, new_AGEMA_signal_7181, add_sub1_1_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, new_AGEMA_signal_6314, addc_in[64]}), .b ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, new_AGEMA_signal_6341, addc_in[67]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, new_AGEMA_signal_7184, add_sub1_1_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, new_AGEMA_signal_6314, addc_in[64]}), .b ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, new_AGEMA_signal_6323, addc_in[65]}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_7189, new_AGEMA_signal_7188, new_AGEMA_signal_7187, add_sub1_1_subc_rom_sbox_0_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_10135, new_AGEMA_signal_10134, new_AGEMA_signal_10133, add_sub1_2_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_10132, new_AGEMA_signal_10131, new_AGEMA_signal_10130, add_sub1_2_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, new_AGEMA_signal_10382, add_sub1_2_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_9277, new_AGEMA_signal_9276, new_AGEMA_signal_9275, add_sub1_2_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_9283, new_AGEMA_signal_9282, new_AGEMA_signal_9281, add_sub1_2_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_10132, new_AGEMA_signal_10131, new_AGEMA_signal_10130, add_sub1_2_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_9286, new_AGEMA_signal_9285, new_AGEMA_signal_9284, add_sub1_2_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_8503, new_AGEMA_signal_8502, new_AGEMA_signal_8501, add_sub1_2_addc_out[2]}), .c ({new_AGEMA_signal_10135, new_AGEMA_signal_10134, new_AGEMA_signal_10133, add_sub1_2_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_9268, new_AGEMA_signal_9267, new_AGEMA_signal_9266, add_sub1_2_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_10138, new_AGEMA_signal_10137, new_AGEMA_signal_10136, add_sub1_2_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, new_AGEMA_signal_10388, subc_out[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_9274, new_AGEMA_signal_9273, new_AGEMA_signal_9272, add_sub1_2_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_8509, new_AGEMA_signal_8508, new_AGEMA_signal_8507, add_sub1_2_addc_out[0]}), .c ({new_AGEMA_signal_10138, new_AGEMA_signal_10137, new_AGEMA_signal_10136, add_sub1_2_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_8506, new_AGEMA_signal_8505, new_AGEMA_signal_8504, add_sub1_2_addc_out[1]}), .b ({new_AGEMA_signal_8503, new_AGEMA_signal_8502, new_AGEMA_signal_8501, add_sub1_2_addc_out[2]}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_9274, new_AGEMA_signal_9273, new_AGEMA_signal_9272, add_sub1_2_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_8506, new_AGEMA_signal_8505, new_AGEMA_signal_8504, add_sub1_2_addc_out[1]}), .b ({new_AGEMA_signal_8500, new_AGEMA_signal_8499, new_AGEMA_signal_8498, add_sub1_2_addc_out[3]}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_9277, new_AGEMA_signal_9276, new_AGEMA_signal_9275, add_sub1_2_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_8503, new_AGEMA_signal_8502, new_AGEMA_signal_8501, add_sub1_2_addc_out[2]}), .b ({new_AGEMA_signal_8500, new_AGEMA_signal_8499, new_AGEMA_signal_8498, add_sub1_2_addc_out[3]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_9280, new_AGEMA_signal_9279, new_AGEMA_signal_9278, add_sub1_2_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_8509, new_AGEMA_signal_8508, new_AGEMA_signal_8507, add_sub1_2_addc_out[0]}), .b ({new_AGEMA_signal_8500, new_AGEMA_signal_8499, new_AGEMA_signal_8498, add_sub1_2_addc_out[3]}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_9283, new_AGEMA_signal_9282, new_AGEMA_signal_9281, add_sub1_2_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_8509, new_AGEMA_signal_8508, new_AGEMA_signal_8507, add_sub1_2_addc_out[0]}), .b ({new_AGEMA_signal_8506, new_AGEMA_signal_8505, new_AGEMA_signal_8504, add_sub1_2_addc_out[1]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_9286, new_AGEMA_signal_9285, new_AGEMA_signal_9284, add_sub1_2_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_7720, new_AGEMA_signal_7719, new_AGEMA_signal_7718, add_sub1_2_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_7717, new_AGEMA_signal_7716, new_AGEMA_signal_7715, add_sub1_2_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_8056, new_AGEMA_signal_8055, new_AGEMA_signal_8054, add_sub1_2_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_7207, new_AGEMA_signal_7206, new_AGEMA_signal_7205, add_sub1_2_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_7213, new_AGEMA_signal_7212, new_AGEMA_signal_7211, add_sub1_2_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_7717, new_AGEMA_signal_7716, new_AGEMA_signal_7715, add_sub1_2_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_7216, new_AGEMA_signal_7215, new_AGEMA_signal_7214, add_sub1_2_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, new_AGEMA_signal_6260, addc_in[58]}), .c ({new_AGEMA_signal_7720, new_AGEMA_signal_7719, new_AGEMA_signal_7718, add_sub1_2_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_7198, new_AGEMA_signal_7197, new_AGEMA_signal_7196, add_sub1_2_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_7723, new_AGEMA_signal_7722, new_AGEMA_signal_7721, add_sub1_2_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_8062, new_AGEMA_signal_8061, new_AGEMA_signal_8060, subc_out[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, new_AGEMA_signal_7202, add_sub1_2_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, new_AGEMA_signal_6242, addc_in[56]}), .c ({new_AGEMA_signal_7723, new_AGEMA_signal_7722, new_AGEMA_signal_7721, add_sub1_2_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, new_AGEMA_signal_6251, addc_in[57]}), .b ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, new_AGEMA_signal_6260, addc_in[58]}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, new_AGEMA_signal_7202, add_sub1_2_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, new_AGEMA_signal_6251, addc_in[57]}), .b ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, new_AGEMA_signal_6269, addc_in[59]}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_7207, new_AGEMA_signal_7206, new_AGEMA_signal_7205, add_sub1_2_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6262, new_AGEMA_signal_6261, new_AGEMA_signal_6260, addc_in[58]}), .b ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, new_AGEMA_signal_6269, addc_in[59]}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_7210, new_AGEMA_signal_7209, new_AGEMA_signal_7208, add_sub1_2_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, new_AGEMA_signal_6242, addc_in[56]}), .b ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, new_AGEMA_signal_6269, addc_in[59]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_7213, new_AGEMA_signal_7212, new_AGEMA_signal_7211, add_sub1_2_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, new_AGEMA_signal_6242, addc_in[56]}), .b ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, new_AGEMA_signal_6251, addc_in[57]}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_7216, new_AGEMA_signal_7215, new_AGEMA_signal_7214, add_sub1_2_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_7735, new_AGEMA_signal_7734, new_AGEMA_signal_7733, add_sub1_2_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_7732, new_AGEMA_signal_7731, new_AGEMA_signal_7730, add_sub1_2_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_8065, new_AGEMA_signal_8064, new_AGEMA_signal_8063, add_sub1_2_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, new_AGEMA_signal_7226, add_sub1_2_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, new_AGEMA_signal_7232, add_sub1_2_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_7732, new_AGEMA_signal_7731, new_AGEMA_signal_7730, add_sub1_2_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_7237, new_AGEMA_signal_7236, new_AGEMA_signal_7235, add_sub1_2_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, new_AGEMA_signal_6224, addc_in[54]}), .c ({new_AGEMA_signal_7735, new_AGEMA_signal_7734, new_AGEMA_signal_7733, add_sub1_2_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_7219, new_AGEMA_signal_7218, new_AGEMA_signal_7217, add_sub1_2_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_7738, new_AGEMA_signal_7737, new_AGEMA_signal_7736, add_sub1_2_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_8071, new_AGEMA_signal_8070, new_AGEMA_signal_8069, subc_out[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_7225, new_AGEMA_signal_7224, new_AGEMA_signal_7223, add_sub1_2_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, new_AGEMA_signal_6206, addc_in[52]}), .c ({new_AGEMA_signal_7738, new_AGEMA_signal_7737, new_AGEMA_signal_7736, add_sub1_2_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, new_AGEMA_signal_6215, addc_in[53]}), .b ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, new_AGEMA_signal_6224, addc_in[54]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_7225, new_AGEMA_signal_7224, new_AGEMA_signal_7223, add_sub1_2_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, new_AGEMA_signal_6215, addc_in[53]}), .b ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, addc_in[55]}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, new_AGEMA_signal_7226, add_sub1_2_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6226, new_AGEMA_signal_6225, new_AGEMA_signal_6224, addc_in[54]}), .b ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, addc_in[55]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_7231, new_AGEMA_signal_7230, new_AGEMA_signal_7229, add_sub1_2_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, new_AGEMA_signal_6206, addc_in[52]}), .b ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, addc_in[55]}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, new_AGEMA_signal_7232, add_sub1_2_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, new_AGEMA_signal_6206, addc_in[52]}), .b ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, new_AGEMA_signal_6215, addc_in[53]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_7237, new_AGEMA_signal_7236, new_AGEMA_signal_7235, add_sub1_2_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_7750, new_AGEMA_signal_7749, new_AGEMA_signal_7748, add_sub1_2_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_7747, new_AGEMA_signal_7746, new_AGEMA_signal_7745, add_sub1_2_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_8074, new_AGEMA_signal_8073, new_AGEMA_signal_8072, add_sub1_2_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_7249, new_AGEMA_signal_7248, new_AGEMA_signal_7247, add_sub1_2_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_7255, new_AGEMA_signal_7254, new_AGEMA_signal_7253, add_sub1_2_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_7747, new_AGEMA_signal_7746, new_AGEMA_signal_7745, add_sub1_2_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_7258, new_AGEMA_signal_7257, new_AGEMA_signal_7256, add_sub1_2_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, addc_in[50]}), .c ({new_AGEMA_signal_7750, new_AGEMA_signal_7749, new_AGEMA_signal_7748, add_sub1_2_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_7240, new_AGEMA_signal_7239, new_AGEMA_signal_7238, add_sub1_2_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_7753, new_AGEMA_signal_7752, new_AGEMA_signal_7751, add_sub1_2_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_8080, new_AGEMA_signal_8079, new_AGEMA_signal_8078, subc_out[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_7246, new_AGEMA_signal_7245, new_AGEMA_signal_7244, add_sub1_2_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_6172, new_AGEMA_signal_6171, new_AGEMA_signal_6170, addc_in[48]}), .c ({new_AGEMA_signal_7753, new_AGEMA_signal_7752, new_AGEMA_signal_7751, add_sub1_2_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, new_AGEMA_signal_6179, addc_in[49]}), .b ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, addc_in[50]}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_7246, new_AGEMA_signal_7245, new_AGEMA_signal_7244, add_sub1_2_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, new_AGEMA_signal_6179, addc_in[49]}), .b ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, new_AGEMA_signal_6197, addc_in[51]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_7249, new_AGEMA_signal_7248, new_AGEMA_signal_7247, add_sub1_2_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6190, new_AGEMA_signal_6189, new_AGEMA_signal_6188, addc_in[50]}), .b ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, new_AGEMA_signal_6197, addc_in[51]}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_7252, new_AGEMA_signal_7251, new_AGEMA_signal_7250, add_sub1_2_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6172, new_AGEMA_signal_6171, new_AGEMA_signal_6170, addc_in[48]}), .b ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, new_AGEMA_signal_6197, addc_in[51]}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_7255, new_AGEMA_signal_7254, new_AGEMA_signal_7253, add_sub1_2_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6172, new_AGEMA_signal_6171, new_AGEMA_signal_6170, addc_in[48]}), .b ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, new_AGEMA_signal_6179, addc_in[49]}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_7258, new_AGEMA_signal_7257, new_AGEMA_signal_7256, add_sub1_2_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_7765, new_AGEMA_signal_7764, new_AGEMA_signal_7763, add_sub1_2_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_7762, new_AGEMA_signal_7761, new_AGEMA_signal_7760, add_sub1_2_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_8083, new_AGEMA_signal_8082, new_AGEMA_signal_8081, add_sub1_2_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_7270, new_AGEMA_signal_7269, new_AGEMA_signal_7268, add_sub1_2_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, new_AGEMA_signal_7274, add_sub1_2_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_7762, new_AGEMA_signal_7761, new_AGEMA_signal_7760, add_sub1_2_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_7279, new_AGEMA_signal_7278, new_AGEMA_signal_7277, add_sub1_2_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, new_AGEMA_signal_6152, addc_in[46]}), .c ({new_AGEMA_signal_7765, new_AGEMA_signal_7764, new_AGEMA_signal_7763, add_sub1_2_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_7261, new_AGEMA_signal_7260, new_AGEMA_signal_7259, add_sub1_2_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_7768, new_AGEMA_signal_7767, new_AGEMA_signal_7766, add_sub1_2_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_8089, new_AGEMA_signal_8088, new_AGEMA_signal_8087, subc_out[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_7267, new_AGEMA_signal_7266, new_AGEMA_signal_7265, add_sub1_2_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, new_AGEMA_signal_6134, addc_in[44]}), .c ({new_AGEMA_signal_7768, new_AGEMA_signal_7767, new_AGEMA_signal_7766, add_sub1_2_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, new_AGEMA_signal_6143, addc_in[45]}), .b ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, new_AGEMA_signal_6152, addc_in[46]}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_7267, new_AGEMA_signal_7266, new_AGEMA_signal_7265, add_sub1_2_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, new_AGEMA_signal_6143, addc_in[45]}), .b ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, new_AGEMA_signal_6161, addc_in[47]}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_7270, new_AGEMA_signal_7269, new_AGEMA_signal_7268, add_sub1_2_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6154, new_AGEMA_signal_6153, new_AGEMA_signal_6152, addc_in[46]}), .b ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, new_AGEMA_signal_6161, addc_in[47]}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_7273, new_AGEMA_signal_7272, new_AGEMA_signal_7271, add_sub1_2_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, new_AGEMA_signal_6134, addc_in[44]}), .b ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, new_AGEMA_signal_6161, addc_in[47]}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, new_AGEMA_signal_7274, add_sub1_2_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, new_AGEMA_signal_6134, addc_in[44]}), .b ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, new_AGEMA_signal_6143, addc_in[45]}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_7279, new_AGEMA_signal_7278, new_AGEMA_signal_7277, add_sub1_2_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_7780, new_AGEMA_signal_7779, new_AGEMA_signal_7778, add_sub1_2_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_7777, new_AGEMA_signal_7776, new_AGEMA_signal_7775, add_sub1_2_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_8092, new_AGEMA_signal_8091, new_AGEMA_signal_8090, add_sub1_2_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_7291, new_AGEMA_signal_7290, new_AGEMA_signal_7289, add_sub1_2_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_7297, new_AGEMA_signal_7296, new_AGEMA_signal_7295, add_sub1_2_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_7777, new_AGEMA_signal_7776, new_AGEMA_signal_7775, add_sub1_2_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_7300, new_AGEMA_signal_7299, new_AGEMA_signal_7298, add_sub1_2_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, new_AGEMA_signal_6116, addc_in[42]}), .c ({new_AGEMA_signal_7780, new_AGEMA_signal_7779, new_AGEMA_signal_7778, add_sub1_2_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_7282, new_AGEMA_signal_7281, new_AGEMA_signal_7280, add_sub1_2_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_7783, new_AGEMA_signal_7782, new_AGEMA_signal_7781, add_sub1_2_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_8098, new_AGEMA_signal_8097, new_AGEMA_signal_8096, subc_out[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, new_AGEMA_signal_7286, add_sub1_2_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, new_AGEMA_signal_6098, addc_in[40]}), .c ({new_AGEMA_signal_7783, new_AGEMA_signal_7782, new_AGEMA_signal_7781, add_sub1_2_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6109, new_AGEMA_signal_6108, new_AGEMA_signal_6107, addc_in[41]}), .b ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, new_AGEMA_signal_6116, addc_in[42]}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, new_AGEMA_signal_7286, add_sub1_2_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6109, new_AGEMA_signal_6108, new_AGEMA_signal_6107, addc_in[41]}), .b ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, new_AGEMA_signal_6125, addc_in[43]}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_7291, new_AGEMA_signal_7290, new_AGEMA_signal_7289, add_sub1_2_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6118, new_AGEMA_signal_6117, new_AGEMA_signal_6116, addc_in[42]}), .b ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, new_AGEMA_signal_6125, addc_in[43]}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_7294, new_AGEMA_signal_7293, new_AGEMA_signal_7292, add_sub1_2_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, new_AGEMA_signal_6098, addc_in[40]}), .b ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, new_AGEMA_signal_6125, addc_in[43]}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_7297, new_AGEMA_signal_7296, new_AGEMA_signal_7295, add_sub1_2_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, new_AGEMA_signal_6098, addc_in[40]}), .b ({new_AGEMA_signal_6109, new_AGEMA_signal_6108, new_AGEMA_signal_6107, addc_in[41]}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_7300, new_AGEMA_signal_7299, new_AGEMA_signal_7298, add_sub1_2_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_7795, new_AGEMA_signal_7794, new_AGEMA_signal_7793, add_sub1_2_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_7792, new_AGEMA_signal_7791, new_AGEMA_signal_7790, add_sub1_2_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_8101, new_AGEMA_signal_8100, new_AGEMA_signal_8099, add_sub1_2_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, new_AGEMA_signal_7310, add_sub1_2_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, new_AGEMA_signal_7316, add_sub1_2_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_7792, new_AGEMA_signal_7791, new_AGEMA_signal_7790, add_sub1_2_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_7321, new_AGEMA_signal_7320, new_AGEMA_signal_7319, add_sub1_2_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, new_AGEMA_signal_6080, addc_in[38]}), .c ({new_AGEMA_signal_7795, new_AGEMA_signal_7794, new_AGEMA_signal_7793, add_sub1_2_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_7303, new_AGEMA_signal_7302, new_AGEMA_signal_7301, add_sub1_2_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_7798, new_AGEMA_signal_7797, new_AGEMA_signal_7796, add_sub1_2_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_8107, new_AGEMA_signal_8106, new_AGEMA_signal_8105, subc_out[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_7309, new_AGEMA_signal_7308, new_AGEMA_signal_7307, add_sub1_2_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, new_AGEMA_signal_6062, addc_in[36]}), .c ({new_AGEMA_signal_7798, new_AGEMA_signal_7797, new_AGEMA_signal_7796, add_sub1_2_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, new_AGEMA_signal_6071, addc_in[37]}), .b ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, new_AGEMA_signal_6080, addc_in[38]}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_7309, new_AGEMA_signal_7308, new_AGEMA_signal_7307, add_sub1_2_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, new_AGEMA_signal_6071, addc_in[37]}), .b ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, new_AGEMA_signal_6089, addc_in[39]}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, new_AGEMA_signal_7310, add_sub1_2_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6082, new_AGEMA_signal_6081, new_AGEMA_signal_6080, addc_in[38]}), .b ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, new_AGEMA_signal_6089, addc_in[39]}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_7315, new_AGEMA_signal_7314, new_AGEMA_signal_7313, add_sub1_2_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, new_AGEMA_signal_6062, addc_in[36]}), .b ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, new_AGEMA_signal_6089, addc_in[39]}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, new_AGEMA_signal_7316, add_sub1_2_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, new_AGEMA_signal_6062, addc_in[36]}), .b ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, new_AGEMA_signal_6071, addc_in[37]}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_7321, new_AGEMA_signal_7320, new_AGEMA_signal_7319, add_sub1_2_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_7810, new_AGEMA_signal_7809, new_AGEMA_signal_7808, add_sub1_2_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_7807, new_AGEMA_signal_7806, new_AGEMA_signal_7805, add_sub1_2_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_8110, new_AGEMA_signal_8109, new_AGEMA_signal_8108, add_sub1_2_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_7333, new_AGEMA_signal_7332, new_AGEMA_signal_7331, add_sub1_2_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_7339, new_AGEMA_signal_7338, new_AGEMA_signal_7337, add_sub1_2_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_7807, new_AGEMA_signal_7806, new_AGEMA_signal_7805, add_sub1_2_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_7342, new_AGEMA_signal_7341, new_AGEMA_signal_7340, add_sub1_2_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, new_AGEMA_signal_6044, addc_in[34]}), .c ({new_AGEMA_signal_7810, new_AGEMA_signal_7809, new_AGEMA_signal_7808, add_sub1_2_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_7324, new_AGEMA_signal_7323, new_AGEMA_signal_7322, add_sub1_2_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_7813, new_AGEMA_signal_7812, new_AGEMA_signal_7811, add_sub1_2_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_8116, new_AGEMA_signal_8115, new_AGEMA_signal_8114, subc_out[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_7330, new_AGEMA_signal_7329, new_AGEMA_signal_7328, add_sub1_2_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, new_AGEMA_signal_6026, addc_in[32]}), .c ({new_AGEMA_signal_7813, new_AGEMA_signal_7812, new_AGEMA_signal_7811, add_sub1_2_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, new_AGEMA_signal_6035, addc_in[33]}), .b ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, new_AGEMA_signal_6044, addc_in[34]}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_7330, new_AGEMA_signal_7329, new_AGEMA_signal_7328, add_sub1_2_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, new_AGEMA_signal_6035, addc_in[33]}), .b ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, new_AGEMA_signal_6053, addc_in[35]}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_7333, new_AGEMA_signal_7332, new_AGEMA_signal_7331, add_sub1_2_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_6046, new_AGEMA_signal_6045, new_AGEMA_signal_6044, addc_in[34]}), .b ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, new_AGEMA_signal_6053, addc_in[35]}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, new_AGEMA_signal_7334, add_sub1_2_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, new_AGEMA_signal_6026, addc_in[32]}), .b ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, new_AGEMA_signal_6053, addc_in[35]}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_7339, new_AGEMA_signal_7338, new_AGEMA_signal_7337, add_sub1_2_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, new_AGEMA_signal_6026, addc_in[32]}), .b ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, new_AGEMA_signal_6035, addc_in[33]}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_7342, new_AGEMA_signal_7341, new_AGEMA_signal_7340, add_sub1_2_subc_rom_sbox_0_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U12 ( .a ({new_AGEMA_signal_10171, new_AGEMA_signal_10170, new_AGEMA_signal_10169, add_sub1_3_subc_rom_sbox_7_ANF_2_n16}), .b ({new_AGEMA_signal_10168, new_AGEMA_signal_10167, new_AGEMA_signal_10166, add_sub1_3_subc_rom_sbox_7_ANF_2_n15}), .c ({new_AGEMA_signal_10393, new_AGEMA_signal_10392, new_AGEMA_signal_10391, add_sub1_3_subc_rom_sbox_7_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U11 ( .a ({new_AGEMA_signal_9340, new_AGEMA_signal_9339, new_AGEMA_signal_9338, add_sub1_3_subc_rom_sbox_7_ANF_2_t1}), .b ({new_AGEMA_signal_9346, new_AGEMA_signal_9345, new_AGEMA_signal_9344, add_sub1_3_subc_rom_sbox_7_ANF_2_t4}), .c ({new_AGEMA_signal_10168, new_AGEMA_signal_10167, new_AGEMA_signal_10166, add_sub1_3_subc_rom_sbox_7_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U10 ( .a ({new_AGEMA_signal_9349, new_AGEMA_signal_9348, new_AGEMA_signal_9347, add_sub1_3_subc_rom_sbox_7_ANF_2_t7}), .b ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, new_AGEMA_signal_8534, add_sub1_3_addc_out[2]}), .c ({new_AGEMA_signal_10171, new_AGEMA_signal_10170, new_AGEMA_signal_10169, add_sub1_3_subc_rom_sbox_7_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U4 ( .a ({new_AGEMA_signal_9331, new_AGEMA_signal_9330, new_AGEMA_signal_9329, add_sub1_3_subc_rom_sbox_7_ANF_2_n12}), .b ({new_AGEMA_signal_10174, new_AGEMA_signal_10173, new_AGEMA_signal_10172, add_sub1_3_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_10399, new_AGEMA_signal_10398, new_AGEMA_signal_10397, subc_out[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U3 ( .a ({new_AGEMA_signal_9337, new_AGEMA_signal_9336, new_AGEMA_signal_9335, add_sub1_3_subc_rom_sbox_7_ANF_2_t0}), .b ({new_AGEMA_signal_8542, new_AGEMA_signal_8541, new_AGEMA_signal_8540, add_sub1_3_addc_out[0]}), .c ({new_AGEMA_signal_10174, new_AGEMA_signal_10173, new_AGEMA_signal_10172, add_sub1_3_subc_rom_sbox_7_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_8539, new_AGEMA_signal_8538, new_AGEMA_signal_8537, add_sub1_3_addc_out[1]}), .b ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, new_AGEMA_signal_8534, add_sub1_3_addc_out[2]}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_9337, new_AGEMA_signal_9336, new_AGEMA_signal_9335, add_sub1_3_subc_rom_sbox_7_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_8539, new_AGEMA_signal_8538, new_AGEMA_signal_8537, add_sub1_3_addc_out[1]}), .b ({new_AGEMA_signal_8533, new_AGEMA_signal_8532, new_AGEMA_signal_8531, add_sub1_3_addc_out[3]}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_9340, new_AGEMA_signal_9339, new_AGEMA_signal_9338, add_sub1_3_subc_rom_sbox_7_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_8536, new_AGEMA_signal_8535, new_AGEMA_signal_8534, add_sub1_3_addc_out[2]}), .b ({new_AGEMA_signal_8533, new_AGEMA_signal_8532, new_AGEMA_signal_8531, add_sub1_3_addc_out[3]}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_9343, new_AGEMA_signal_9342, new_AGEMA_signal_9341, add_sub1_3_subc_rom_sbox_7_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_8542, new_AGEMA_signal_8541, new_AGEMA_signal_8540, add_sub1_3_addc_out[0]}), .b ({new_AGEMA_signal_8533, new_AGEMA_signal_8532, new_AGEMA_signal_8531, add_sub1_3_addc_out[3]}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_9346, new_AGEMA_signal_9345, new_AGEMA_signal_9344, add_sub1_3_subc_rom_sbox_7_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_8542, new_AGEMA_signal_8541, new_AGEMA_signal_8540, add_sub1_3_addc_out[0]}), .b ({new_AGEMA_signal_8539, new_AGEMA_signal_8538, new_AGEMA_signal_8537, add_sub1_3_addc_out[1]}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_9349, new_AGEMA_signal_9348, new_AGEMA_signal_9347, add_sub1_3_subc_rom_sbox_7_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U12 ( .a ({new_AGEMA_signal_7828, new_AGEMA_signal_7827, new_AGEMA_signal_7826, add_sub1_3_subc_rom_sbox_6_ANF_2_n16}), .b ({new_AGEMA_signal_7825, new_AGEMA_signal_7824, new_AGEMA_signal_7823, add_sub1_3_subc_rom_sbox_6_ANF_2_n15}), .c ({new_AGEMA_signal_8119, new_AGEMA_signal_8118, new_AGEMA_signal_8117, add_sub1_3_subc_rom_sbox_6_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U11 ( .a ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, new_AGEMA_signal_7358, add_sub1_3_subc_rom_sbox_6_ANF_2_t1}), .b ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, new_AGEMA_signal_7364, add_sub1_3_subc_rom_sbox_6_ANF_2_t4}), .c ({new_AGEMA_signal_7825, new_AGEMA_signal_7824, new_AGEMA_signal_7823, add_sub1_3_subc_rom_sbox_6_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U10 ( .a ({new_AGEMA_signal_7369, new_AGEMA_signal_7368, new_AGEMA_signal_7367, add_sub1_3_subc_rom_sbox_6_ANF_2_t7}), .b ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, new_AGEMA_signal_5972, addc_in[26]}), .c ({new_AGEMA_signal_7828, new_AGEMA_signal_7827, new_AGEMA_signal_7826, add_sub1_3_subc_rom_sbox_6_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U4 ( .a ({new_AGEMA_signal_7351, new_AGEMA_signal_7350, new_AGEMA_signal_7349, add_sub1_3_subc_rom_sbox_6_ANF_2_n12}), .b ({new_AGEMA_signal_7831, new_AGEMA_signal_7830, new_AGEMA_signal_7829, add_sub1_3_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_8125, new_AGEMA_signal_8124, new_AGEMA_signal_8123, subc_out[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U3 ( .a ({new_AGEMA_signal_7357, new_AGEMA_signal_7356, new_AGEMA_signal_7355, add_sub1_3_subc_rom_sbox_6_ANF_2_t0}), .b ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, new_AGEMA_signal_5954, addc_in[24]}), .c ({new_AGEMA_signal_7831, new_AGEMA_signal_7830, new_AGEMA_signal_7829, add_sub1_3_subc_rom_sbox_6_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, new_AGEMA_signal_5963, addc_in[25]}), .b ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, new_AGEMA_signal_5972, addc_in[26]}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_7357, new_AGEMA_signal_7356, new_AGEMA_signal_7355, add_sub1_3_subc_rom_sbox_6_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, new_AGEMA_signal_5963, addc_in[25]}), .b ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, new_AGEMA_signal_5981, addc_in[27]}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, new_AGEMA_signal_7358, add_sub1_3_subc_rom_sbox_6_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5974, new_AGEMA_signal_5973, new_AGEMA_signal_5972, addc_in[26]}), .b ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, new_AGEMA_signal_5981, addc_in[27]}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_7363, new_AGEMA_signal_7362, new_AGEMA_signal_7361, add_sub1_3_subc_rom_sbox_6_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, new_AGEMA_signal_5954, addc_in[24]}), .b ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, new_AGEMA_signal_5981, addc_in[27]}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, new_AGEMA_signal_7364, add_sub1_3_subc_rom_sbox_6_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, new_AGEMA_signal_5954, addc_in[24]}), .b ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, new_AGEMA_signal_5963, addc_in[25]}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_7369, new_AGEMA_signal_7368, new_AGEMA_signal_7367, add_sub1_3_subc_rom_sbox_6_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U12 ( .a ({new_AGEMA_signal_7843, new_AGEMA_signal_7842, new_AGEMA_signal_7841, add_sub1_3_subc_rom_sbox_5_ANF_2_n16}), .b ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, new_AGEMA_signal_7838, add_sub1_3_subc_rom_sbox_5_ANF_2_n15}), .c ({new_AGEMA_signal_8128, new_AGEMA_signal_8127, new_AGEMA_signal_8126, add_sub1_3_subc_rom_sbox_5_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U11 ( .a ({new_AGEMA_signal_7381, new_AGEMA_signal_7380, new_AGEMA_signal_7379, add_sub1_3_subc_rom_sbox_5_ANF_2_t1}), .b ({new_AGEMA_signal_7387, new_AGEMA_signal_7386, new_AGEMA_signal_7385, add_sub1_3_subc_rom_sbox_5_ANF_2_t4}), .c ({new_AGEMA_signal_7840, new_AGEMA_signal_7839, new_AGEMA_signal_7838, add_sub1_3_subc_rom_sbox_5_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U10 ( .a ({new_AGEMA_signal_7390, new_AGEMA_signal_7389, new_AGEMA_signal_7388, add_sub1_3_subc_rom_sbox_5_ANF_2_t7}), .b ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, new_AGEMA_signal_5936, addc_in[22]}), .c ({new_AGEMA_signal_7843, new_AGEMA_signal_7842, new_AGEMA_signal_7841, add_sub1_3_subc_rom_sbox_5_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U4 ( .a ({new_AGEMA_signal_7372, new_AGEMA_signal_7371, new_AGEMA_signal_7370, add_sub1_3_subc_rom_sbox_5_ANF_2_n12}), .b ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, new_AGEMA_signal_7844, add_sub1_3_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_8134, new_AGEMA_signal_8133, new_AGEMA_signal_8132, subc_out[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U3 ( .a ({new_AGEMA_signal_7378, new_AGEMA_signal_7377, new_AGEMA_signal_7376, add_sub1_3_subc_rom_sbox_5_ANF_2_t0}), .b ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, new_AGEMA_signal_5918, addc_in[20]}), .c ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, new_AGEMA_signal_7844, add_sub1_3_subc_rom_sbox_5_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, new_AGEMA_signal_5927, addc_in[21]}), .b ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, new_AGEMA_signal_5936, addc_in[22]}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_7378, new_AGEMA_signal_7377, new_AGEMA_signal_7376, add_sub1_3_subc_rom_sbox_5_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, new_AGEMA_signal_5927, addc_in[21]}), .b ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, new_AGEMA_signal_5945, addc_in[23]}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_7381, new_AGEMA_signal_7380, new_AGEMA_signal_7379, add_sub1_3_subc_rom_sbox_5_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5938, new_AGEMA_signal_5937, new_AGEMA_signal_5936, addc_in[22]}), .b ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, new_AGEMA_signal_5945, addc_in[23]}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, new_AGEMA_signal_7382, add_sub1_3_subc_rom_sbox_5_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, new_AGEMA_signal_5918, addc_in[20]}), .b ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, new_AGEMA_signal_5945, addc_in[23]}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_7387, new_AGEMA_signal_7386, new_AGEMA_signal_7385, add_sub1_3_subc_rom_sbox_5_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, new_AGEMA_signal_5918, addc_in[20]}), .b ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, new_AGEMA_signal_5927, addc_in[21]}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_7390, new_AGEMA_signal_7389, new_AGEMA_signal_7388, add_sub1_3_subc_rom_sbox_5_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U12 ( .a ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, new_AGEMA_signal_7856, add_sub1_3_subc_rom_sbox_4_ANF_2_n16}), .b ({new_AGEMA_signal_7855, new_AGEMA_signal_7854, new_AGEMA_signal_7853, add_sub1_3_subc_rom_sbox_4_ANF_2_n15}), .c ({new_AGEMA_signal_8137, new_AGEMA_signal_8136, new_AGEMA_signal_8135, add_sub1_3_subc_rom_sbox_4_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U11 ( .a ({new_AGEMA_signal_7402, new_AGEMA_signal_7401, new_AGEMA_signal_7400, add_sub1_3_subc_rom_sbox_4_ANF_2_t1}), .b ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, new_AGEMA_signal_7406, add_sub1_3_subc_rom_sbox_4_ANF_2_t4}), .c ({new_AGEMA_signal_7855, new_AGEMA_signal_7854, new_AGEMA_signal_7853, add_sub1_3_subc_rom_sbox_4_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U10 ( .a ({new_AGEMA_signal_7411, new_AGEMA_signal_7410, new_AGEMA_signal_7409, add_sub1_3_subc_rom_sbox_4_ANF_2_t7}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, new_AGEMA_signal_5900, addc_in[18]}), .c ({new_AGEMA_signal_7858, new_AGEMA_signal_7857, new_AGEMA_signal_7856, add_sub1_3_subc_rom_sbox_4_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U4 ( .a ({new_AGEMA_signal_7393, new_AGEMA_signal_7392, new_AGEMA_signal_7391, add_sub1_3_subc_rom_sbox_4_ANF_2_n12}), .b ({new_AGEMA_signal_7861, new_AGEMA_signal_7860, new_AGEMA_signal_7859, add_sub1_3_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_8143, new_AGEMA_signal_8142, new_AGEMA_signal_8141, subc_out[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U3 ( .a ({new_AGEMA_signal_7399, new_AGEMA_signal_7398, new_AGEMA_signal_7397, add_sub1_3_subc_rom_sbox_4_ANF_2_t0}), .b ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, new_AGEMA_signal_5882, addc_in[16]}), .c ({new_AGEMA_signal_7861, new_AGEMA_signal_7860, new_AGEMA_signal_7859, add_sub1_3_subc_rom_sbox_4_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, new_AGEMA_signal_5891, addc_in[17]}), .b ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, new_AGEMA_signal_5900, addc_in[18]}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_7399, new_AGEMA_signal_7398, new_AGEMA_signal_7397, add_sub1_3_subc_rom_sbox_4_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, new_AGEMA_signal_5891, addc_in[17]}), .b ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, new_AGEMA_signal_5909, addc_in[19]}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_7402, new_AGEMA_signal_7401, new_AGEMA_signal_7400, add_sub1_3_subc_rom_sbox_4_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5902, new_AGEMA_signal_5901, new_AGEMA_signal_5900, addc_in[18]}), .b ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, new_AGEMA_signal_5909, addc_in[19]}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_7405, new_AGEMA_signal_7404, new_AGEMA_signal_7403, add_sub1_3_subc_rom_sbox_4_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, new_AGEMA_signal_5882, addc_in[16]}), .b ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, new_AGEMA_signal_5909, addc_in[19]}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, new_AGEMA_signal_7406, add_sub1_3_subc_rom_sbox_4_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, new_AGEMA_signal_5882, addc_in[16]}), .b ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, new_AGEMA_signal_5891, addc_in[17]}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_7411, new_AGEMA_signal_7410, new_AGEMA_signal_7409, add_sub1_3_subc_rom_sbox_4_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U12 ( .a ({new_AGEMA_signal_7873, new_AGEMA_signal_7872, new_AGEMA_signal_7871, add_sub1_3_subc_rom_sbox_3_ANF_2_n16}), .b ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, new_AGEMA_signal_7868, add_sub1_3_subc_rom_sbox_3_ANF_2_n15}), .c ({new_AGEMA_signal_8146, new_AGEMA_signal_8145, new_AGEMA_signal_8144, add_sub1_3_subc_rom_sbox_3_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U11 ( .a ({new_AGEMA_signal_7423, new_AGEMA_signal_7422, new_AGEMA_signal_7421, add_sub1_3_subc_rom_sbox_3_ANF_2_t1}), .b ({new_AGEMA_signal_7429, new_AGEMA_signal_7428, new_AGEMA_signal_7427, add_sub1_3_subc_rom_sbox_3_ANF_2_t4}), .c ({new_AGEMA_signal_7870, new_AGEMA_signal_7869, new_AGEMA_signal_7868, add_sub1_3_subc_rom_sbox_3_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U10 ( .a ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, new_AGEMA_signal_7430, add_sub1_3_subc_rom_sbox_3_ANF_2_t7}), .b ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, new_AGEMA_signal_5864, addc_in[14]}), .c ({new_AGEMA_signal_7873, new_AGEMA_signal_7872, new_AGEMA_signal_7871, add_sub1_3_subc_rom_sbox_3_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U4 ( .a ({new_AGEMA_signal_7414, new_AGEMA_signal_7413, new_AGEMA_signal_7412, add_sub1_3_subc_rom_sbox_3_ANF_2_n12}), .b ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, new_AGEMA_signal_7874, add_sub1_3_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_8152, new_AGEMA_signal_8151, new_AGEMA_signal_8150, subc_out[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U3 ( .a ({new_AGEMA_signal_7420, new_AGEMA_signal_7419, new_AGEMA_signal_7418, add_sub1_3_subc_rom_sbox_3_ANF_2_t0}), .b ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, new_AGEMA_signal_5846, addc_in[12]}), .c ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, new_AGEMA_signal_7874, add_sub1_3_subc_rom_sbox_3_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, new_AGEMA_signal_5855, addc_in[13]}), .b ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, new_AGEMA_signal_5864, addc_in[14]}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_7420, new_AGEMA_signal_7419, new_AGEMA_signal_7418, add_sub1_3_subc_rom_sbox_3_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, new_AGEMA_signal_5855, addc_in[13]}), .b ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, new_AGEMA_signal_5873, addc_in[15]}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_7423, new_AGEMA_signal_7422, new_AGEMA_signal_7421, add_sub1_3_subc_rom_sbox_3_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5866, new_AGEMA_signal_5865, new_AGEMA_signal_5864, addc_in[14]}), .b ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, new_AGEMA_signal_5873, addc_in[15]}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_7426, new_AGEMA_signal_7425, new_AGEMA_signal_7424, add_sub1_3_subc_rom_sbox_3_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, new_AGEMA_signal_5846, addc_in[12]}), .b ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, new_AGEMA_signal_5873, addc_in[15]}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_7429, new_AGEMA_signal_7428, new_AGEMA_signal_7427, add_sub1_3_subc_rom_sbox_3_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, new_AGEMA_signal_5846, addc_in[12]}), .b ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, new_AGEMA_signal_5855, addc_in[13]}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_7432, new_AGEMA_signal_7431, new_AGEMA_signal_7430, add_sub1_3_subc_rom_sbox_3_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U12 ( .a ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, new_AGEMA_signal_7886, add_sub1_3_subc_rom_sbox_2_ANF_2_n16}), .b ({new_AGEMA_signal_7885, new_AGEMA_signal_7884, new_AGEMA_signal_7883, add_sub1_3_subc_rom_sbox_2_ANF_2_n15}), .c ({new_AGEMA_signal_8155, new_AGEMA_signal_8154, new_AGEMA_signal_8153, add_sub1_3_subc_rom_sbox_2_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U11 ( .a ({new_AGEMA_signal_7444, new_AGEMA_signal_7443, new_AGEMA_signal_7442, add_sub1_3_subc_rom_sbox_2_ANF_2_t1}), .b ({new_AGEMA_signal_7450, new_AGEMA_signal_7449, new_AGEMA_signal_7448, add_sub1_3_subc_rom_sbox_2_ANF_2_t4}), .c ({new_AGEMA_signal_7885, new_AGEMA_signal_7884, new_AGEMA_signal_7883, add_sub1_3_subc_rom_sbox_2_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U10 ( .a ({new_AGEMA_signal_7453, new_AGEMA_signal_7452, new_AGEMA_signal_7451, add_sub1_3_subc_rom_sbox_2_ANF_2_t7}), .b ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, new_AGEMA_signal_5828, addc_in[10]}), .c ({new_AGEMA_signal_7888, new_AGEMA_signal_7887, new_AGEMA_signal_7886, add_sub1_3_subc_rom_sbox_2_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U4 ( .a ({new_AGEMA_signal_7435, new_AGEMA_signal_7434, new_AGEMA_signal_7433, add_sub1_3_subc_rom_sbox_2_ANF_2_n12}), .b ({new_AGEMA_signal_7891, new_AGEMA_signal_7890, new_AGEMA_signal_7889, add_sub1_3_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_8161, new_AGEMA_signal_8160, new_AGEMA_signal_8159, subc_out[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U3 ( .a ({new_AGEMA_signal_7441, new_AGEMA_signal_7440, new_AGEMA_signal_7439, add_sub1_3_subc_rom_sbox_2_ANF_2_t0}), .b ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, new_AGEMA_signal_5810, addc_in[8]}), .c ({new_AGEMA_signal_7891, new_AGEMA_signal_7890, new_AGEMA_signal_7889, add_sub1_3_subc_rom_sbox_2_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, new_AGEMA_signal_5819, addc_in[9]}), .b ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, new_AGEMA_signal_5828, addc_in[10]}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_7441, new_AGEMA_signal_7440, new_AGEMA_signal_7439, add_sub1_3_subc_rom_sbox_2_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, new_AGEMA_signal_5819, addc_in[9]}), .b ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, new_AGEMA_signal_5837, addc_in[11]}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_7444, new_AGEMA_signal_7443, new_AGEMA_signal_7442, add_sub1_3_subc_rom_sbox_2_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5830, new_AGEMA_signal_5829, new_AGEMA_signal_5828, addc_in[10]}), .b ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, new_AGEMA_signal_5837, addc_in[11]}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_7447, new_AGEMA_signal_7446, new_AGEMA_signal_7445, add_sub1_3_subc_rom_sbox_2_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, new_AGEMA_signal_5810, addc_in[8]}), .b ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, new_AGEMA_signal_5837, addc_in[11]}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_7450, new_AGEMA_signal_7449, new_AGEMA_signal_7448, add_sub1_3_subc_rom_sbox_2_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, new_AGEMA_signal_5810, addc_in[8]}), .b ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, new_AGEMA_signal_5819, addc_in[9]}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_7453, new_AGEMA_signal_7452, new_AGEMA_signal_7451, add_sub1_3_subc_rom_sbox_2_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U12 ( .a ({new_AGEMA_signal_7903, new_AGEMA_signal_7902, new_AGEMA_signal_7901, add_sub1_3_subc_rom_sbox_1_ANF_2_n16}), .b ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, new_AGEMA_signal_7898, add_sub1_3_subc_rom_sbox_1_ANF_2_n15}), .c ({new_AGEMA_signal_8164, new_AGEMA_signal_8163, new_AGEMA_signal_8162, add_sub1_3_subc_rom_sbox_1_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U11 ( .a ({new_AGEMA_signal_7465, new_AGEMA_signal_7464, new_AGEMA_signal_7463, add_sub1_3_subc_rom_sbox_1_ANF_2_t1}), .b ({new_AGEMA_signal_7471, new_AGEMA_signal_7470, new_AGEMA_signal_7469, add_sub1_3_subc_rom_sbox_1_ANF_2_t4}), .c ({new_AGEMA_signal_7900, new_AGEMA_signal_7899, new_AGEMA_signal_7898, add_sub1_3_subc_rom_sbox_1_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U10 ( .a ({new_AGEMA_signal_7474, new_AGEMA_signal_7473, new_AGEMA_signal_7472, add_sub1_3_subc_rom_sbox_1_ANF_2_t7}), .b ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, new_AGEMA_signal_5792, addc_in[6]}), .c ({new_AGEMA_signal_7903, new_AGEMA_signal_7902, new_AGEMA_signal_7901, add_sub1_3_subc_rom_sbox_1_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U4 ( .a ({new_AGEMA_signal_7456, new_AGEMA_signal_7455, new_AGEMA_signal_7454, add_sub1_3_subc_rom_sbox_1_ANF_2_n12}), .b ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, new_AGEMA_signal_7904, add_sub1_3_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_8170, new_AGEMA_signal_8169, new_AGEMA_signal_8168, subc_out[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U3 ( .a ({new_AGEMA_signal_7462, new_AGEMA_signal_7461, new_AGEMA_signal_7460, add_sub1_3_subc_rom_sbox_1_ANF_2_t0}), .b ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, new_AGEMA_signal_5774, addc_in[4]}), .c ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, new_AGEMA_signal_7904, add_sub1_3_subc_rom_sbox_1_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, new_AGEMA_signal_5783, addc_in[5]}), .b ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, new_AGEMA_signal_5792, addc_in[6]}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_7462, new_AGEMA_signal_7461, new_AGEMA_signal_7460, add_sub1_3_subc_rom_sbox_1_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, new_AGEMA_signal_5783, addc_in[5]}), .b ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, new_AGEMA_signal_5801, addc_in[7]}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_7465, new_AGEMA_signal_7464, new_AGEMA_signal_7463, add_sub1_3_subc_rom_sbox_1_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5794, new_AGEMA_signal_5793, new_AGEMA_signal_5792, addc_in[6]}), .b ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, new_AGEMA_signal_5801, addc_in[7]}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_7468, new_AGEMA_signal_7467, new_AGEMA_signal_7466, add_sub1_3_subc_rom_sbox_1_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, new_AGEMA_signal_5774, addc_in[4]}), .b ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, new_AGEMA_signal_5801, addc_in[7]}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_7471, new_AGEMA_signal_7470, new_AGEMA_signal_7469, add_sub1_3_subc_rom_sbox_1_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, new_AGEMA_signal_5774, addc_in[4]}), .b ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, new_AGEMA_signal_5783, addc_in[5]}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_7474, new_AGEMA_signal_7473, new_AGEMA_signal_7472, add_sub1_3_subc_rom_sbox_1_ANF_2_t7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U12 ( .a ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, new_AGEMA_signal_7916, add_sub1_3_subc_rom_sbox_0_ANF_2_n16}), .b ({new_AGEMA_signal_7915, new_AGEMA_signal_7914, new_AGEMA_signal_7913, add_sub1_3_subc_rom_sbox_0_ANF_2_n15}), .c ({new_AGEMA_signal_8173, new_AGEMA_signal_8172, new_AGEMA_signal_8171, add_sub1_3_subc_rom_sbox_0_ANF_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U11 ( .a ({new_AGEMA_signal_7486, new_AGEMA_signal_7485, new_AGEMA_signal_7484, add_sub1_3_subc_rom_sbox_0_ANF_2_t1}), .b ({new_AGEMA_signal_7492, new_AGEMA_signal_7491, new_AGEMA_signal_7490, add_sub1_3_subc_rom_sbox_0_ANF_2_t4}), .c ({new_AGEMA_signal_7915, new_AGEMA_signal_7914, new_AGEMA_signal_7913, add_sub1_3_subc_rom_sbox_0_ANF_2_n15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U10 ( .a ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, new_AGEMA_signal_7493, add_sub1_3_subc_rom_sbox_0_ANF_2_t7}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, new_AGEMA_signal_5756, addc_in[2]}), .c ({new_AGEMA_signal_7918, new_AGEMA_signal_7917, new_AGEMA_signal_7916, add_sub1_3_subc_rom_sbox_0_ANF_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U4 ( .a ({new_AGEMA_signal_7477, new_AGEMA_signal_7476, new_AGEMA_signal_7475, add_sub1_3_subc_rom_sbox_0_ANF_2_n12}), .b ({new_AGEMA_signal_7921, new_AGEMA_signal_7920, new_AGEMA_signal_7919, add_sub1_3_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_8179, new_AGEMA_signal_8178, new_AGEMA_signal_8177, subc_out[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U3 ( .a ({new_AGEMA_signal_7483, new_AGEMA_signal_7482, new_AGEMA_signal_7481, add_sub1_3_subc_rom_sbox_0_ANF_2_t0}), .b ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, new_AGEMA_signal_5738, addc_in[0]}), .c ({new_AGEMA_signal_7921, new_AGEMA_signal_7920, new_AGEMA_signal_7919, add_sub1_3_subc_rom_sbox_0_ANF_2_n19}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t0_AND_U1 ( .a ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, new_AGEMA_signal_5747, addc_in[1]}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, new_AGEMA_signal_5756, addc_in[2]}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_7483, new_AGEMA_signal_7482, new_AGEMA_signal_7481, add_sub1_3_subc_rom_sbox_0_ANF_2_t0}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t1_AND_U1 ( .a ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, new_AGEMA_signal_5747, addc_in[1]}), .b ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, new_AGEMA_signal_5765, addc_in[3]}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_7486, new_AGEMA_signal_7485, new_AGEMA_signal_7484, add_sub1_3_subc_rom_sbox_0_ANF_2_t1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t2_AND_U1 ( .a ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, new_AGEMA_signal_5756, addc_in[2]}), .b ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, new_AGEMA_signal_5765, addc_in[3]}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, new_AGEMA_signal_7487, add_sub1_3_subc_rom_sbox_0_ANF_2_t2}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t4_AND_U1 ( .a ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, new_AGEMA_signal_5738, addc_in[0]}), .b ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, new_AGEMA_signal_5765, addc_in[3]}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_7492, new_AGEMA_signal_7491, new_AGEMA_signal_7490, add_sub1_3_subc_rom_sbox_0_ANF_2_t4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t7_AND_U1 ( .a ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, new_AGEMA_signal_5738, addc_in[0]}), .b ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, new_AGEMA_signal_5747, addc_in[1]}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_7495, new_AGEMA_signal_7494, new_AGEMA_signal_7493, add_sub1_3_subc_rom_sbox_0_ANF_2_t7}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, new_AGEMA_signal_7988, subc_out[96]}), .a ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, new_AGEMA_signal_7952, subc_out[112]}), .c ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7981, new_AGEMA_signal_7980, new_AGEMA_signal_7979, subc_out[100]}), .a ({new_AGEMA_signal_7945, new_AGEMA_signal_7944, new_AGEMA_signal_7943, subc_out[116]}), .c ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, new_AGEMA_signal_7970, subc_out[104]}), .a ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, new_AGEMA_signal_7934, subc_out[120]}), .c ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7963, new_AGEMA_signal_7962, new_AGEMA_signal_7961, subc_out[108]}), .a ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, new_AGEMA_signal_10370, subc_out[124]}), .c ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7954, new_AGEMA_signal_7953, new_AGEMA_signal_7952, subc_out[112]}), .a ({new_AGEMA_signal_7990, new_AGEMA_signal_7989, new_AGEMA_signal_7988, subc_out[96]}), .c ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7945, new_AGEMA_signal_7944, new_AGEMA_signal_7943, subc_out[116]}), .a ({new_AGEMA_signal_7981, new_AGEMA_signal_7980, new_AGEMA_signal_7979, subc_out[100]}), .c ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7936, new_AGEMA_signal_7935, new_AGEMA_signal_7934, subc_out[120]}), .a ({new_AGEMA_signal_7972, new_AGEMA_signal_7971, new_AGEMA_signal_7970, subc_out[104]}), .c ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10372, new_AGEMA_signal_10371, new_AGEMA_signal_10370, subc_out[124]}), .a ({new_AGEMA_signal_7963, new_AGEMA_signal_7962, new_AGEMA_signal_7961, subc_out[108]}), .c ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10381, new_AGEMA_signal_10380, new_AGEMA_signal_10379, subc_out[92]}), .a ({new_AGEMA_signal_8026, new_AGEMA_signal_8025, new_AGEMA_signal_8024, subc_out[76]}), .c ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8053, new_AGEMA_signal_8052, new_AGEMA_signal_8051, subc_out[64]}), .a ({new_AGEMA_signal_8017, new_AGEMA_signal_8016, new_AGEMA_signal_8015, subc_out[80]}), .c ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8044, new_AGEMA_signal_8043, new_AGEMA_signal_8042, subc_out[68]}), .a ({new_AGEMA_signal_8008, new_AGEMA_signal_8007, new_AGEMA_signal_8006, subc_out[84]}), .c ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8035, new_AGEMA_signal_8034, new_AGEMA_signal_8033, subc_out[72]}), .a ({new_AGEMA_signal_7999, new_AGEMA_signal_7998, new_AGEMA_signal_7997, subc_out[88]}), .c ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8026, new_AGEMA_signal_8025, new_AGEMA_signal_8024, subc_out[76]}), .a ({new_AGEMA_signal_10381, new_AGEMA_signal_10380, new_AGEMA_signal_10379, subc_out[92]}), .c ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8017, new_AGEMA_signal_8016, new_AGEMA_signal_8015, subc_out[80]}), .a ({new_AGEMA_signal_8053, new_AGEMA_signal_8052, new_AGEMA_signal_8051, subc_out[64]}), .c ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8008, new_AGEMA_signal_8007, new_AGEMA_signal_8006, subc_out[84]}), .a ({new_AGEMA_signal_8044, new_AGEMA_signal_8043, new_AGEMA_signal_8042, subc_out[68]}), .c ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_7999, new_AGEMA_signal_7998, new_AGEMA_signal_7997, subc_out[88]}), .a ({new_AGEMA_signal_8035, new_AGEMA_signal_8034, new_AGEMA_signal_8033, subc_out[72]}), .c ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8062, new_AGEMA_signal_8061, new_AGEMA_signal_8060, subc_out[56]}), .a ({new_AGEMA_signal_8098, new_AGEMA_signal_8097, new_AGEMA_signal_8096, subc_out[40]}), .c ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, new_AGEMA_signal_10388, subc_out[60]}), .a ({new_AGEMA_signal_8089, new_AGEMA_signal_8088, new_AGEMA_signal_8087, subc_out[44]}), .c ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8116, new_AGEMA_signal_8115, new_AGEMA_signal_8114, subc_out[32]}), .a ({new_AGEMA_signal_8080, new_AGEMA_signal_8079, new_AGEMA_signal_8078, subc_out[48]}), .c ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8107, new_AGEMA_signal_8106, new_AGEMA_signal_8105, subc_out[36]}), .a ({new_AGEMA_signal_8071, new_AGEMA_signal_8070, new_AGEMA_signal_8069, subc_out[52]}), .c ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8098, new_AGEMA_signal_8097, new_AGEMA_signal_8096, subc_out[40]}), .a ({new_AGEMA_signal_8062, new_AGEMA_signal_8061, new_AGEMA_signal_8060, subc_out[56]}), .c ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8089, new_AGEMA_signal_8088, new_AGEMA_signal_8087, subc_out[44]}), .a ({new_AGEMA_signal_10390, new_AGEMA_signal_10389, new_AGEMA_signal_10388, subc_out[60]}), .c ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8080, new_AGEMA_signal_8079, new_AGEMA_signal_8078, subc_out[48]}), .a ({new_AGEMA_signal_8116, new_AGEMA_signal_8115, new_AGEMA_signal_8114, subc_out[32]}), .c ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8071, new_AGEMA_signal_8070, new_AGEMA_signal_8069, subc_out[52]}), .a ({new_AGEMA_signal_8107, new_AGEMA_signal_8106, new_AGEMA_signal_8105, subc_out[36]}), .c ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8134, new_AGEMA_signal_8133, new_AGEMA_signal_8132, subc_out[20]}), .a ({new_AGEMA_signal_8170, new_AGEMA_signal_8169, new_AGEMA_signal_8168, subc_out[4]}), .c ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8125, new_AGEMA_signal_8124, new_AGEMA_signal_8123, subc_out[24]}), .a ({new_AGEMA_signal_8161, new_AGEMA_signal_8160, new_AGEMA_signal_8159, subc_out[8]}), .c ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10399, new_AGEMA_signal_10398, new_AGEMA_signal_10397, subc_out[28]}), .a ({new_AGEMA_signal_8152, new_AGEMA_signal_8151, new_AGEMA_signal_8150, subc_out[12]}), .c ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8179, new_AGEMA_signal_8178, new_AGEMA_signal_8177, subc_out[0]}), .a ({new_AGEMA_signal_8143, new_AGEMA_signal_8142, new_AGEMA_signal_8141, subc_out[16]}), .c ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8170, new_AGEMA_signal_8169, new_AGEMA_signal_8168, subc_out[4]}), .a ({new_AGEMA_signal_8134, new_AGEMA_signal_8133, new_AGEMA_signal_8132, subc_out[20]}), .c ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8161, new_AGEMA_signal_8160, new_AGEMA_signal_8159, subc_out[8]}), .a ({new_AGEMA_signal_8125, new_AGEMA_signal_8124, new_AGEMA_signal_8123, subc_out[24]}), .c ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8152, new_AGEMA_signal_8151, new_AGEMA_signal_8150, subc_out[12]}), .a ({new_AGEMA_signal_10399, new_AGEMA_signal_10398, new_AGEMA_signal_10397, subc_out[28]}), .c ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8143, new_AGEMA_signal_8142, new_AGEMA_signal_8141, subc_out[16]}), .a ({new_AGEMA_signal_8179, new_AGEMA_signal_8178, new_AGEMA_signal_8177, subc_out[0]}), .c ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_12808, new_AGEMA_signal_12807, new_AGEMA_signal_12806, add_sub1_0_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_10066, new_AGEMA_signal_10065, new_AGEMA_signal_10064, add_sub1_0_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_14254, new_AGEMA_signal_14253, new_AGEMA_signal_14252, subc_out[127]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_10369, new_AGEMA_signal_10368, new_AGEMA_signal_10367, add_sub1_0_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_10366, new_AGEMA_signal_10365, new_AGEMA_signal_10364, add_sub1_0_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_11356, new_AGEMA_signal_11355, new_AGEMA_signal_11354, subc_out[126]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_14257, new_AGEMA_signal_14256, new_AGEMA_signal_14255, add_sub1_0_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_9154, new_AGEMA_signal_9153, new_AGEMA_signal_9152, add_sub1_0_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_15682, new_AGEMA_signal_15681, new_AGEMA_signal_15680, subc_out[125]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_12808, new_AGEMA_signal_12807, new_AGEMA_signal_12806, add_sub1_0_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_9151, new_AGEMA_signal_9150, new_AGEMA_signal_9149, add_sub1_0_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_14257, new_AGEMA_signal_14256, new_AGEMA_signal_14255, add_sub1_0_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_11359, new_AGEMA_signal_11358, new_AGEMA_signal_11357, add_sub1_0_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_8440, new_AGEMA_signal_8439, new_AGEMA_signal_8438, add_sub1_0_addc_out[1]}), .c ({new_AGEMA_signal_12808, new_AGEMA_signal_12807, new_AGEMA_signal_12806, add_sub1_0_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_10369, new_AGEMA_signal_10368, new_AGEMA_signal_10367, add_sub1_0_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_10069, new_AGEMA_signal_10068, new_AGEMA_signal_10067, add_sub1_0_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_11359, new_AGEMA_signal_11358, new_AGEMA_signal_11357, add_sub1_0_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_10072, new_AGEMA_signal_10071, new_AGEMA_signal_10070, add_sub1_0_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_8434, new_AGEMA_signal_8433, new_AGEMA_signal_8432, add_sub1_0_addc_out[3]}), .c ({new_AGEMA_signal_10369, new_AGEMA_signal_10368, new_AGEMA_signal_10367, add_sub1_0_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_8443, new_AGEMA_signal_8442, new_AGEMA_signal_8441, add_sub1_0_addc_out[0]}), .b ({new_AGEMA_signal_9148, new_AGEMA_signal_9147, new_AGEMA_signal_9146, add_sub1_0_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_10069, new_AGEMA_signal_10068, new_AGEMA_signal_10067, add_sub1_0_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_9145, new_AGEMA_signal_9144, new_AGEMA_signal_9143, add_sub1_0_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_9157, new_AGEMA_signal_9156, new_AGEMA_signal_9155, add_sub1_0_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_10072, new_AGEMA_signal_10071, new_AGEMA_signal_10070, add_sub1_0_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_8446, new_AGEMA_signal_8445, new_AGEMA_signal_8444, add_sub1_0_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_7507, new_AGEMA_signal_7506, new_AGEMA_signal_7505, add_sub1_0_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_9163, new_AGEMA_signal_9162, new_AGEMA_signal_9161, subc_out[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_7933, new_AGEMA_signal_7932, new_AGEMA_signal_7931, add_sub1_0_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7930, new_AGEMA_signal_7929, new_AGEMA_signal_7928, add_sub1_0_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_8185, new_AGEMA_signal_8184, new_AGEMA_signal_8183, subc_out[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_9166, new_AGEMA_signal_9165, new_AGEMA_signal_9164, add_sub1_0_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_6904, new_AGEMA_signal_6903, new_AGEMA_signal_6902, add_sub1_0_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_10075, new_AGEMA_signal_10074, new_AGEMA_signal_10073, subc_out[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_8446, new_AGEMA_signal_8445, new_AGEMA_signal_8444, add_sub1_0_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_6901, new_AGEMA_signal_6900, new_AGEMA_signal_6899, add_sub1_0_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_9166, new_AGEMA_signal_9165, new_AGEMA_signal_9164, add_sub1_0_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_8188, new_AGEMA_signal_8187, new_AGEMA_signal_8186, add_sub1_0_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_6829, new_AGEMA_signal_6828, new_AGEMA_signal_6827, addc_in[121]}), .c ({new_AGEMA_signal_8446, new_AGEMA_signal_8445, new_AGEMA_signal_8444, add_sub1_0_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_7933, new_AGEMA_signal_7932, new_AGEMA_signal_7931, add_sub1_0_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7510, new_AGEMA_signal_7509, new_AGEMA_signal_7508, add_sub1_0_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_8188, new_AGEMA_signal_8187, new_AGEMA_signal_8186, add_sub1_0_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, new_AGEMA_signal_7511, add_sub1_0_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_6847, new_AGEMA_signal_6846, new_AGEMA_signal_6845, addc_in[123]}), .c ({new_AGEMA_signal_7933, new_AGEMA_signal_7932, new_AGEMA_signal_7931, add_sub1_0_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6820, new_AGEMA_signal_6819, new_AGEMA_signal_6818, addc_in[120]}), .b ({new_AGEMA_signal_6898, new_AGEMA_signal_6897, new_AGEMA_signal_6896, add_sub1_0_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_7510, new_AGEMA_signal_7509, new_AGEMA_signal_7508, add_sub1_0_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6895, new_AGEMA_signal_6894, new_AGEMA_signal_6893, add_sub1_0_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_6907, new_AGEMA_signal_6906, new_AGEMA_signal_6905, add_sub1_0_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_7513, new_AGEMA_signal_7512, new_AGEMA_signal_7511, add_sub1_0_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_8449, new_AGEMA_signal_8448, new_AGEMA_signal_8447, add_sub1_0_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_7522, new_AGEMA_signal_7521, new_AGEMA_signal_7520, add_sub1_0_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_9169, new_AGEMA_signal_9168, new_AGEMA_signal_9167, subc_out[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, new_AGEMA_signal_7940, add_sub1_0_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7939, new_AGEMA_signal_7938, new_AGEMA_signal_7937, add_sub1_0_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_8191, new_AGEMA_signal_8190, new_AGEMA_signal_8189, subc_out[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_9172, new_AGEMA_signal_9171, new_AGEMA_signal_9170, add_sub1_0_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_6925, new_AGEMA_signal_6924, new_AGEMA_signal_6923, add_sub1_0_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_10078, new_AGEMA_signal_10077, new_AGEMA_signal_10076, subc_out[117]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_8449, new_AGEMA_signal_8448, new_AGEMA_signal_8447, add_sub1_0_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_6922, new_AGEMA_signal_6921, new_AGEMA_signal_6920, add_sub1_0_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_9172, new_AGEMA_signal_9171, new_AGEMA_signal_9170, add_sub1_0_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_8194, new_AGEMA_signal_8193, new_AGEMA_signal_8192, add_sub1_0_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_6793, new_AGEMA_signal_6792, new_AGEMA_signal_6791, addc_in[117]}), .c ({new_AGEMA_signal_8449, new_AGEMA_signal_8448, new_AGEMA_signal_8447, add_sub1_0_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, new_AGEMA_signal_7940, add_sub1_0_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, new_AGEMA_signal_7523, add_sub1_0_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_8194, new_AGEMA_signal_8193, new_AGEMA_signal_8192, add_sub1_0_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_7528, new_AGEMA_signal_7527, new_AGEMA_signal_7526, add_sub1_0_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_6811, new_AGEMA_signal_6810, new_AGEMA_signal_6809, addc_in[119]}), .c ({new_AGEMA_signal_7942, new_AGEMA_signal_7941, new_AGEMA_signal_7940, add_sub1_0_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6784, new_AGEMA_signal_6783, new_AGEMA_signal_6782, addc_in[116]}), .b ({new_AGEMA_signal_6919, new_AGEMA_signal_6918, new_AGEMA_signal_6917, add_sub1_0_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_7525, new_AGEMA_signal_7524, new_AGEMA_signal_7523, add_sub1_0_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6916, new_AGEMA_signal_6915, new_AGEMA_signal_6914, add_sub1_0_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_6928, new_AGEMA_signal_6927, new_AGEMA_signal_6926, add_sub1_0_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_7528, new_AGEMA_signal_7527, new_AGEMA_signal_7526, add_sub1_0_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_8452, new_AGEMA_signal_8451, new_AGEMA_signal_8450, add_sub1_0_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_7537, new_AGEMA_signal_7536, new_AGEMA_signal_7535, add_sub1_0_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_9175, new_AGEMA_signal_9174, new_AGEMA_signal_9173, subc_out[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_7951, new_AGEMA_signal_7950, new_AGEMA_signal_7949, add_sub1_0_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7948, new_AGEMA_signal_7947, new_AGEMA_signal_7946, add_sub1_0_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_8197, new_AGEMA_signal_8196, new_AGEMA_signal_8195, subc_out[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_9178, new_AGEMA_signal_9177, new_AGEMA_signal_9176, add_sub1_0_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_6946, new_AGEMA_signal_6945, new_AGEMA_signal_6944, add_sub1_0_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_10081, new_AGEMA_signal_10080, new_AGEMA_signal_10079, subc_out[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_8452, new_AGEMA_signal_8451, new_AGEMA_signal_8450, add_sub1_0_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_6943, new_AGEMA_signal_6942, new_AGEMA_signal_6941, add_sub1_0_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_9178, new_AGEMA_signal_9177, new_AGEMA_signal_9176, add_sub1_0_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_8200, new_AGEMA_signal_8199, new_AGEMA_signal_8198, add_sub1_0_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_6757, new_AGEMA_signal_6756, new_AGEMA_signal_6755, addc_in[113]}), .c ({new_AGEMA_signal_8452, new_AGEMA_signal_8451, new_AGEMA_signal_8450, add_sub1_0_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_7951, new_AGEMA_signal_7950, new_AGEMA_signal_7949, add_sub1_0_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7540, new_AGEMA_signal_7539, new_AGEMA_signal_7538, add_sub1_0_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_8200, new_AGEMA_signal_8199, new_AGEMA_signal_8198, add_sub1_0_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_7543, new_AGEMA_signal_7542, new_AGEMA_signal_7541, add_sub1_0_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_6775, new_AGEMA_signal_6774, new_AGEMA_signal_6773, addc_in[115]}), .c ({new_AGEMA_signal_7951, new_AGEMA_signal_7950, new_AGEMA_signal_7949, add_sub1_0_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6748, new_AGEMA_signal_6747, new_AGEMA_signal_6746, addc_in[112]}), .b ({new_AGEMA_signal_6940, new_AGEMA_signal_6939, new_AGEMA_signal_6938, add_sub1_0_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_7540, new_AGEMA_signal_7539, new_AGEMA_signal_7538, add_sub1_0_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6937, new_AGEMA_signal_6936, new_AGEMA_signal_6935, add_sub1_0_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_6949, new_AGEMA_signal_6948, new_AGEMA_signal_6947, add_sub1_0_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_7543, new_AGEMA_signal_7542, new_AGEMA_signal_7541, add_sub1_0_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_8455, new_AGEMA_signal_8454, new_AGEMA_signal_8453, add_sub1_0_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_7552, new_AGEMA_signal_7551, new_AGEMA_signal_7550, add_sub1_0_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_9181, new_AGEMA_signal_9180, new_AGEMA_signal_9179, subc_out[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, new_AGEMA_signal_7958, add_sub1_0_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7957, new_AGEMA_signal_7956, new_AGEMA_signal_7955, add_sub1_0_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_8203, new_AGEMA_signal_8202, new_AGEMA_signal_8201, subc_out[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_9184, new_AGEMA_signal_9183, new_AGEMA_signal_9182, add_sub1_0_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_6967, new_AGEMA_signal_6966, new_AGEMA_signal_6965, add_sub1_0_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_10084, new_AGEMA_signal_10083, new_AGEMA_signal_10082, subc_out[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_8455, new_AGEMA_signal_8454, new_AGEMA_signal_8453, add_sub1_0_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_6964, new_AGEMA_signal_6963, new_AGEMA_signal_6962, add_sub1_0_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_9184, new_AGEMA_signal_9183, new_AGEMA_signal_9182, add_sub1_0_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_8206, new_AGEMA_signal_8205, new_AGEMA_signal_8204, add_sub1_0_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_6721, new_AGEMA_signal_6720, new_AGEMA_signal_6719, addc_in[109]}), .c ({new_AGEMA_signal_8455, new_AGEMA_signal_8454, new_AGEMA_signal_8453, add_sub1_0_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, new_AGEMA_signal_7958, add_sub1_0_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7555, new_AGEMA_signal_7554, new_AGEMA_signal_7553, add_sub1_0_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_8206, new_AGEMA_signal_8205, new_AGEMA_signal_8204, add_sub1_0_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_7558, new_AGEMA_signal_7557, new_AGEMA_signal_7556, add_sub1_0_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_6739, new_AGEMA_signal_6738, new_AGEMA_signal_6737, addc_in[111]}), .c ({new_AGEMA_signal_7960, new_AGEMA_signal_7959, new_AGEMA_signal_7958, add_sub1_0_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6712, new_AGEMA_signal_6711, new_AGEMA_signal_6710, addc_in[108]}), .b ({new_AGEMA_signal_6961, new_AGEMA_signal_6960, new_AGEMA_signal_6959, add_sub1_0_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_7555, new_AGEMA_signal_7554, new_AGEMA_signal_7553, add_sub1_0_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6958, new_AGEMA_signal_6957, new_AGEMA_signal_6956, add_sub1_0_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_6970, new_AGEMA_signal_6969, new_AGEMA_signal_6968, add_sub1_0_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_7558, new_AGEMA_signal_7557, new_AGEMA_signal_7556, add_sub1_0_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_8458, new_AGEMA_signal_8457, new_AGEMA_signal_8456, add_sub1_0_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_7567, new_AGEMA_signal_7566, new_AGEMA_signal_7565, add_sub1_0_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_9187, new_AGEMA_signal_9186, new_AGEMA_signal_9185, subc_out[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_7969, new_AGEMA_signal_7968, new_AGEMA_signal_7967, add_sub1_0_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7966, new_AGEMA_signal_7965, new_AGEMA_signal_7964, add_sub1_0_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_8209, new_AGEMA_signal_8208, new_AGEMA_signal_8207, subc_out[106]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_9190, new_AGEMA_signal_9189, new_AGEMA_signal_9188, add_sub1_0_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_6988, new_AGEMA_signal_6987, new_AGEMA_signal_6986, add_sub1_0_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_10087, new_AGEMA_signal_10086, new_AGEMA_signal_10085, subc_out[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_8458, new_AGEMA_signal_8457, new_AGEMA_signal_8456, add_sub1_0_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_6985, new_AGEMA_signal_6984, new_AGEMA_signal_6983, add_sub1_0_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_9190, new_AGEMA_signal_9189, new_AGEMA_signal_9188, add_sub1_0_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_8212, new_AGEMA_signal_8211, new_AGEMA_signal_8210, add_sub1_0_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_6685, new_AGEMA_signal_6684, new_AGEMA_signal_6683, addc_in[105]}), .c ({new_AGEMA_signal_8458, new_AGEMA_signal_8457, new_AGEMA_signal_8456, add_sub1_0_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_7969, new_AGEMA_signal_7968, new_AGEMA_signal_7967, add_sub1_0_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7570, new_AGEMA_signal_7569, new_AGEMA_signal_7568, add_sub1_0_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_8212, new_AGEMA_signal_8211, new_AGEMA_signal_8210, add_sub1_0_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_7573, new_AGEMA_signal_7572, new_AGEMA_signal_7571, add_sub1_0_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_6703, new_AGEMA_signal_6702, new_AGEMA_signal_6701, addc_in[107]}), .c ({new_AGEMA_signal_7969, new_AGEMA_signal_7968, new_AGEMA_signal_7967, add_sub1_0_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6676, new_AGEMA_signal_6675, new_AGEMA_signal_6674, addc_in[104]}), .b ({new_AGEMA_signal_6982, new_AGEMA_signal_6981, new_AGEMA_signal_6980, add_sub1_0_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_7570, new_AGEMA_signal_7569, new_AGEMA_signal_7568, add_sub1_0_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_6979, new_AGEMA_signal_6978, new_AGEMA_signal_6977, add_sub1_0_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_6991, new_AGEMA_signal_6990, new_AGEMA_signal_6989, add_sub1_0_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_7573, new_AGEMA_signal_7572, new_AGEMA_signal_7571, add_sub1_0_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_8461, new_AGEMA_signal_8460, new_AGEMA_signal_8459, add_sub1_0_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7582, new_AGEMA_signal_7581, new_AGEMA_signal_7580, add_sub1_0_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_9193, new_AGEMA_signal_9192, new_AGEMA_signal_9191, subc_out[103]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, new_AGEMA_signal_7976, add_sub1_0_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7975, new_AGEMA_signal_7974, new_AGEMA_signal_7973, add_sub1_0_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_8215, new_AGEMA_signal_8214, new_AGEMA_signal_8213, subc_out[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_9196, new_AGEMA_signal_9195, new_AGEMA_signal_9194, add_sub1_0_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_7009, new_AGEMA_signal_7008, new_AGEMA_signal_7007, add_sub1_0_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, new_AGEMA_signal_10088, subc_out[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_8461, new_AGEMA_signal_8460, new_AGEMA_signal_8459, add_sub1_0_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7006, new_AGEMA_signal_7005, new_AGEMA_signal_7004, add_sub1_0_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_9196, new_AGEMA_signal_9195, new_AGEMA_signal_9194, add_sub1_0_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_8218, new_AGEMA_signal_8217, new_AGEMA_signal_8216, add_sub1_0_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_6649, new_AGEMA_signal_6648, new_AGEMA_signal_6647, addc_in[101]}), .c ({new_AGEMA_signal_8461, new_AGEMA_signal_8460, new_AGEMA_signal_8459, add_sub1_0_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, new_AGEMA_signal_7976, add_sub1_0_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7585, new_AGEMA_signal_7584, new_AGEMA_signal_7583, add_sub1_0_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_8218, new_AGEMA_signal_8217, new_AGEMA_signal_8216, add_sub1_0_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_7588, new_AGEMA_signal_7587, new_AGEMA_signal_7586, add_sub1_0_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_6667, new_AGEMA_signal_6666, new_AGEMA_signal_6665, addc_in[103]}), .c ({new_AGEMA_signal_7978, new_AGEMA_signal_7977, new_AGEMA_signal_7976, add_sub1_0_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6640, new_AGEMA_signal_6639, new_AGEMA_signal_6638, addc_in[100]}), .b ({new_AGEMA_signal_7003, new_AGEMA_signal_7002, new_AGEMA_signal_7001, add_sub1_0_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_7585, new_AGEMA_signal_7584, new_AGEMA_signal_7583, add_sub1_0_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7000, new_AGEMA_signal_6999, new_AGEMA_signal_6998, add_sub1_0_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_7012, new_AGEMA_signal_7011, new_AGEMA_signal_7010, add_sub1_0_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_7588, new_AGEMA_signal_7587, new_AGEMA_signal_7586, add_sub1_0_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_8464, new_AGEMA_signal_8463, new_AGEMA_signal_8462, add_sub1_0_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7597, new_AGEMA_signal_7596, new_AGEMA_signal_7595, add_sub1_0_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_9199, new_AGEMA_signal_9198, new_AGEMA_signal_9197, subc_out[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_7987, new_AGEMA_signal_7986, new_AGEMA_signal_7985, add_sub1_0_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7984, new_AGEMA_signal_7983, new_AGEMA_signal_7982, add_sub1_0_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_8221, new_AGEMA_signal_8220, new_AGEMA_signal_8219, subc_out[98]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_9202, new_AGEMA_signal_9201, new_AGEMA_signal_9200, add_sub1_0_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_7030, new_AGEMA_signal_7029, new_AGEMA_signal_7028, add_sub1_0_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_10093, new_AGEMA_signal_10092, new_AGEMA_signal_10091, subc_out[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_8464, new_AGEMA_signal_8463, new_AGEMA_signal_8462, add_sub1_0_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7027, new_AGEMA_signal_7026, new_AGEMA_signal_7025, add_sub1_0_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_9202, new_AGEMA_signal_9201, new_AGEMA_signal_9200, add_sub1_0_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_8224, new_AGEMA_signal_8223, new_AGEMA_signal_8222, add_sub1_0_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_6613, new_AGEMA_signal_6612, new_AGEMA_signal_6611, addc_in[97]}), .c ({new_AGEMA_signal_8464, new_AGEMA_signal_8463, new_AGEMA_signal_8462, add_sub1_0_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_7987, new_AGEMA_signal_7986, new_AGEMA_signal_7985, add_sub1_0_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7600, new_AGEMA_signal_7599, new_AGEMA_signal_7598, add_sub1_0_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_8224, new_AGEMA_signal_8223, new_AGEMA_signal_8222, add_sub1_0_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_7603, new_AGEMA_signal_7602, new_AGEMA_signal_7601, add_sub1_0_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_6631, new_AGEMA_signal_6630, new_AGEMA_signal_6629, addc_in[99]}), .c ({new_AGEMA_signal_7987, new_AGEMA_signal_7986, new_AGEMA_signal_7985, add_sub1_0_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6604, new_AGEMA_signal_6603, new_AGEMA_signal_6602, addc_in[96]}), .b ({new_AGEMA_signal_7024, new_AGEMA_signal_7023, new_AGEMA_signal_7022, add_sub1_0_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_7600, new_AGEMA_signal_7599, new_AGEMA_signal_7598, add_sub1_0_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_0_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7021, new_AGEMA_signal_7020, new_AGEMA_signal_7019, add_sub1_0_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_7033, new_AGEMA_signal_7032, new_AGEMA_signal_7031, add_sub1_0_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_7603, new_AGEMA_signal_7602, new_AGEMA_signal_7601, add_sub1_0_subc_rom_sbox_0_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_12811, new_AGEMA_signal_12810, new_AGEMA_signal_12809, add_sub1_1_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_10102, new_AGEMA_signal_10101, new_AGEMA_signal_10100, add_sub1_1_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_14260, new_AGEMA_signal_14259, new_AGEMA_signal_14258, subc_out[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, new_AGEMA_signal_10376, add_sub1_1_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_10375, new_AGEMA_signal_10374, new_AGEMA_signal_10373, add_sub1_1_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_11362, new_AGEMA_signal_11361, new_AGEMA_signal_11360, subc_out[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_14263, new_AGEMA_signal_14262, new_AGEMA_signal_14261, add_sub1_1_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_9217, new_AGEMA_signal_9216, new_AGEMA_signal_9215, add_sub1_1_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_15685, new_AGEMA_signal_15684, new_AGEMA_signal_15683, subc_out[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_12811, new_AGEMA_signal_12810, new_AGEMA_signal_12809, add_sub1_1_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_9214, new_AGEMA_signal_9213, new_AGEMA_signal_9212, add_sub1_1_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_14263, new_AGEMA_signal_14262, new_AGEMA_signal_14261, add_sub1_1_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_11365, new_AGEMA_signal_11364, new_AGEMA_signal_11363, add_sub1_1_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_8473, new_AGEMA_signal_8472, new_AGEMA_signal_8471, add_sub1_1_addc_out[1]}), .c ({new_AGEMA_signal_12811, new_AGEMA_signal_12810, new_AGEMA_signal_12809, add_sub1_1_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, new_AGEMA_signal_10376, add_sub1_1_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_10105, new_AGEMA_signal_10104, new_AGEMA_signal_10103, add_sub1_1_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_11365, new_AGEMA_signal_11364, new_AGEMA_signal_11363, add_sub1_1_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_10108, new_AGEMA_signal_10107, new_AGEMA_signal_10106, add_sub1_1_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_8467, new_AGEMA_signal_8466, new_AGEMA_signal_8465, add_sub1_1_addc_out[3]}), .c ({new_AGEMA_signal_10378, new_AGEMA_signal_10377, new_AGEMA_signal_10376, add_sub1_1_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_8476, new_AGEMA_signal_8475, new_AGEMA_signal_8474, add_sub1_1_addc_out[0]}), .b ({new_AGEMA_signal_9211, new_AGEMA_signal_9210, new_AGEMA_signal_9209, add_sub1_1_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_10105, new_AGEMA_signal_10104, new_AGEMA_signal_10103, add_sub1_1_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_9208, new_AGEMA_signal_9207, new_AGEMA_signal_9206, add_sub1_1_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_9220, new_AGEMA_signal_9219, new_AGEMA_signal_9218, add_sub1_1_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_10108, new_AGEMA_signal_10107, new_AGEMA_signal_10106, add_sub1_1_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_8479, new_AGEMA_signal_8478, new_AGEMA_signal_8477, add_sub1_1_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_7615, new_AGEMA_signal_7614, new_AGEMA_signal_7613, add_sub1_1_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_9226, new_AGEMA_signal_9225, new_AGEMA_signal_9224, subc_out[91]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, new_AGEMA_signal_7994, add_sub1_1_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7993, new_AGEMA_signal_7992, new_AGEMA_signal_7991, add_sub1_1_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_8230, new_AGEMA_signal_8229, new_AGEMA_signal_8228, subc_out[90]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_9229, new_AGEMA_signal_9228, new_AGEMA_signal_9227, add_sub1_1_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_7057, new_AGEMA_signal_7056, new_AGEMA_signal_7055, add_sub1_1_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_10111, new_AGEMA_signal_10110, new_AGEMA_signal_10109, subc_out[89]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_8479, new_AGEMA_signal_8478, new_AGEMA_signal_8477, add_sub1_1_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_7054, new_AGEMA_signal_7053, new_AGEMA_signal_7052, add_sub1_1_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_9229, new_AGEMA_signal_9228, new_AGEMA_signal_9227, add_sub1_1_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_8233, new_AGEMA_signal_8232, new_AGEMA_signal_8231, add_sub1_1_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_6541, new_AGEMA_signal_6540, new_AGEMA_signal_6539, addc_in[89]}), .c ({new_AGEMA_signal_8479, new_AGEMA_signal_8478, new_AGEMA_signal_8477, add_sub1_1_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, new_AGEMA_signal_7994, add_sub1_1_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7618, new_AGEMA_signal_7617, new_AGEMA_signal_7616, add_sub1_1_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_8233, new_AGEMA_signal_8232, new_AGEMA_signal_8231, add_sub1_1_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, new_AGEMA_signal_7619, add_sub1_1_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_6559, new_AGEMA_signal_6558, new_AGEMA_signal_6557, addc_in[91]}), .c ({new_AGEMA_signal_7996, new_AGEMA_signal_7995, new_AGEMA_signal_7994, add_sub1_1_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6532, new_AGEMA_signal_6531, new_AGEMA_signal_6530, addc_in[88]}), .b ({new_AGEMA_signal_7051, new_AGEMA_signal_7050, new_AGEMA_signal_7049, add_sub1_1_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_7618, new_AGEMA_signal_7617, new_AGEMA_signal_7616, add_sub1_1_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7048, new_AGEMA_signal_7047, new_AGEMA_signal_7046, add_sub1_1_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_7060, new_AGEMA_signal_7059, new_AGEMA_signal_7058, add_sub1_1_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_7621, new_AGEMA_signal_7620, new_AGEMA_signal_7619, add_sub1_1_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_8482, new_AGEMA_signal_8481, new_AGEMA_signal_8480, add_sub1_1_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_7630, new_AGEMA_signal_7629, new_AGEMA_signal_7628, add_sub1_1_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_9232, new_AGEMA_signal_9231, new_AGEMA_signal_9230, subc_out[87]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_8005, new_AGEMA_signal_8004, new_AGEMA_signal_8003, add_sub1_1_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_8002, new_AGEMA_signal_8001, new_AGEMA_signal_8000, add_sub1_1_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_8236, new_AGEMA_signal_8235, new_AGEMA_signal_8234, subc_out[86]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_9235, new_AGEMA_signal_9234, new_AGEMA_signal_9233, add_sub1_1_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_7078, new_AGEMA_signal_7077, new_AGEMA_signal_7076, add_sub1_1_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_10114, new_AGEMA_signal_10113, new_AGEMA_signal_10112, subc_out[85]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_8482, new_AGEMA_signal_8481, new_AGEMA_signal_8480, add_sub1_1_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_7075, new_AGEMA_signal_7074, new_AGEMA_signal_7073, add_sub1_1_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_9235, new_AGEMA_signal_9234, new_AGEMA_signal_9233, add_sub1_1_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_8239, new_AGEMA_signal_8238, new_AGEMA_signal_8237, add_sub1_1_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_6505, new_AGEMA_signal_6504, new_AGEMA_signal_6503, addc_in[85]}), .c ({new_AGEMA_signal_8482, new_AGEMA_signal_8481, new_AGEMA_signal_8480, add_sub1_1_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_8005, new_AGEMA_signal_8004, new_AGEMA_signal_8003, add_sub1_1_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, new_AGEMA_signal_7631, add_sub1_1_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_8239, new_AGEMA_signal_8238, new_AGEMA_signal_8237, add_sub1_1_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_7636, new_AGEMA_signal_7635, new_AGEMA_signal_7634, add_sub1_1_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_6523, new_AGEMA_signal_6522, new_AGEMA_signal_6521, addc_in[87]}), .c ({new_AGEMA_signal_8005, new_AGEMA_signal_8004, new_AGEMA_signal_8003, add_sub1_1_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6496, new_AGEMA_signal_6495, new_AGEMA_signal_6494, addc_in[84]}), .b ({new_AGEMA_signal_7072, new_AGEMA_signal_7071, new_AGEMA_signal_7070, add_sub1_1_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_7633, new_AGEMA_signal_7632, new_AGEMA_signal_7631, add_sub1_1_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7069, new_AGEMA_signal_7068, new_AGEMA_signal_7067, add_sub1_1_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_7081, new_AGEMA_signal_7080, new_AGEMA_signal_7079, add_sub1_1_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_7636, new_AGEMA_signal_7635, new_AGEMA_signal_7634, add_sub1_1_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_8485, new_AGEMA_signal_8484, new_AGEMA_signal_8483, add_sub1_1_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_7645, new_AGEMA_signal_7644, new_AGEMA_signal_7643, add_sub1_1_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_9238, new_AGEMA_signal_9237, new_AGEMA_signal_9236, subc_out[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_8014, new_AGEMA_signal_8013, new_AGEMA_signal_8012, add_sub1_1_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_8011, new_AGEMA_signal_8010, new_AGEMA_signal_8009, add_sub1_1_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_8242, new_AGEMA_signal_8241, new_AGEMA_signal_8240, subc_out[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_9241, new_AGEMA_signal_9240, new_AGEMA_signal_9239, add_sub1_1_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_7099, new_AGEMA_signal_7098, new_AGEMA_signal_7097, add_sub1_1_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_10117, new_AGEMA_signal_10116, new_AGEMA_signal_10115, subc_out[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_8485, new_AGEMA_signal_8484, new_AGEMA_signal_8483, add_sub1_1_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_7096, new_AGEMA_signal_7095, new_AGEMA_signal_7094, add_sub1_1_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_9241, new_AGEMA_signal_9240, new_AGEMA_signal_9239, add_sub1_1_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_8245, new_AGEMA_signal_8244, new_AGEMA_signal_8243, add_sub1_1_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_6469, new_AGEMA_signal_6468, new_AGEMA_signal_6467, addc_in[81]}), .c ({new_AGEMA_signal_8485, new_AGEMA_signal_8484, new_AGEMA_signal_8483, add_sub1_1_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_8014, new_AGEMA_signal_8013, new_AGEMA_signal_8012, add_sub1_1_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7648, new_AGEMA_signal_7647, new_AGEMA_signal_7646, add_sub1_1_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_8245, new_AGEMA_signal_8244, new_AGEMA_signal_8243, add_sub1_1_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, new_AGEMA_signal_7649, add_sub1_1_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_6487, new_AGEMA_signal_6486, new_AGEMA_signal_6485, addc_in[83]}), .c ({new_AGEMA_signal_8014, new_AGEMA_signal_8013, new_AGEMA_signal_8012, add_sub1_1_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6460, new_AGEMA_signal_6459, new_AGEMA_signal_6458, addc_in[80]}), .b ({new_AGEMA_signal_7093, new_AGEMA_signal_7092, new_AGEMA_signal_7091, add_sub1_1_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_7648, new_AGEMA_signal_7647, new_AGEMA_signal_7646, add_sub1_1_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7090, new_AGEMA_signal_7089, new_AGEMA_signal_7088, add_sub1_1_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_7102, new_AGEMA_signal_7101, new_AGEMA_signal_7100, add_sub1_1_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_7651, new_AGEMA_signal_7650, new_AGEMA_signal_7649, add_sub1_1_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_8488, new_AGEMA_signal_8487, new_AGEMA_signal_8486, add_sub1_1_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_7660, new_AGEMA_signal_7659, new_AGEMA_signal_7658, add_sub1_1_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_9244, new_AGEMA_signal_9243, new_AGEMA_signal_9242, subc_out[79]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_8023, new_AGEMA_signal_8022, new_AGEMA_signal_8021, add_sub1_1_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_8020, new_AGEMA_signal_8019, new_AGEMA_signal_8018, add_sub1_1_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_8248, new_AGEMA_signal_8247, new_AGEMA_signal_8246, subc_out[78]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_9247, new_AGEMA_signal_9246, new_AGEMA_signal_9245, add_sub1_1_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_7120, new_AGEMA_signal_7119, new_AGEMA_signal_7118, add_sub1_1_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_10120, new_AGEMA_signal_10119, new_AGEMA_signal_10118, subc_out[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_8488, new_AGEMA_signal_8487, new_AGEMA_signal_8486, add_sub1_1_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_7117, new_AGEMA_signal_7116, new_AGEMA_signal_7115, add_sub1_1_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_9247, new_AGEMA_signal_9246, new_AGEMA_signal_9245, add_sub1_1_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_8251, new_AGEMA_signal_8250, new_AGEMA_signal_8249, add_sub1_1_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_6433, new_AGEMA_signal_6432, new_AGEMA_signal_6431, addc_in[77]}), .c ({new_AGEMA_signal_8488, new_AGEMA_signal_8487, new_AGEMA_signal_8486, add_sub1_1_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_8023, new_AGEMA_signal_8022, new_AGEMA_signal_8021, add_sub1_1_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, new_AGEMA_signal_7661, add_sub1_1_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_8251, new_AGEMA_signal_8250, new_AGEMA_signal_8249, add_sub1_1_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_7666, new_AGEMA_signal_7665, new_AGEMA_signal_7664, add_sub1_1_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_6451, new_AGEMA_signal_6450, new_AGEMA_signal_6449, addc_in[79]}), .c ({new_AGEMA_signal_8023, new_AGEMA_signal_8022, new_AGEMA_signal_8021, add_sub1_1_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6424, new_AGEMA_signal_6423, new_AGEMA_signal_6422, addc_in[76]}), .b ({new_AGEMA_signal_7114, new_AGEMA_signal_7113, new_AGEMA_signal_7112, add_sub1_1_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_7663, new_AGEMA_signal_7662, new_AGEMA_signal_7661, add_sub1_1_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7111, new_AGEMA_signal_7110, new_AGEMA_signal_7109, add_sub1_1_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_7123, new_AGEMA_signal_7122, new_AGEMA_signal_7121, add_sub1_1_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_7666, new_AGEMA_signal_7665, new_AGEMA_signal_7664, add_sub1_1_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_8491, new_AGEMA_signal_8490, new_AGEMA_signal_8489, add_sub1_1_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_7675, new_AGEMA_signal_7674, new_AGEMA_signal_7673, add_sub1_1_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_9250, new_AGEMA_signal_9249, new_AGEMA_signal_9248, subc_out[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_8032, new_AGEMA_signal_8031, new_AGEMA_signal_8030, add_sub1_1_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_8029, new_AGEMA_signal_8028, new_AGEMA_signal_8027, add_sub1_1_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_8254, new_AGEMA_signal_8253, new_AGEMA_signal_8252, subc_out[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_9253, new_AGEMA_signal_9252, new_AGEMA_signal_9251, add_sub1_1_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_7141, new_AGEMA_signal_7140, new_AGEMA_signal_7139, add_sub1_1_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_10123, new_AGEMA_signal_10122, new_AGEMA_signal_10121, subc_out[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_8491, new_AGEMA_signal_8490, new_AGEMA_signal_8489, add_sub1_1_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_7138, new_AGEMA_signal_7137, new_AGEMA_signal_7136, add_sub1_1_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_9253, new_AGEMA_signal_9252, new_AGEMA_signal_9251, add_sub1_1_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_8257, new_AGEMA_signal_8256, new_AGEMA_signal_8255, add_sub1_1_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_6397, new_AGEMA_signal_6396, new_AGEMA_signal_6395, addc_in[73]}), .c ({new_AGEMA_signal_8491, new_AGEMA_signal_8490, new_AGEMA_signal_8489, add_sub1_1_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_8032, new_AGEMA_signal_8031, new_AGEMA_signal_8030, add_sub1_1_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7678, new_AGEMA_signal_7677, new_AGEMA_signal_7676, add_sub1_1_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_8257, new_AGEMA_signal_8256, new_AGEMA_signal_8255, add_sub1_1_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_7681, new_AGEMA_signal_7680, new_AGEMA_signal_7679, add_sub1_1_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_6415, new_AGEMA_signal_6414, new_AGEMA_signal_6413, addc_in[75]}), .c ({new_AGEMA_signal_8032, new_AGEMA_signal_8031, new_AGEMA_signal_8030, add_sub1_1_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6388, new_AGEMA_signal_6387, new_AGEMA_signal_6386, addc_in[72]}), .b ({new_AGEMA_signal_7135, new_AGEMA_signal_7134, new_AGEMA_signal_7133, add_sub1_1_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_7678, new_AGEMA_signal_7677, new_AGEMA_signal_7676, add_sub1_1_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7132, new_AGEMA_signal_7131, new_AGEMA_signal_7130, add_sub1_1_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_7144, new_AGEMA_signal_7143, new_AGEMA_signal_7142, add_sub1_1_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_7681, new_AGEMA_signal_7680, new_AGEMA_signal_7679, add_sub1_1_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_8494, new_AGEMA_signal_8493, new_AGEMA_signal_8492, add_sub1_1_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7690, new_AGEMA_signal_7689, new_AGEMA_signal_7688, add_sub1_1_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_9256, new_AGEMA_signal_9255, new_AGEMA_signal_9254, subc_out[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_8041, new_AGEMA_signal_8040, new_AGEMA_signal_8039, add_sub1_1_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_8038, new_AGEMA_signal_8037, new_AGEMA_signal_8036, add_sub1_1_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_8260, new_AGEMA_signal_8259, new_AGEMA_signal_8258, subc_out[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_9259, new_AGEMA_signal_9258, new_AGEMA_signal_9257, add_sub1_1_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_7162, new_AGEMA_signal_7161, new_AGEMA_signal_7160, add_sub1_1_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_10126, new_AGEMA_signal_10125, new_AGEMA_signal_10124, subc_out[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_8494, new_AGEMA_signal_8493, new_AGEMA_signal_8492, add_sub1_1_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7159, new_AGEMA_signal_7158, new_AGEMA_signal_7157, add_sub1_1_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_9259, new_AGEMA_signal_9258, new_AGEMA_signal_9257, add_sub1_1_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_8263, new_AGEMA_signal_8262, new_AGEMA_signal_8261, add_sub1_1_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_6361, new_AGEMA_signal_6360, new_AGEMA_signal_6359, addc_in[69]}), .c ({new_AGEMA_signal_8494, new_AGEMA_signal_8493, new_AGEMA_signal_8492, add_sub1_1_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_8041, new_AGEMA_signal_8040, new_AGEMA_signal_8039, add_sub1_1_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7693, new_AGEMA_signal_7692, new_AGEMA_signal_7691, add_sub1_1_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_8263, new_AGEMA_signal_8262, new_AGEMA_signal_8261, add_sub1_1_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_7696, new_AGEMA_signal_7695, new_AGEMA_signal_7694, add_sub1_1_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_6379, new_AGEMA_signal_6378, new_AGEMA_signal_6377, addc_in[71]}), .c ({new_AGEMA_signal_8041, new_AGEMA_signal_8040, new_AGEMA_signal_8039, add_sub1_1_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6352, new_AGEMA_signal_6351, new_AGEMA_signal_6350, addc_in[68]}), .b ({new_AGEMA_signal_7156, new_AGEMA_signal_7155, new_AGEMA_signal_7154, add_sub1_1_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_7693, new_AGEMA_signal_7692, new_AGEMA_signal_7691, add_sub1_1_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7153, new_AGEMA_signal_7152, new_AGEMA_signal_7151, add_sub1_1_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_7165, new_AGEMA_signal_7164, new_AGEMA_signal_7163, add_sub1_1_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_7696, new_AGEMA_signal_7695, new_AGEMA_signal_7694, add_sub1_1_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_8497, new_AGEMA_signal_8496, new_AGEMA_signal_8495, add_sub1_1_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7705, new_AGEMA_signal_7704, new_AGEMA_signal_7703, add_sub1_1_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_9262, new_AGEMA_signal_9261, new_AGEMA_signal_9260, subc_out[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_8050, new_AGEMA_signal_8049, new_AGEMA_signal_8048, add_sub1_1_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_8047, new_AGEMA_signal_8046, new_AGEMA_signal_8045, add_sub1_1_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_8266, new_AGEMA_signal_8265, new_AGEMA_signal_8264, subc_out[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_9265, new_AGEMA_signal_9264, new_AGEMA_signal_9263, add_sub1_1_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_7183, new_AGEMA_signal_7182, new_AGEMA_signal_7181, add_sub1_1_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_10129, new_AGEMA_signal_10128, new_AGEMA_signal_10127, subc_out[65]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_8497, new_AGEMA_signal_8496, new_AGEMA_signal_8495, add_sub1_1_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7180, new_AGEMA_signal_7179, new_AGEMA_signal_7178, add_sub1_1_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_9265, new_AGEMA_signal_9264, new_AGEMA_signal_9263, add_sub1_1_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_8269, new_AGEMA_signal_8268, new_AGEMA_signal_8267, add_sub1_1_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_6325, new_AGEMA_signal_6324, new_AGEMA_signal_6323, addc_in[65]}), .c ({new_AGEMA_signal_8497, new_AGEMA_signal_8496, new_AGEMA_signal_8495, add_sub1_1_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_8050, new_AGEMA_signal_8049, new_AGEMA_signal_8048, add_sub1_1_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7708, new_AGEMA_signal_7707, new_AGEMA_signal_7706, add_sub1_1_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_8269, new_AGEMA_signal_8268, new_AGEMA_signal_8267, add_sub1_1_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_7711, new_AGEMA_signal_7710, new_AGEMA_signal_7709, add_sub1_1_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_6343, new_AGEMA_signal_6342, new_AGEMA_signal_6341, addc_in[67]}), .c ({new_AGEMA_signal_8050, new_AGEMA_signal_8049, new_AGEMA_signal_8048, add_sub1_1_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6316, new_AGEMA_signal_6315, new_AGEMA_signal_6314, addc_in[64]}), .b ({new_AGEMA_signal_7177, new_AGEMA_signal_7176, new_AGEMA_signal_7175, add_sub1_1_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_7708, new_AGEMA_signal_7707, new_AGEMA_signal_7706, add_sub1_1_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_1_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7174, new_AGEMA_signal_7173, new_AGEMA_signal_7172, add_sub1_1_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_7186, new_AGEMA_signal_7185, new_AGEMA_signal_7184, add_sub1_1_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_7711, new_AGEMA_signal_7710, new_AGEMA_signal_7709, add_sub1_1_subc_rom_sbox_0_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_12814, new_AGEMA_signal_12813, new_AGEMA_signal_12812, add_sub1_2_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_10138, new_AGEMA_signal_10137, new_AGEMA_signal_10136, add_sub1_2_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_14266, new_AGEMA_signal_14265, new_AGEMA_signal_14264, subc_out[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_10387, new_AGEMA_signal_10386, new_AGEMA_signal_10385, add_sub1_2_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_10384, new_AGEMA_signal_10383, new_AGEMA_signal_10382, add_sub1_2_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_11368, new_AGEMA_signal_11367, new_AGEMA_signal_11366, subc_out[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_14269, new_AGEMA_signal_14268, new_AGEMA_signal_14267, add_sub1_2_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_9280, new_AGEMA_signal_9279, new_AGEMA_signal_9278, add_sub1_2_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_15688, new_AGEMA_signal_15687, new_AGEMA_signal_15686, subc_out[61]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_12814, new_AGEMA_signal_12813, new_AGEMA_signal_12812, add_sub1_2_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_9277, new_AGEMA_signal_9276, new_AGEMA_signal_9275, add_sub1_2_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_14269, new_AGEMA_signal_14268, new_AGEMA_signal_14267, add_sub1_2_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_11371, new_AGEMA_signal_11370, new_AGEMA_signal_11369, add_sub1_2_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_8506, new_AGEMA_signal_8505, new_AGEMA_signal_8504, add_sub1_2_addc_out[1]}), .c ({new_AGEMA_signal_12814, new_AGEMA_signal_12813, new_AGEMA_signal_12812, add_sub1_2_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_10387, new_AGEMA_signal_10386, new_AGEMA_signal_10385, add_sub1_2_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_10141, new_AGEMA_signal_10140, new_AGEMA_signal_10139, add_sub1_2_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_11371, new_AGEMA_signal_11370, new_AGEMA_signal_11369, add_sub1_2_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_10144, new_AGEMA_signal_10143, new_AGEMA_signal_10142, add_sub1_2_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_8500, new_AGEMA_signal_8499, new_AGEMA_signal_8498, add_sub1_2_addc_out[3]}), .c ({new_AGEMA_signal_10387, new_AGEMA_signal_10386, new_AGEMA_signal_10385, add_sub1_2_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_8509, new_AGEMA_signal_8508, new_AGEMA_signal_8507, add_sub1_2_addc_out[0]}), .b ({new_AGEMA_signal_9274, new_AGEMA_signal_9273, new_AGEMA_signal_9272, add_sub1_2_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_10141, new_AGEMA_signal_10140, new_AGEMA_signal_10139, add_sub1_2_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_9271, new_AGEMA_signal_9270, new_AGEMA_signal_9269, add_sub1_2_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_9283, new_AGEMA_signal_9282, new_AGEMA_signal_9281, add_sub1_2_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_10144, new_AGEMA_signal_10143, new_AGEMA_signal_10142, add_sub1_2_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_8512, new_AGEMA_signal_8511, new_AGEMA_signal_8510, add_sub1_2_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_7723, new_AGEMA_signal_7722, new_AGEMA_signal_7721, add_sub1_2_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_9289, new_AGEMA_signal_9288, new_AGEMA_signal_9287, subc_out[59]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_8059, new_AGEMA_signal_8058, new_AGEMA_signal_8057, add_sub1_2_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_8056, new_AGEMA_signal_8055, new_AGEMA_signal_8054, add_sub1_2_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_8275, new_AGEMA_signal_8274, new_AGEMA_signal_8273, subc_out[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_9292, new_AGEMA_signal_9291, new_AGEMA_signal_9290, add_sub1_2_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_7210, new_AGEMA_signal_7209, new_AGEMA_signal_7208, add_sub1_2_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_10147, new_AGEMA_signal_10146, new_AGEMA_signal_10145, subc_out[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_8512, new_AGEMA_signal_8511, new_AGEMA_signal_8510, add_sub1_2_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_7207, new_AGEMA_signal_7206, new_AGEMA_signal_7205, add_sub1_2_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_9292, new_AGEMA_signal_9291, new_AGEMA_signal_9290, add_sub1_2_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_8278, new_AGEMA_signal_8277, new_AGEMA_signal_8276, add_sub1_2_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, new_AGEMA_signal_6251, addc_in[57]}), .c ({new_AGEMA_signal_8512, new_AGEMA_signal_8511, new_AGEMA_signal_8510, add_sub1_2_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_8059, new_AGEMA_signal_8058, new_AGEMA_signal_8057, add_sub1_2_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7726, new_AGEMA_signal_7725, new_AGEMA_signal_7724, add_sub1_2_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_8278, new_AGEMA_signal_8277, new_AGEMA_signal_8276, add_sub1_2_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_7729, new_AGEMA_signal_7728, new_AGEMA_signal_7727, add_sub1_2_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_6271, new_AGEMA_signal_6270, new_AGEMA_signal_6269, addc_in[59]}), .c ({new_AGEMA_signal_8059, new_AGEMA_signal_8058, new_AGEMA_signal_8057, add_sub1_2_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6244, new_AGEMA_signal_6243, new_AGEMA_signal_6242, addc_in[56]}), .b ({new_AGEMA_signal_7204, new_AGEMA_signal_7203, new_AGEMA_signal_7202, add_sub1_2_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_7726, new_AGEMA_signal_7725, new_AGEMA_signal_7724, add_sub1_2_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7201, new_AGEMA_signal_7200, new_AGEMA_signal_7199, add_sub1_2_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_7213, new_AGEMA_signal_7212, new_AGEMA_signal_7211, add_sub1_2_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_7729, new_AGEMA_signal_7728, new_AGEMA_signal_7727, add_sub1_2_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_8515, new_AGEMA_signal_8514, new_AGEMA_signal_8513, add_sub1_2_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_7738, new_AGEMA_signal_7737, new_AGEMA_signal_7736, add_sub1_2_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_9295, new_AGEMA_signal_9294, new_AGEMA_signal_9293, subc_out[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_8068, new_AGEMA_signal_8067, new_AGEMA_signal_8066, add_sub1_2_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_8065, new_AGEMA_signal_8064, new_AGEMA_signal_8063, add_sub1_2_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_8281, new_AGEMA_signal_8280, new_AGEMA_signal_8279, subc_out[54]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_9298, new_AGEMA_signal_9297, new_AGEMA_signal_9296, add_sub1_2_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_7231, new_AGEMA_signal_7230, new_AGEMA_signal_7229, add_sub1_2_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_10150, new_AGEMA_signal_10149, new_AGEMA_signal_10148, subc_out[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_8515, new_AGEMA_signal_8514, new_AGEMA_signal_8513, add_sub1_2_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_7228, new_AGEMA_signal_7227, new_AGEMA_signal_7226, add_sub1_2_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_9298, new_AGEMA_signal_9297, new_AGEMA_signal_9296, add_sub1_2_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_8284, new_AGEMA_signal_8283, new_AGEMA_signal_8282, add_sub1_2_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, new_AGEMA_signal_6215, addc_in[53]}), .c ({new_AGEMA_signal_8515, new_AGEMA_signal_8514, new_AGEMA_signal_8513, add_sub1_2_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_8068, new_AGEMA_signal_8067, new_AGEMA_signal_8066, add_sub1_2_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7741, new_AGEMA_signal_7740, new_AGEMA_signal_7739, add_sub1_2_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_8284, new_AGEMA_signal_8283, new_AGEMA_signal_8282, add_sub1_2_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_7744, new_AGEMA_signal_7743, new_AGEMA_signal_7742, add_sub1_2_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_6235, new_AGEMA_signal_6234, new_AGEMA_signal_6233, addc_in[55]}), .c ({new_AGEMA_signal_8068, new_AGEMA_signal_8067, new_AGEMA_signal_8066, add_sub1_2_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6208, new_AGEMA_signal_6207, new_AGEMA_signal_6206, addc_in[52]}), .b ({new_AGEMA_signal_7225, new_AGEMA_signal_7224, new_AGEMA_signal_7223, add_sub1_2_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_7741, new_AGEMA_signal_7740, new_AGEMA_signal_7739, add_sub1_2_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7222, new_AGEMA_signal_7221, new_AGEMA_signal_7220, add_sub1_2_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_7234, new_AGEMA_signal_7233, new_AGEMA_signal_7232, add_sub1_2_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_7744, new_AGEMA_signal_7743, new_AGEMA_signal_7742, add_sub1_2_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_8518, new_AGEMA_signal_8517, new_AGEMA_signal_8516, add_sub1_2_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_7753, new_AGEMA_signal_7752, new_AGEMA_signal_7751, add_sub1_2_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_9301, new_AGEMA_signal_9300, new_AGEMA_signal_9299, subc_out[51]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_8077, new_AGEMA_signal_8076, new_AGEMA_signal_8075, add_sub1_2_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_8074, new_AGEMA_signal_8073, new_AGEMA_signal_8072, add_sub1_2_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_8287, new_AGEMA_signal_8286, new_AGEMA_signal_8285, subc_out[50]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_9304, new_AGEMA_signal_9303, new_AGEMA_signal_9302, add_sub1_2_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_7252, new_AGEMA_signal_7251, new_AGEMA_signal_7250, add_sub1_2_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_10153, new_AGEMA_signal_10152, new_AGEMA_signal_10151, subc_out[49]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_8518, new_AGEMA_signal_8517, new_AGEMA_signal_8516, add_sub1_2_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_7249, new_AGEMA_signal_7248, new_AGEMA_signal_7247, add_sub1_2_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_9304, new_AGEMA_signal_9303, new_AGEMA_signal_9302, add_sub1_2_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_8290, new_AGEMA_signal_8289, new_AGEMA_signal_8288, add_sub1_2_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_6181, new_AGEMA_signal_6180, new_AGEMA_signal_6179, addc_in[49]}), .c ({new_AGEMA_signal_8518, new_AGEMA_signal_8517, new_AGEMA_signal_8516, add_sub1_2_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_8077, new_AGEMA_signal_8076, new_AGEMA_signal_8075, add_sub1_2_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7756, new_AGEMA_signal_7755, new_AGEMA_signal_7754, add_sub1_2_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_8290, new_AGEMA_signal_8289, new_AGEMA_signal_8288, add_sub1_2_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_7759, new_AGEMA_signal_7758, new_AGEMA_signal_7757, add_sub1_2_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, new_AGEMA_signal_6197, addc_in[51]}), .c ({new_AGEMA_signal_8077, new_AGEMA_signal_8076, new_AGEMA_signal_8075, add_sub1_2_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6172, new_AGEMA_signal_6171, new_AGEMA_signal_6170, addc_in[48]}), .b ({new_AGEMA_signal_7246, new_AGEMA_signal_7245, new_AGEMA_signal_7244, add_sub1_2_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_7756, new_AGEMA_signal_7755, new_AGEMA_signal_7754, add_sub1_2_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7243, new_AGEMA_signal_7242, new_AGEMA_signal_7241, add_sub1_2_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_7255, new_AGEMA_signal_7254, new_AGEMA_signal_7253, add_sub1_2_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_7759, new_AGEMA_signal_7758, new_AGEMA_signal_7757, add_sub1_2_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_8521, new_AGEMA_signal_8520, new_AGEMA_signal_8519, add_sub1_2_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_7768, new_AGEMA_signal_7767, new_AGEMA_signal_7766, add_sub1_2_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_9307, new_AGEMA_signal_9306, new_AGEMA_signal_9305, subc_out[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_8086, new_AGEMA_signal_8085, new_AGEMA_signal_8084, add_sub1_2_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_8083, new_AGEMA_signal_8082, new_AGEMA_signal_8081, add_sub1_2_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_8293, new_AGEMA_signal_8292, new_AGEMA_signal_8291, subc_out[46]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_9310, new_AGEMA_signal_9309, new_AGEMA_signal_9308, add_sub1_2_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_7273, new_AGEMA_signal_7272, new_AGEMA_signal_7271, add_sub1_2_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, new_AGEMA_signal_10154, subc_out[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_8521, new_AGEMA_signal_8520, new_AGEMA_signal_8519, add_sub1_2_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_7270, new_AGEMA_signal_7269, new_AGEMA_signal_7268, add_sub1_2_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_9310, new_AGEMA_signal_9309, new_AGEMA_signal_9308, add_sub1_2_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_8296, new_AGEMA_signal_8295, new_AGEMA_signal_8294, add_sub1_2_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_6145, new_AGEMA_signal_6144, new_AGEMA_signal_6143, addc_in[45]}), .c ({new_AGEMA_signal_8521, new_AGEMA_signal_8520, new_AGEMA_signal_8519, add_sub1_2_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_8086, new_AGEMA_signal_8085, new_AGEMA_signal_8084, add_sub1_2_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7771, new_AGEMA_signal_7770, new_AGEMA_signal_7769, add_sub1_2_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_8296, new_AGEMA_signal_8295, new_AGEMA_signal_8294, add_sub1_2_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_7774, new_AGEMA_signal_7773, new_AGEMA_signal_7772, add_sub1_2_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, new_AGEMA_signal_6161, addc_in[47]}), .c ({new_AGEMA_signal_8086, new_AGEMA_signal_8085, new_AGEMA_signal_8084, add_sub1_2_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6136, new_AGEMA_signal_6135, new_AGEMA_signal_6134, addc_in[44]}), .b ({new_AGEMA_signal_7267, new_AGEMA_signal_7266, new_AGEMA_signal_7265, add_sub1_2_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_7771, new_AGEMA_signal_7770, new_AGEMA_signal_7769, add_sub1_2_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7264, new_AGEMA_signal_7263, new_AGEMA_signal_7262, add_sub1_2_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_7276, new_AGEMA_signal_7275, new_AGEMA_signal_7274, add_sub1_2_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_7774, new_AGEMA_signal_7773, new_AGEMA_signal_7772, add_sub1_2_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_8524, new_AGEMA_signal_8523, new_AGEMA_signal_8522, add_sub1_2_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_7783, new_AGEMA_signal_7782, new_AGEMA_signal_7781, add_sub1_2_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_9313, new_AGEMA_signal_9312, new_AGEMA_signal_9311, subc_out[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_8095, new_AGEMA_signal_8094, new_AGEMA_signal_8093, add_sub1_2_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_8092, new_AGEMA_signal_8091, new_AGEMA_signal_8090, add_sub1_2_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_8299, new_AGEMA_signal_8298, new_AGEMA_signal_8297, subc_out[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_9316, new_AGEMA_signal_9315, new_AGEMA_signal_9314, add_sub1_2_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_7294, new_AGEMA_signal_7293, new_AGEMA_signal_7292, add_sub1_2_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_10159, new_AGEMA_signal_10158, new_AGEMA_signal_10157, subc_out[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_8524, new_AGEMA_signal_8523, new_AGEMA_signal_8522, add_sub1_2_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_7291, new_AGEMA_signal_7290, new_AGEMA_signal_7289, add_sub1_2_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_9316, new_AGEMA_signal_9315, new_AGEMA_signal_9314, add_sub1_2_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_8302, new_AGEMA_signal_8301, new_AGEMA_signal_8300, add_sub1_2_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_6109, new_AGEMA_signal_6108, new_AGEMA_signal_6107, addc_in[41]}), .c ({new_AGEMA_signal_8524, new_AGEMA_signal_8523, new_AGEMA_signal_8522, add_sub1_2_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_8095, new_AGEMA_signal_8094, new_AGEMA_signal_8093, add_sub1_2_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7786, new_AGEMA_signal_7785, new_AGEMA_signal_7784, add_sub1_2_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_8302, new_AGEMA_signal_8301, new_AGEMA_signal_8300, add_sub1_2_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_7789, new_AGEMA_signal_7788, new_AGEMA_signal_7787, add_sub1_2_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, new_AGEMA_signal_6125, addc_in[43]}), .c ({new_AGEMA_signal_8095, new_AGEMA_signal_8094, new_AGEMA_signal_8093, add_sub1_2_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6100, new_AGEMA_signal_6099, new_AGEMA_signal_6098, addc_in[40]}), .b ({new_AGEMA_signal_7288, new_AGEMA_signal_7287, new_AGEMA_signal_7286, add_sub1_2_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_7786, new_AGEMA_signal_7785, new_AGEMA_signal_7784, add_sub1_2_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7285, new_AGEMA_signal_7284, new_AGEMA_signal_7283, add_sub1_2_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_7297, new_AGEMA_signal_7296, new_AGEMA_signal_7295, add_sub1_2_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_7789, new_AGEMA_signal_7788, new_AGEMA_signal_7787, add_sub1_2_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_8527, new_AGEMA_signal_8526, new_AGEMA_signal_8525, add_sub1_2_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7798, new_AGEMA_signal_7797, new_AGEMA_signal_7796, add_sub1_2_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_9319, new_AGEMA_signal_9318, new_AGEMA_signal_9317, subc_out[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_8104, new_AGEMA_signal_8103, new_AGEMA_signal_8102, add_sub1_2_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_8101, new_AGEMA_signal_8100, new_AGEMA_signal_8099, add_sub1_2_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_8305, new_AGEMA_signal_8304, new_AGEMA_signal_8303, subc_out[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_9322, new_AGEMA_signal_9321, new_AGEMA_signal_9320, add_sub1_2_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_7315, new_AGEMA_signal_7314, new_AGEMA_signal_7313, add_sub1_2_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_10162, new_AGEMA_signal_10161, new_AGEMA_signal_10160, subc_out[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_8527, new_AGEMA_signal_8526, new_AGEMA_signal_8525, add_sub1_2_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7312, new_AGEMA_signal_7311, new_AGEMA_signal_7310, add_sub1_2_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_9322, new_AGEMA_signal_9321, new_AGEMA_signal_9320, add_sub1_2_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_8308, new_AGEMA_signal_8307, new_AGEMA_signal_8306, add_sub1_2_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, new_AGEMA_signal_6071, addc_in[37]}), .c ({new_AGEMA_signal_8527, new_AGEMA_signal_8526, new_AGEMA_signal_8525, add_sub1_2_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_8104, new_AGEMA_signal_8103, new_AGEMA_signal_8102, add_sub1_2_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7801, new_AGEMA_signal_7800, new_AGEMA_signal_7799, add_sub1_2_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_8308, new_AGEMA_signal_8307, new_AGEMA_signal_8306, add_sub1_2_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_7804, new_AGEMA_signal_7803, new_AGEMA_signal_7802, add_sub1_2_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, new_AGEMA_signal_6089, addc_in[39]}), .c ({new_AGEMA_signal_8104, new_AGEMA_signal_8103, new_AGEMA_signal_8102, add_sub1_2_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6064, new_AGEMA_signal_6063, new_AGEMA_signal_6062, addc_in[36]}), .b ({new_AGEMA_signal_7309, new_AGEMA_signal_7308, new_AGEMA_signal_7307, add_sub1_2_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_7801, new_AGEMA_signal_7800, new_AGEMA_signal_7799, add_sub1_2_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7306, new_AGEMA_signal_7305, new_AGEMA_signal_7304, add_sub1_2_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_7318, new_AGEMA_signal_7317, new_AGEMA_signal_7316, add_sub1_2_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_7804, new_AGEMA_signal_7803, new_AGEMA_signal_7802, add_sub1_2_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_8530, new_AGEMA_signal_8529, new_AGEMA_signal_8528, add_sub1_2_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7813, new_AGEMA_signal_7812, new_AGEMA_signal_7811, add_sub1_2_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_9325, new_AGEMA_signal_9324, new_AGEMA_signal_9323, subc_out[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_8113, new_AGEMA_signal_8112, new_AGEMA_signal_8111, add_sub1_2_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_8110, new_AGEMA_signal_8109, new_AGEMA_signal_8108, add_sub1_2_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_8311, new_AGEMA_signal_8310, new_AGEMA_signal_8309, subc_out[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_9328, new_AGEMA_signal_9327, new_AGEMA_signal_9326, add_sub1_2_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_7336, new_AGEMA_signal_7335, new_AGEMA_signal_7334, add_sub1_2_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_10165, new_AGEMA_signal_10164, new_AGEMA_signal_10163, subc_out[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_8530, new_AGEMA_signal_8529, new_AGEMA_signal_8528, add_sub1_2_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7333, new_AGEMA_signal_7332, new_AGEMA_signal_7331, add_sub1_2_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_9328, new_AGEMA_signal_9327, new_AGEMA_signal_9326, add_sub1_2_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_8314, new_AGEMA_signal_8313, new_AGEMA_signal_8312, add_sub1_2_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_6037, new_AGEMA_signal_6036, new_AGEMA_signal_6035, addc_in[33]}), .c ({new_AGEMA_signal_8530, new_AGEMA_signal_8529, new_AGEMA_signal_8528, add_sub1_2_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_8113, new_AGEMA_signal_8112, new_AGEMA_signal_8111, add_sub1_2_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7816, new_AGEMA_signal_7815, new_AGEMA_signal_7814, add_sub1_2_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_8314, new_AGEMA_signal_8313, new_AGEMA_signal_8312, add_sub1_2_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_7819, new_AGEMA_signal_7818, new_AGEMA_signal_7817, add_sub1_2_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, new_AGEMA_signal_6053, addc_in[35]}), .c ({new_AGEMA_signal_8113, new_AGEMA_signal_8112, new_AGEMA_signal_8111, add_sub1_2_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_6028, new_AGEMA_signal_6027, new_AGEMA_signal_6026, addc_in[32]}), .b ({new_AGEMA_signal_7330, new_AGEMA_signal_7329, new_AGEMA_signal_7328, add_sub1_2_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_7816, new_AGEMA_signal_7815, new_AGEMA_signal_7814, add_sub1_2_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_2_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7327, new_AGEMA_signal_7326, new_AGEMA_signal_7325, add_sub1_2_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_7339, new_AGEMA_signal_7338, new_AGEMA_signal_7337, add_sub1_2_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_7819, new_AGEMA_signal_7818, new_AGEMA_signal_7817, add_sub1_2_subc_rom_sbox_0_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U14 ( .a ({new_AGEMA_signal_12817, new_AGEMA_signal_12816, new_AGEMA_signal_12815, add_sub1_3_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_10174, new_AGEMA_signal_10173, new_AGEMA_signal_10172, add_sub1_3_subc_rom_sbox_7_ANF_2_n19}), .c ({new_AGEMA_signal_14272, new_AGEMA_signal_14271, new_AGEMA_signal_14270, subc_out[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U13 ( .a ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, new_AGEMA_signal_10394, add_sub1_3_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_10393, new_AGEMA_signal_10392, new_AGEMA_signal_10391, add_sub1_3_subc_rom_sbox_7_ANF_2_n17}), .c ({new_AGEMA_signal_11374, new_AGEMA_signal_11373, new_AGEMA_signal_11372, subc_out[30]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U9 ( .a ({new_AGEMA_signal_14275, new_AGEMA_signal_14274, new_AGEMA_signal_14273, add_sub1_3_subc_rom_sbox_7_ANF_2_n14}), .b ({new_AGEMA_signal_9343, new_AGEMA_signal_9342, new_AGEMA_signal_9341, add_sub1_3_subc_rom_sbox_7_ANF_2_t2}), .c ({new_AGEMA_signal_15691, new_AGEMA_signal_15690, new_AGEMA_signal_15689, subc_out[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U8 ( .a ({new_AGEMA_signal_12817, new_AGEMA_signal_12816, new_AGEMA_signal_12815, add_sub1_3_subc_rom_sbox_7_ANF_2_n20}), .b ({new_AGEMA_signal_9340, new_AGEMA_signal_9339, new_AGEMA_signal_9338, add_sub1_3_subc_rom_sbox_7_ANF_2_t1}), .c ({new_AGEMA_signal_14275, new_AGEMA_signal_14274, new_AGEMA_signal_14273, add_sub1_3_subc_rom_sbox_7_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U7 ( .a ({new_AGEMA_signal_11377, new_AGEMA_signal_11376, new_AGEMA_signal_11375, add_sub1_3_subc_rom_sbox_7_ANF_2_n13}), .b ({new_AGEMA_signal_8539, new_AGEMA_signal_8538, new_AGEMA_signal_8537, add_sub1_3_addc_out[1]}), .c ({new_AGEMA_signal_12817, new_AGEMA_signal_12816, new_AGEMA_signal_12815, add_sub1_3_subc_rom_sbox_7_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U6 ( .a ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, new_AGEMA_signal_10394, add_sub1_3_subc_rom_sbox_7_ANF_2_n18}), .b ({new_AGEMA_signal_10177, new_AGEMA_signal_10176, new_AGEMA_signal_10175, add_sub1_3_subc_rom_sbox_7_ANF_2_t3}), .c ({new_AGEMA_signal_11377, new_AGEMA_signal_11376, new_AGEMA_signal_11375, add_sub1_3_subc_rom_sbox_7_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_U5 ( .a ({new_AGEMA_signal_10180, new_AGEMA_signal_10179, new_AGEMA_signal_10178, add_sub1_3_subc_rom_sbox_7_ANF_2_t6}), .b ({new_AGEMA_signal_8533, new_AGEMA_signal_8532, new_AGEMA_signal_8531, add_sub1_3_addc_out[3]}), .c ({new_AGEMA_signal_10396, new_AGEMA_signal_10395, new_AGEMA_signal_10394, add_sub1_3_subc_rom_sbox_7_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_8542, new_AGEMA_signal_8541, new_AGEMA_signal_8540, add_sub1_3_addc_out[0]}), .b ({new_AGEMA_signal_9337, new_AGEMA_signal_9336, new_AGEMA_signal_9335, add_sub1_3_subc_rom_sbox_7_ANF_2_t0}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_10177, new_AGEMA_signal_10176, new_AGEMA_signal_10175, add_sub1_3_subc_rom_sbox_7_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_7_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_9334, new_AGEMA_signal_9333, new_AGEMA_signal_9332, add_sub1_3_subc_rom_sbox_7_ANF_2_t5}), .b ({new_AGEMA_signal_9346, new_AGEMA_signal_9345, new_AGEMA_signal_9344, add_sub1_3_subc_rom_sbox_7_ANF_2_t4}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_10180, new_AGEMA_signal_10179, new_AGEMA_signal_10178, add_sub1_3_subc_rom_sbox_7_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U14 ( .a ({new_AGEMA_signal_8545, new_AGEMA_signal_8544, new_AGEMA_signal_8543, add_sub1_3_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_7831, new_AGEMA_signal_7830, new_AGEMA_signal_7829, add_sub1_3_subc_rom_sbox_6_ANF_2_n19}), .c ({new_AGEMA_signal_9352, new_AGEMA_signal_9351, new_AGEMA_signal_9350, subc_out[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U13 ( .a ({new_AGEMA_signal_8122, new_AGEMA_signal_8121, new_AGEMA_signal_8120, add_sub1_3_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_8119, new_AGEMA_signal_8118, new_AGEMA_signal_8117, add_sub1_3_subc_rom_sbox_6_ANF_2_n17}), .c ({new_AGEMA_signal_8320, new_AGEMA_signal_8319, new_AGEMA_signal_8318, subc_out[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U9 ( .a ({new_AGEMA_signal_9355, new_AGEMA_signal_9354, new_AGEMA_signal_9353, add_sub1_3_subc_rom_sbox_6_ANF_2_n14}), .b ({new_AGEMA_signal_7363, new_AGEMA_signal_7362, new_AGEMA_signal_7361, add_sub1_3_subc_rom_sbox_6_ANF_2_t2}), .c ({new_AGEMA_signal_10183, new_AGEMA_signal_10182, new_AGEMA_signal_10181, subc_out[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U8 ( .a ({new_AGEMA_signal_8545, new_AGEMA_signal_8544, new_AGEMA_signal_8543, add_sub1_3_subc_rom_sbox_6_ANF_2_n20}), .b ({new_AGEMA_signal_7360, new_AGEMA_signal_7359, new_AGEMA_signal_7358, add_sub1_3_subc_rom_sbox_6_ANF_2_t1}), .c ({new_AGEMA_signal_9355, new_AGEMA_signal_9354, new_AGEMA_signal_9353, add_sub1_3_subc_rom_sbox_6_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U7 ( .a ({new_AGEMA_signal_8323, new_AGEMA_signal_8322, new_AGEMA_signal_8321, add_sub1_3_subc_rom_sbox_6_ANF_2_n13}), .b ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, new_AGEMA_signal_5963, addc_in[25]}), .c ({new_AGEMA_signal_8545, new_AGEMA_signal_8544, new_AGEMA_signal_8543, add_sub1_3_subc_rom_sbox_6_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U6 ( .a ({new_AGEMA_signal_8122, new_AGEMA_signal_8121, new_AGEMA_signal_8120, add_sub1_3_subc_rom_sbox_6_ANF_2_n18}), .b ({new_AGEMA_signal_7834, new_AGEMA_signal_7833, new_AGEMA_signal_7832, add_sub1_3_subc_rom_sbox_6_ANF_2_t3}), .c ({new_AGEMA_signal_8323, new_AGEMA_signal_8322, new_AGEMA_signal_8321, add_sub1_3_subc_rom_sbox_6_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_U5 ( .a ({new_AGEMA_signal_7837, new_AGEMA_signal_7836, new_AGEMA_signal_7835, add_sub1_3_subc_rom_sbox_6_ANF_2_t6}), .b ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, new_AGEMA_signal_5981, addc_in[27]}), .c ({new_AGEMA_signal_8122, new_AGEMA_signal_8121, new_AGEMA_signal_8120, add_sub1_3_subc_rom_sbox_6_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5956, new_AGEMA_signal_5955, new_AGEMA_signal_5954, addc_in[24]}), .b ({new_AGEMA_signal_7357, new_AGEMA_signal_7356, new_AGEMA_signal_7355, add_sub1_3_subc_rom_sbox_6_ANF_2_t0}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_7834, new_AGEMA_signal_7833, new_AGEMA_signal_7832, add_sub1_3_subc_rom_sbox_6_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_6_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7354, new_AGEMA_signal_7353, new_AGEMA_signal_7352, add_sub1_3_subc_rom_sbox_6_ANF_2_t5}), .b ({new_AGEMA_signal_7366, new_AGEMA_signal_7365, new_AGEMA_signal_7364, add_sub1_3_subc_rom_sbox_6_ANF_2_t4}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_7837, new_AGEMA_signal_7836, new_AGEMA_signal_7835, add_sub1_3_subc_rom_sbox_6_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U14 ( .a ({new_AGEMA_signal_8548, new_AGEMA_signal_8547, new_AGEMA_signal_8546, add_sub1_3_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_7846, new_AGEMA_signal_7845, new_AGEMA_signal_7844, add_sub1_3_subc_rom_sbox_5_ANF_2_n19}), .c ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, new_AGEMA_signal_9356, subc_out[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U13 ( .a ({new_AGEMA_signal_8131, new_AGEMA_signal_8130, new_AGEMA_signal_8129, add_sub1_3_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_8128, new_AGEMA_signal_8127, new_AGEMA_signal_8126, add_sub1_3_subc_rom_sbox_5_ANF_2_n17}), .c ({new_AGEMA_signal_8326, new_AGEMA_signal_8325, new_AGEMA_signal_8324, subc_out[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U9 ( .a ({new_AGEMA_signal_9361, new_AGEMA_signal_9360, new_AGEMA_signal_9359, add_sub1_3_subc_rom_sbox_5_ANF_2_n14}), .b ({new_AGEMA_signal_7384, new_AGEMA_signal_7383, new_AGEMA_signal_7382, add_sub1_3_subc_rom_sbox_5_ANF_2_t2}), .c ({new_AGEMA_signal_10186, new_AGEMA_signal_10185, new_AGEMA_signal_10184, subc_out[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U8 ( .a ({new_AGEMA_signal_8548, new_AGEMA_signal_8547, new_AGEMA_signal_8546, add_sub1_3_subc_rom_sbox_5_ANF_2_n20}), .b ({new_AGEMA_signal_7381, new_AGEMA_signal_7380, new_AGEMA_signal_7379, add_sub1_3_subc_rom_sbox_5_ANF_2_t1}), .c ({new_AGEMA_signal_9361, new_AGEMA_signal_9360, new_AGEMA_signal_9359, add_sub1_3_subc_rom_sbox_5_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U7 ( .a ({new_AGEMA_signal_8329, new_AGEMA_signal_8328, new_AGEMA_signal_8327, add_sub1_3_subc_rom_sbox_5_ANF_2_n13}), .b ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, new_AGEMA_signal_5927, addc_in[21]}), .c ({new_AGEMA_signal_8548, new_AGEMA_signal_8547, new_AGEMA_signal_8546, add_sub1_3_subc_rom_sbox_5_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U6 ( .a ({new_AGEMA_signal_8131, new_AGEMA_signal_8130, new_AGEMA_signal_8129, add_sub1_3_subc_rom_sbox_5_ANF_2_n18}), .b ({new_AGEMA_signal_7849, new_AGEMA_signal_7848, new_AGEMA_signal_7847, add_sub1_3_subc_rom_sbox_5_ANF_2_t3}), .c ({new_AGEMA_signal_8329, new_AGEMA_signal_8328, new_AGEMA_signal_8327, add_sub1_3_subc_rom_sbox_5_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_U5 ( .a ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, new_AGEMA_signal_7850, add_sub1_3_subc_rom_sbox_5_ANF_2_t6}), .b ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, new_AGEMA_signal_5945, addc_in[23]}), .c ({new_AGEMA_signal_8131, new_AGEMA_signal_8130, new_AGEMA_signal_8129, add_sub1_3_subc_rom_sbox_5_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5920, new_AGEMA_signal_5919, new_AGEMA_signal_5918, addc_in[20]}), .b ({new_AGEMA_signal_7378, new_AGEMA_signal_7377, new_AGEMA_signal_7376, add_sub1_3_subc_rom_sbox_5_ANF_2_t0}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_7849, new_AGEMA_signal_7848, new_AGEMA_signal_7847, add_sub1_3_subc_rom_sbox_5_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_5_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7375, new_AGEMA_signal_7374, new_AGEMA_signal_7373, add_sub1_3_subc_rom_sbox_5_ANF_2_t5}), .b ({new_AGEMA_signal_7387, new_AGEMA_signal_7386, new_AGEMA_signal_7385, add_sub1_3_subc_rom_sbox_5_ANF_2_t4}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_7852, new_AGEMA_signal_7851, new_AGEMA_signal_7850, add_sub1_3_subc_rom_sbox_5_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U14 ( .a ({new_AGEMA_signal_8551, new_AGEMA_signal_8550, new_AGEMA_signal_8549, add_sub1_3_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_7861, new_AGEMA_signal_7860, new_AGEMA_signal_7859, add_sub1_3_subc_rom_sbox_4_ANF_2_n19}), .c ({new_AGEMA_signal_9364, new_AGEMA_signal_9363, new_AGEMA_signal_9362, subc_out[19]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U13 ( .a ({new_AGEMA_signal_8140, new_AGEMA_signal_8139, new_AGEMA_signal_8138, add_sub1_3_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_8137, new_AGEMA_signal_8136, new_AGEMA_signal_8135, add_sub1_3_subc_rom_sbox_4_ANF_2_n17}), .c ({new_AGEMA_signal_8332, new_AGEMA_signal_8331, new_AGEMA_signal_8330, subc_out[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U9 ( .a ({new_AGEMA_signal_9367, new_AGEMA_signal_9366, new_AGEMA_signal_9365, add_sub1_3_subc_rom_sbox_4_ANF_2_n14}), .b ({new_AGEMA_signal_7405, new_AGEMA_signal_7404, new_AGEMA_signal_7403, add_sub1_3_subc_rom_sbox_4_ANF_2_t2}), .c ({new_AGEMA_signal_10189, new_AGEMA_signal_10188, new_AGEMA_signal_10187, subc_out[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U8 ( .a ({new_AGEMA_signal_8551, new_AGEMA_signal_8550, new_AGEMA_signal_8549, add_sub1_3_subc_rom_sbox_4_ANF_2_n20}), .b ({new_AGEMA_signal_7402, new_AGEMA_signal_7401, new_AGEMA_signal_7400, add_sub1_3_subc_rom_sbox_4_ANF_2_t1}), .c ({new_AGEMA_signal_9367, new_AGEMA_signal_9366, new_AGEMA_signal_9365, add_sub1_3_subc_rom_sbox_4_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U7 ( .a ({new_AGEMA_signal_8335, new_AGEMA_signal_8334, new_AGEMA_signal_8333, add_sub1_3_subc_rom_sbox_4_ANF_2_n13}), .b ({new_AGEMA_signal_5893, new_AGEMA_signal_5892, new_AGEMA_signal_5891, addc_in[17]}), .c ({new_AGEMA_signal_8551, new_AGEMA_signal_8550, new_AGEMA_signal_8549, add_sub1_3_subc_rom_sbox_4_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U6 ( .a ({new_AGEMA_signal_8140, new_AGEMA_signal_8139, new_AGEMA_signal_8138, add_sub1_3_subc_rom_sbox_4_ANF_2_n18}), .b ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, new_AGEMA_signal_7862, add_sub1_3_subc_rom_sbox_4_ANF_2_t3}), .c ({new_AGEMA_signal_8335, new_AGEMA_signal_8334, new_AGEMA_signal_8333, add_sub1_3_subc_rom_sbox_4_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_U5 ( .a ({new_AGEMA_signal_7867, new_AGEMA_signal_7866, new_AGEMA_signal_7865, add_sub1_3_subc_rom_sbox_4_ANF_2_t6}), .b ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, new_AGEMA_signal_5909, addc_in[19]}), .c ({new_AGEMA_signal_8140, new_AGEMA_signal_8139, new_AGEMA_signal_8138, add_sub1_3_subc_rom_sbox_4_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5884, new_AGEMA_signal_5883, new_AGEMA_signal_5882, addc_in[16]}), .b ({new_AGEMA_signal_7399, new_AGEMA_signal_7398, new_AGEMA_signal_7397, add_sub1_3_subc_rom_sbox_4_ANF_2_t0}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_7864, new_AGEMA_signal_7863, new_AGEMA_signal_7862, add_sub1_3_subc_rom_sbox_4_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_4_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7396, new_AGEMA_signal_7395, new_AGEMA_signal_7394, add_sub1_3_subc_rom_sbox_4_ANF_2_t5}), .b ({new_AGEMA_signal_7408, new_AGEMA_signal_7407, new_AGEMA_signal_7406, add_sub1_3_subc_rom_sbox_4_ANF_2_t4}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_7867, new_AGEMA_signal_7866, new_AGEMA_signal_7865, add_sub1_3_subc_rom_sbox_4_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U14 ( .a ({new_AGEMA_signal_8554, new_AGEMA_signal_8553, new_AGEMA_signal_8552, add_sub1_3_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_7876, new_AGEMA_signal_7875, new_AGEMA_signal_7874, add_sub1_3_subc_rom_sbox_3_ANF_2_n19}), .c ({new_AGEMA_signal_9370, new_AGEMA_signal_9369, new_AGEMA_signal_9368, subc_out[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U13 ( .a ({new_AGEMA_signal_8149, new_AGEMA_signal_8148, new_AGEMA_signal_8147, add_sub1_3_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_8146, new_AGEMA_signal_8145, new_AGEMA_signal_8144, add_sub1_3_subc_rom_sbox_3_ANF_2_n17}), .c ({new_AGEMA_signal_8338, new_AGEMA_signal_8337, new_AGEMA_signal_8336, subc_out[14]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U9 ( .a ({new_AGEMA_signal_9373, new_AGEMA_signal_9372, new_AGEMA_signal_9371, add_sub1_3_subc_rom_sbox_3_ANF_2_n14}), .b ({new_AGEMA_signal_7426, new_AGEMA_signal_7425, new_AGEMA_signal_7424, add_sub1_3_subc_rom_sbox_3_ANF_2_t2}), .c ({new_AGEMA_signal_10192, new_AGEMA_signal_10191, new_AGEMA_signal_10190, subc_out[13]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U8 ( .a ({new_AGEMA_signal_8554, new_AGEMA_signal_8553, new_AGEMA_signal_8552, add_sub1_3_subc_rom_sbox_3_ANF_2_n20}), .b ({new_AGEMA_signal_7423, new_AGEMA_signal_7422, new_AGEMA_signal_7421, add_sub1_3_subc_rom_sbox_3_ANF_2_t1}), .c ({new_AGEMA_signal_9373, new_AGEMA_signal_9372, new_AGEMA_signal_9371, add_sub1_3_subc_rom_sbox_3_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U7 ( .a ({new_AGEMA_signal_8341, new_AGEMA_signal_8340, new_AGEMA_signal_8339, add_sub1_3_subc_rom_sbox_3_ANF_2_n13}), .b ({new_AGEMA_signal_5857, new_AGEMA_signal_5856, new_AGEMA_signal_5855, addc_in[13]}), .c ({new_AGEMA_signal_8554, new_AGEMA_signal_8553, new_AGEMA_signal_8552, add_sub1_3_subc_rom_sbox_3_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U6 ( .a ({new_AGEMA_signal_8149, new_AGEMA_signal_8148, new_AGEMA_signal_8147, add_sub1_3_subc_rom_sbox_3_ANF_2_n18}), .b ({new_AGEMA_signal_7879, new_AGEMA_signal_7878, new_AGEMA_signal_7877, add_sub1_3_subc_rom_sbox_3_ANF_2_t3}), .c ({new_AGEMA_signal_8341, new_AGEMA_signal_8340, new_AGEMA_signal_8339, add_sub1_3_subc_rom_sbox_3_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_U5 ( .a ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, new_AGEMA_signal_7880, add_sub1_3_subc_rom_sbox_3_ANF_2_t6}), .b ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, new_AGEMA_signal_5873, addc_in[15]}), .c ({new_AGEMA_signal_8149, new_AGEMA_signal_8148, new_AGEMA_signal_8147, add_sub1_3_subc_rom_sbox_3_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5848, new_AGEMA_signal_5847, new_AGEMA_signal_5846, addc_in[12]}), .b ({new_AGEMA_signal_7420, new_AGEMA_signal_7419, new_AGEMA_signal_7418, add_sub1_3_subc_rom_sbox_3_ANF_2_t0}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_7879, new_AGEMA_signal_7878, new_AGEMA_signal_7877, add_sub1_3_subc_rom_sbox_3_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_3_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7417, new_AGEMA_signal_7416, new_AGEMA_signal_7415, add_sub1_3_subc_rom_sbox_3_ANF_2_t5}), .b ({new_AGEMA_signal_7429, new_AGEMA_signal_7428, new_AGEMA_signal_7427, add_sub1_3_subc_rom_sbox_3_ANF_2_t4}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_7882, new_AGEMA_signal_7881, new_AGEMA_signal_7880, add_sub1_3_subc_rom_sbox_3_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U14 ( .a ({new_AGEMA_signal_8557, new_AGEMA_signal_8556, new_AGEMA_signal_8555, add_sub1_3_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_7891, new_AGEMA_signal_7890, new_AGEMA_signal_7889, add_sub1_3_subc_rom_sbox_2_ANF_2_n19}), .c ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, new_AGEMA_signal_9374, subc_out[11]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U13 ( .a ({new_AGEMA_signal_8158, new_AGEMA_signal_8157, new_AGEMA_signal_8156, add_sub1_3_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_8155, new_AGEMA_signal_8154, new_AGEMA_signal_8153, add_sub1_3_subc_rom_sbox_2_ANF_2_n17}), .c ({new_AGEMA_signal_8344, new_AGEMA_signal_8343, new_AGEMA_signal_8342, subc_out[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U9 ( .a ({new_AGEMA_signal_9379, new_AGEMA_signal_9378, new_AGEMA_signal_9377, add_sub1_3_subc_rom_sbox_2_ANF_2_n14}), .b ({new_AGEMA_signal_7447, new_AGEMA_signal_7446, new_AGEMA_signal_7445, add_sub1_3_subc_rom_sbox_2_ANF_2_t2}), .c ({new_AGEMA_signal_10195, new_AGEMA_signal_10194, new_AGEMA_signal_10193, subc_out[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U8 ( .a ({new_AGEMA_signal_8557, new_AGEMA_signal_8556, new_AGEMA_signal_8555, add_sub1_3_subc_rom_sbox_2_ANF_2_n20}), .b ({new_AGEMA_signal_7444, new_AGEMA_signal_7443, new_AGEMA_signal_7442, add_sub1_3_subc_rom_sbox_2_ANF_2_t1}), .c ({new_AGEMA_signal_9379, new_AGEMA_signal_9378, new_AGEMA_signal_9377, add_sub1_3_subc_rom_sbox_2_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U7 ( .a ({new_AGEMA_signal_8347, new_AGEMA_signal_8346, new_AGEMA_signal_8345, add_sub1_3_subc_rom_sbox_2_ANF_2_n13}), .b ({new_AGEMA_signal_5821, new_AGEMA_signal_5820, new_AGEMA_signal_5819, addc_in[9]}), .c ({new_AGEMA_signal_8557, new_AGEMA_signal_8556, new_AGEMA_signal_8555, add_sub1_3_subc_rom_sbox_2_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U6 ( .a ({new_AGEMA_signal_8158, new_AGEMA_signal_8157, new_AGEMA_signal_8156, add_sub1_3_subc_rom_sbox_2_ANF_2_n18}), .b ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, new_AGEMA_signal_7892, add_sub1_3_subc_rom_sbox_2_ANF_2_t3}), .c ({new_AGEMA_signal_8347, new_AGEMA_signal_8346, new_AGEMA_signal_8345, add_sub1_3_subc_rom_sbox_2_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_U5 ( .a ({new_AGEMA_signal_7897, new_AGEMA_signal_7896, new_AGEMA_signal_7895, add_sub1_3_subc_rom_sbox_2_ANF_2_t6}), .b ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, new_AGEMA_signal_5837, addc_in[11]}), .c ({new_AGEMA_signal_8158, new_AGEMA_signal_8157, new_AGEMA_signal_8156, add_sub1_3_subc_rom_sbox_2_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5812, new_AGEMA_signal_5811, new_AGEMA_signal_5810, addc_in[8]}), .b ({new_AGEMA_signal_7441, new_AGEMA_signal_7440, new_AGEMA_signal_7439, add_sub1_3_subc_rom_sbox_2_ANF_2_t0}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_7894, new_AGEMA_signal_7893, new_AGEMA_signal_7892, add_sub1_3_subc_rom_sbox_2_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_2_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7438, new_AGEMA_signal_7437, new_AGEMA_signal_7436, add_sub1_3_subc_rom_sbox_2_ANF_2_t5}), .b ({new_AGEMA_signal_7450, new_AGEMA_signal_7449, new_AGEMA_signal_7448, add_sub1_3_subc_rom_sbox_2_ANF_2_t4}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_7897, new_AGEMA_signal_7896, new_AGEMA_signal_7895, add_sub1_3_subc_rom_sbox_2_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U14 ( .a ({new_AGEMA_signal_8560, new_AGEMA_signal_8559, new_AGEMA_signal_8558, add_sub1_3_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7906, new_AGEMA_signal_7905, new_AGEMA_signal_7904, add_sub1_3_subc_rom_sbox_1_ANF_2_n19}), .c ({new_AGEMA_signal_9382, new_AGEMA_signal_9381, new_AGEMA_signal_9380, subc_out[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U13 ( .a ({new_AGEMA_signal_8167, new_AGEMA_signal_8166, new_AGEMA_signal_8165, add_sub1_3_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_8164, new_AGEMA_signal_8163, new_AGEMA_signal_8162, add_sub1_3_subc_rom_sbox_1_ANF_2_n17}), .c ({new_AGEMA_signal_8350, new_AGEMA_signal_8349, new_AGEMA_signal_8348, subc_out[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U9 ( .a ({new_AGEMA_signal_9385, new_AGEMA_signal_9384, new_AGEMA_signal_9383, add_sub1_3_subc_rom_sbox_1_ANF_2_n14}), .b ({new_AGEMA_signal_7468, new_AGEMA_signal_7467, new_AGEMA_signal_7466, add_sub1_3_subc_rom_sbox_1_ANF_2_t2}), .c ({new_AGEMA_signal_10198, new_AGEMA_signal_10197, new_AGEMA_signal_10196, subc_out[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U8 ( .a ({new_AGEMA_signal_8560, new_AGEMA_signal_8559, new_AGEMA_signal_8558, add_sub1_3_subc_rom_sbox_1_ANF_2_n20}), .b ({new_AGEMA_signal_7465, new_AGEMA_signal_7464, new_AGEMA_signal_7463, add_sub1_3_subc_rom_sbox_1_ANF_2_t1}), .c ({new_AGEMA_signal_9385, new_AGEMA_signal_9384, new_AGEMA_signal_9383, add_sub1_3_subc_rom_sbox_1_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U7 ( .a ({new_AGEMA_signal_8353, new_AGEMA_signal_8352, new_AGEMA_signal_8351, add_sub1_3_subc_rom_sbox_1_ANF_2_n13}), .b ({new_AGEMA_signal_5785, new_AGEMA_signal_5784, new_AGEMA_signal_5783, addc_in[5]}), .c ({new_AGEMA_signal_8560, new_AGEMA_signal_8559, new_AGEMA_signal_8558, add_sub1_3_subc_rom_sbox_1_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U6 ( .a ({new_AGEMA_signal_8167, new_AGEMA_signal_8166, new_AGEMA_signal_8165, add_sub1_3_subc_rom_sbox_1_ANF_2_n18}), .b ({new_AGEMA_signal_7909, new_AGEMA_signal_7908, new_AGEMA_signal_7907, add_sub1_3_subc_rom_sbox_1_ANF_2_t3}), .c ({new_AGEMA_signal_8353, new_AGEMA_signal_8352, new_AGEMA_signal_8351, add_sub1_3_subc_rom_sbox_1_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_U5 ( .a ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, new_AGEMA_signal_7910, add_sub1_3_subc_rom_sbox_1_ANF_2_t6}), .b ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, new_AGEMA_signal_5801, addc_in[7]}), .c ({new_AGEMA_signal_8167, new_AGEMA_signal_8166, new_AGEMA_signal_8165, add_sub1_3_subc_rom_sbox_1_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, new_AGEMA_signal_5774, addc_in[4]}), .b ({new_AGEMA_signal_7462, new_AGEMA_signal_7461, new_AGEMA_signal_7460, add_sub1_3_subc_rom_sbox_1_ANF_2_t0}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_7909, new_AGEMA_signal_7908, new_AGEMA_signal_7907, add_sub1_3_subc_rom_sbox_1_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_1_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7459, new_AGEMA_signal_7458, new_AGEMA_signal_7457, add_sub1_3_subc_rom_sbox_1_ANF_2_t5}), .b ({new_AGEMA_signal_7471, new_AGEMA_signal_7470, new_AGEMA_signal_7469, add_sub1_3_subc_rom_sbox_1_ANF_2_t4}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_7912, new_AGEMA_signal_7911, new_AGEMA_signal_7910, add_sub1_3_subc_rom_sbox_1_ANF_2_t6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U14 ( .a ({new_AGEMA_signal_8563, new_AGEMA_signal_8562, new_AGEMA_signal_8561, add_sub1_3_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7921, new_AGEMA_signal_7920, new_AGEMA_signal_7919, add_sub1_3_subc_rom_sbox_0_ANF_2_n19}), .c ({new_AGEMA_signal_9388, new_AGEMA_signal_9387, new_AGEMA_signal_9386, subc_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U13 ( .a ({new_AGEMA_signal_8176, new_AGEMA_signal_8175, new_AGEMA_signal_8174, add_sub1_3_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_8173, new_AGEMA_signal_8172, new_AGEMA_signal_8171, add_sub1_3_subc_rom_sbox_0_ANF_2_n17}), .c ({new_AGEMA_signal_8356, new_AGEMA_signal_8355, new_AGEMA_signal_8354, subc_out[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U9 ( .a ({new_AGEMA_signal_9391, new_AGEMA_signal_9390, new_AGEMA_signal_9389, add_sub1_3_subc_rom_sbox_0_ANF_2_n14}), .b ({new_AGEMA_signal_7489, new_AGEMA_signal_7488, new_AGEMA_signal_7487, add_sub1_3_subc_rom_sbox_0_ANF_2_t2}), .c ({new_AGEMA_signal_10201, new_AGEMA_signal_10200, new_AGEMA_signal_10199, subc_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U8 ( .a ({new_AGEMA_signal_8563, new_AGEMA_signal_8562, new_AGEMA_signal_8561, add_sub1_3_subc_rom_sbox_0_ANF_2_n20}), .b ({new_AGEMA_signal_7486, new_AGEMA_signal_7485, new_AGEMA_signal_7484, add_sub1_3_subc_rom_sbox_0_ANF_2_t1}), .c ({new_AGEMA_signal_9391, new_AGEMA_signal_9390, new_AGEMA_signal_9389, add_sub1_3_subc_rom_sbox_0_ANF_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U7 ( .a ({new_AGEMA_signal_8359, new_AGEMA_signal_8358, new_AGEMA_signal_8357, add_sub1_3_subc_rom_sbox_0_ANF_2_n13}), .b ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, new_AGEMA_signal_5747, addc_in[1]}), .c ({new_AGEMA_signal_8563, new_AGEMA_signal_8562, new_AGEMA_signal_8561, add_sub1_3_subc_rom_sbox_0_ANF_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U6 ( .a ({new_AGEMA_signal_8176, new_AGEMA_signal_8175, new_AGEMA_signal_8174, add_sub1_3_subc_rom_sbox_0_ANF_2_n18}), .b ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, new_AGEMA_signal_7922, add_sub1_3_subc_rom_sbox_0_ANF_2_t3}), .c ({new_AGEMA_signal_8359, new_AGEMA_signal_8358, new_AGEMA_signal_8357, add_sub1_3_subc_rom_sbox_0_ANF_2_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_U5 ( .a ({new_AGEMA_signal_7927, new_AGEMA_signal_7926, new_AGEMA_signal_7925, add_sub1_3_subc_rom_sbox_0_ANF_2_t6}), .b ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, new_AGEMA_signal_5765, addc_in[3]}), .c ({new_AGEMA_signal_8176, new_AGEMA_signal_8175, new_AGEMA_signal_8174, add_sub1_3_subc_rom_sbox_0_ANF_2_n18}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t3_AND_U1 ( .a ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, new_AGEMA_signal_5738, addc_in[0]}), .b ({new_AGEMA_signal_7483, new_AGEMA_signal_7482, new_AGEMA_signal_7481, add_sub1_3_subc_rom_sbox_0_ANF_2_t0}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_7924, new_AGEMA_signal_7923, new_AGEMA_signal_7922, add_sub1_3_subc_rom_sbox_0_ANF_2_t3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) add_sub1_3_subc_rom_sbox_0_ANF_2_t6_AND_U1 ( .a ({new_AGEMA_signal_7480, new_AGEMA_signal_7479, new_AGEMA_signal_7478, add_sub1_3_subc_rom_sbox_0_ANF_2_t5}), .b ({new_AGEMA_signal_7492, new_AGEMA_signal_7491, new_AGEMA_signal_7490, add_sub1_3_subc_rom_sbox_0_ANF_2_t4}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_7927, new_AGEMA_signal_7926, new_AGEMA_signal_7925, add_sub1_3_subc_rom_sbox_0_ANF_2_t6}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10093, new_AGEMA_signal_10092, new_AGEMA_signal_10091, subc_out[97]}), .a ({new_AGEMA_signal_10081, new_AGEMA_signal_10080, new_AGEMA_signal_10079, subc_out[113]}), .c ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8221, new_AGEMA_signal_8220, new_AGEMA_signal_8219, subc_out[98]}), .a ({new_AGEMA_signal_8197, new_AGEMA_signal_8196, new_AGEMA_signal_8195, subc_out[114]}), .c ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9199, new_AGEMA_signal_9198, new_AGEMA_signal_9197, subc_out[99]}), .a ({new_AGEMA_signal_9175, new_AGEMA_signal_9174, new_AGEMA_signal_9173, subc_out[115]}), .c ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, new_AGEMA_signal_10088, subc_out[101]}), .a ({new_AGEMA_signal_10078, new_AGEMA_signal_10077, new_AGEMA_signal_10076, subc_out[117]}), .c ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8215, new_AGEMA_signal_8214, new_AGEMA_signal_8213, subc_out[102]}), .a ({new_AGEMA_signal_8191, new_AGEMA_signal_8190, new_AGEMA_signal_8189, subc_out[118]}), .c ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9193, new_AGEMA_signal_9192, new_AGEMA_signal_9191, subc_out[103]}), .a ({new_AGEMA_signal_9169, new_AGEMA_signal_9168, new_AGEMA_signal_9167, subc_out[119]}), .c ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10087, new_AGEMA_signal_10086, new_AGEMA_signal_10085, subc_out[105]}), .a ({new_AGEMA_signal_10075, new_AGEMA_signal_10074, new_AGEMA_signal_10073, subc_out[121]}), .c ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8209, new_AGEMA_signal_8208, new_AGEMA_signal_8207, subc_out[106]}), .a ({new_AGEMA_signal_8185, new_AGEMA_signal_8184, new_AGEMA_signal_8183, subc_out[122]}), .c ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9187, new_AGEMA_signal_9186, new_AGEMA_signal_9185, subc_out[107]}), .a ({new_AGEMA_signal_9163, new_AGEMA_signal_9162, new_AGEMA_signal_9161, subc_out[123]}), .c ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10084, new_AGEMA_signal_10083, new_AGEMA_signal_10082, subc_out[109]}), .a ({new_AGEMA_signal_15682, new_AGEMA_signal_15681, new_AGEMA_signal_15680, subc_out[125]}), .c ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8203, new_AGEMA_signal_8202, new_AGEMA_signal_8201, subc_out[110]}), .a ({new_AGEMA_signal_11356, new_AGEMA_signal_11355, new_AGEMA_signal_11354, subc_out[126]}), .c ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9181, new_AGEMA_signal_9180, new_AGEMA_signal_9179, subc_out[111]}), .a ({new_AGEMA_signal_14254, new_AGEMA_signal_14253, new_AGEMA_signal_14252, subc_out[127]}), .c ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10081, new_AGEMA_signal_10080, new_AGEMA_signal_10079, subc_out[113]}), .a ({new_AGEMA_signal_10093, new_AGEMA_signal_10092, new_AGEMA_signal_10091, subc_out[97]}), .c ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8197, new_AGEMA_signal_8196, new_AGEMA_signal_8195, subc_out[114]}), .a ({new_AGEMA_signal_8221, new_AGEMA_signal_8220, new_AGEMA_signal_8219, subc_out[98]}), .c ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9175, new_AGEMA_signal_9174, new_AGEMA_signal_9173, subc_out[115]}), .a ({new_AGEMA_signal_9199, new_AGEMA_signal_9198, new_AGEMA_signal_9197, subc_out[99]}), .c ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10078, new_AGEMA_signal_10077, new_AGEMA_signal_10076, subc_out[117]}), .a ({new_AGEMA_signal_10090, new_AGEMA_signal_10089, new_AGEMA_signal_10088, subc_out[101]}), .c ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8191, new_AGEMA_signal_8190, new_AGEMA_signal_8189, subc_out[118]}), .a ({new_AGEMA_signal_8215, new_AGEMA_signal_8214, new_AGEMA_signal_8213, subc_out[102]}), .c ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9169, new_AGEMA_signal_9168, new_AGEMA_signal_9167, subc_out[119]}), .a ({new_AGEMA_signal_9193, new_AGEMA_signal_9192, new_AGEMA_signal_9191, subc_out[103]}), .c ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10075, new_AGEMA_signal_10074, new_AGEMA_signal_10073, subc_out[121]}), .a ({new_AGEMA_signal_10087, new_AGEMA_signal_10086, new_AGEMA_signal_10085, subc_out[105]}), .c ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8185, new_AGEMA_signal_8184, new_AGEMA_signal_8183, subc_out[122]}), .a ({new_AGEMA_signal_8209, new_AGEMA_signal_8208, new_AGEMA_signal_8207, subc_out[106]}), .c ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9163, new_AGEMA_signal_9162, new_AGEMA_signal_9161, subc_out[123]}), .a ({new_AGEMA_signal_9187, new_AGEMA_signal_9186, new_AGEMA_signal_9185, subc_out[107]}), .c ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15682, new_AGEMA_signal_15681, new_AGEMA_signal_15680, subc_out[125]}), .a ({new_AGEMA_signal_10084, new_AGEMA_signal_10083, new_AGEMA_signal_10082, subc_out[109]}), .c ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11356, new_AGEMA_signal_11355, new_AGEMA_signal_11354, subc_out[126]}), .a ({new_AGEMA_signal_8203, new_AGEMA_signal_8202, new_AGEMA_signal_8201, subc_out[110]}), .c ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_0_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14254, new_AGEMA_signal_14253, new_AGEMA_signal_14252, subc_out[127]}), .a ({new_AGEMA_signal_9181, new_AGEMA_signal_9180, new_AGEMA_signal_9179, subc_out[111]}), .c ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15685, new_AGEMA_signal_15684, new_AGEMA_signal_15683, subc_out[93]}), .a ({new_AGEMA_signal_10120, new_AGEMA_signal_10119, new_AGEMA_signal_10118, subc_out[77]}), .c ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11362, new_AGEMA_signal_11361, new_AGEMA_signal_11360, subc_out[94]}), .a ({new_AGEMA_signal_8248, new_AGEMA_signal_8247, new_AGEMA_signal_8246, subc_out[78]}), .c ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14260, new_AGEMA_signal_14259, new_AGEMA_signal_14258, subc_out[95]}), .a ({new_AGEMA_signal_9244, new_AGEMA_signal_9243, new_AGEMA_signal_9242, subc_out[79]}), .c ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10129, new_AGEMA_signal_10128, new_AGEMA_signal_10127, subc_out[65]}), .a ({new_AGEMA_signal_10117, new_AGEMA_signal_10116, new_AGEMA_signal_10115, subc_out[81]}), .c ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8266, new_AGEMA_signal_8265, new_AGEMA_signal_8264, subc_out[66]}), .a ({new_AGEMA_signal_8242, new_AGEMA_signal_8241, new_AGEMA_signal_8240, subc_out[82]}), .c ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9262, new_AGEMA_signal_9261, new_AGEMA_signal_9260, subc_out[67]}), .a ({new_AGEMA_signal_9238, new_AGEMA_signal_9237, new_AGEMA_signal_9236, subc_out[83]}), .c ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10126, new_AGEMA_signal_10125, new_AGEMA_signal_10124, subc_out[69]}), .a ({new_AGEMA_signal_10114, new_AGEMA_signal_10113, new_AGEMA_signal_10112, subc_out[85]}), .c ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8260, new_AGEMA_signal_8259, new_AGEMA_signal_8258, subc_out[70]}), .a ({new_AGEMA_signal_8236, new_AGEMA_signal_8235, new_AGEMA_signal_8234, subc_out[86]}), .c ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9256, new_AGEMA_signal_9255, new_AGEMA_signal_9254, subc_out[71]}), .a ({new_AGEMA_signal_9232, new_AGEMA_signal_9231, new_AGEMA_signal_9230, subc_out[87]}), .c ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10123, new_AGEMA_signal_10122, new_AGEMA_signal_10121, subc_out[73]}), .a ({new_AGEMA_signal_10111, new_AGEMA_signal_10110, new_AGEMA_signal_10109, subc_out[89]}), .c ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8254, new_AGEMA_signal_8253, new_AGEMA_signal_8252, subc_out[74]}), .a ({new_AGEMA_signal_8230, new_AGEMA_signal_8229, new_AGEMA_signal_8228, subc_out[90]}), .c ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9250, new_AGEMA_signal_9249, new_AGEMA_signal_9248, subc_out[75]}), .a ({new_AGEMA_signal_9226, new_AGEMA_signal_9225, new_AGEMA_signal_9224, subc_out[91]}), .c ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10120, new_AGEMA_signal_10119, new_AGEMA_signal_10118, subc_out[77]}), .a ({new_AGEMA_signal_15685, new_AGEMA_signal_15684, new_AGEMA_signal_15683, subc_out[93]}), .c ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8248, new_AGEMA_signal_8247, new_AGEMA_signal_8246, subc_out[78]}), .a ({new_AGEMA_signal_11362, new_AGEMA_signal_11361, new_AGEMA_signal_11360, subc_out[94]}), .c ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9244, new_AGEMA_signal_9243, new_AGEMA_signal_9242, subc_out[79]}), .a ({new_AGEMA_signal_14260, new_AGEMA_signal_14259, new_AGEMA_signal_14258, subc_out[95]}), .c ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10117, new_AGEMA_signal_10116, new_AGEMA_signal_10115, subc_out[81]}), .a ({new_AGEMA_signal_10129, new_AGEMA_signal_10128, new_AGEMA_signal_10127, subc_out[65]}), .c ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8242, new_AGEMA_signal_8241, new_AGEMA_signal_8240, subc_out[82]}), .a ({new_AGEMA_signal_8266, new_AGEMA_signal_8265, new_AGEMA_signal_8264, subc_out[66]}), .c ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9238, new_AGEMA_signal_9237, new_AGEMA_signal_9236, subc_out[83]}), .a ({new_AGEMA_signal_9262, new_AGEMA_signal_9261, new_AGEMA_signal_9260, subc_out[67]}), .c ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10114, new_AGEMA_signal_10113, new_AGEMA_signal_10112, subc_out[85]}), .a ({new_AGEMA_signal_10126, new_AGEMA_signal_10125, new_AGEMA_signal_10124, subc_out[69]}), .c ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8236, new_AGEMA_signal_8235, new_AGEMA_signal_8234, subc_out[86]}), .a ({new_AGEMA_signal_8260, new_AGEMA_signal_8259, new_AGEMA_signal_8258, subc_out[70]}), .c ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9232, new_AGEMA_signal_9231, new_AGEMA_signal_9230, subc_out[87]}), .a ({new_AGEMA_signal_9256, new_AGEMA_signal_9255, new_AGEMA_signal_9254, subc_out[71]}), .c ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10111, new_AGEMA_signal_10110, new_AGEMA_signal_10109, subc_out[89]}), .a ({new_AGEMA_signal_10123, new_AGEMA_signal_10122, new_AGEMA_signal_10121, subc_out[73]}), .c ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8230, new_AGEMA_signal_8229, new_AGEMA_signal_8228, subc_out[90]}), .a ({new_AGEMA_signal_8254, new_AGEMA_signal_8253, new_AGEMA_signal_8252, subc_out[74]}), .c ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_1_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9226, new_AGEMA_signal_9225, new_AGEMA_signal_9224, subc_out[91]}), .a ({new_AGEMA_signal_9250, new_AGEMA_signal_9249, new_AGEMA_signal_9248, subc_out[75]}), .c ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10147, new_AGEMA_signal_10146, new_AGEMA_signal_10145, subc_out[57]}), .a ({new_AGEMA_signal_10159, new_AGEMA_signal_10158, new_AGEMA_signal_10157, subc_out[41]}), .c ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8275, new_AGEMA_signal_8274, new_AGEMA_signal_8273, subc_out[58]}), .a ({new_AGEMA_signal_8299, new_AGEMA_signal_8298, new_AGEMA_signal_8297, subc_out[42]}), .c ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9289, new_AGEMA_signal_9288, new_AGEMA_signal_9287, subc_out[59]}), .a ({new_AGEMA_signal_9313, new_AGEMA_signal_9312, new_AGEMA_signal_9311, subc_out[43]}), .c ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15688, new_AGEMA_signal_15687, new_AGEMA_signal_15686, subc_out[61]}), .a ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, new_AGEMA_signal_10154, subc_out[45]}), .c ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11368, new_AGEMA_signal_11367, new_AGEMA_signal_11366, subc_out[62]}), .a ({new_AGEMA_signal_8293, new_AGEMA_signal_8292, new_AGEMA_signal_8291, subc_out[46]}), .c ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14266, new_AGEMA_signal_14265, new_AGEMA_signal_14264, subc_out[63]}), .a ({new_AGEMA_signal_9307, new_AGEMA_signal_9306, new_AGEMA_signal_9305, subc_out[47]}), .c ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10165, new_AGEMA_signal_10164, new_AGEMA_signal_10163, subc_out[33]}), .a ({new_AGEMA_signal_10153, new_AGEMA_signal_10152, new_AGEMA_signal_10151, subc_out[49]}), .c ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8311, new_AGEMA_signal_8310, new_AGEMA_signal_8309, subc_out[34]}), .a ({new_AGEMA_signal_8287, new_AGEMA_signal_8286, new_AGEMA_signal_8285, subc_out[50]}), .c ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9325, new_AGEMA_signal_9324, new_AGEMA_signal_9323, subc_out[35]}), .a ({new_AGEMA_signal_9301, new_AGEMA_signal_9300, new_AGEMA_signal_9299, subc_out[51]}), .c ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10162, new_AGEMA_signal_10161, new_AGEMA_signal_10160, subc_out[37]}), .a ({new_AGEMA_signal_10150, new_AGEMA_signal_10149, new_AGEMA_signal_10148, subc_out[53]}), .c ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8305, new_AGEMA_signal_8304, new_AGEMA_signal_8303, subc_out[38]}), .a ({new_AGEMA_signal_8281, new_AGEMA_signal_8280, new_AGEMA_signal_8279, subc_out[54]}), .c ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9319, new_AGEMA_signal_9318, new_AGEMA_signal_9317, subc_out[39]}), .a ({new_AGEMA_signal_9295, new_AGEMA_signal_9294, new_AGEMA_signal_9293, subc_out[55]}), .c ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10159, new_AGEMA_signal_10158, new_AGEMA_signal_10157, subc_out[41]}), .a ({new_AGEMA_signal_10147, new_AGEMA_signal_10146, new_AGEMA_signal_10145, subc_out[57]}), .c ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8299, new_AGEMA_signal_8298, new_AGEMA_signal_8297, subc_out[42]}), .a ({new_AGEMA_signal_8275, new_AGEMA_signal_8274, new_AGEMA_signal_8273, subc_out[58]}), .c ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9313, new_AGEMA_signal_9312, new_AGEMA_signal_9311, subc_out[43]}), .a ({new_AGEMA_signal_9289, new_AGEMA_signal_9288, new_AGEMA_signal_9287, subc_out[59]}), .c ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10156, new_AGEMA_signal_10155, new_AGEMA_signal_10154, subc_out[45]}), .a ({new_AGEMA_signal_15688, new_AGEMA_signal_15687, new_AGEMA_signal_15686, subc_out[61]}), .c ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8293, new_AGEMA_signal_8292, new_AGEMA_signal_8291, subc_out[46]}), .a ({new_AGEMA_signal_11368, new_AGEMA_signal_11367, new_AGEMA_signal_11366, subc_out[62]}), .c ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9307, new_AGEMA_signal_9306, new_AGEMA_signal_9305, subc_out[47]}), .a ({new_AGEMA_signal_14266, new_AGEMA_signal_14265, new_AGEMA_signal_14264, subc_out[63]}), .c ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10153, new_AGEMA_signal_10152, new_AGEMA_signal_10151, subc_out[49]}), .a ({new_AGEMA_signal_10165, new_AGEMA_signal_10164, new_AGEMA_signal_10163, subc_out[33]}), .c ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8287, new_AGEMA_signal_8286, new_AGEMA_signal_8285, subc_out[50]}), .a ({new_AGEMA_signal_8311, new_AGEMA_signal_8310, new_AGEMA_signal_8309, subc_out[34]}), .c ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9301, new_AGEMA_signal_9300, new_AGEMA_signal_9299, subc_out[51]}), .a ({new_AGEMA_signal_9325, new_AGEMA_signal_9324, new_AGEMA_signal_9323, subc_out[35]}), .c ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10150, new_AGEMA_signal_10149, new_AGEMA_signal_10148, subc_out[53]}), .a ({new_AGEMA_signal_10162, new_AGEMA_signal_10161, new_AGEMA_signal_10160, subc_out[37]}), .c ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8281, new_AGEMA_signal_8280, new_AGEMA_signal_8279, subc_out[54]}), .a ({new_AGEMA_signal_8305, new_AGEMA_signal_8304, new_AGEMA_signal_8303, subc_out[38]}), .c ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_2_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9295, new_AGEMA_signal_9294, new_AGEMA_signal_9293, subc_out[55]}), .a ({new_AGEMA_signal_9319, new_AGEMA_signal_9318, new_AGEMA_signal_9317, subc_out[39]}), .c ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10186, new_AGEMA_signal_10185, new_AGEMA_signal_10184, subc_out[21]}), .a ({new_AGEMA_signal_10198, new_AGEMA_signal_10197, new_AGEMA_signal_10196, subc_out[5]}), .c ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8326, new_AGEMA_signal_8325, new_AGEMA_signal_8324, subc_out[22]}), .a ({new_AGEMA_signal_8350, new_AGEMA_signal_8349, new_AGEMA_signal_8348, subc_out[6]}), .c ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, new_AGEMA_signal_9356, subc_out[23]}), .a ({new_AGEMA_signal_9382, new_AGEMA_signal_9381, new_AGEMA_signal_9380, subc_out[7]}), .c ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10183, new_AGEMA_signal_10182, new_AGEMA_signal_10181, subc_out[25]}), .a ({new_AGEMA_signal_10195, new_AGEMA_signal_10194, new_AGEMA_signal_10193, subc_out[9]}), .c ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8320, new_AGEMA_signal_8319, new_AGEMA_signal_8318, subc_out[26]}), .a ({new_AGEMA_signal_8344, new_AGEMA_signal_8343, new_AGEMA_signal_8342, subc_out[10]}), .c ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9352, new_AGEMA_signal_9351, new_AGEMA_signal_9350, subc_out[27]}), .a ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, new_AGEMA_signal_9374, subc_out[11]}), .c ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15691, new_AGEMA_signal_15690, new_AGEMA_signal_15689, subc_out[29]}), .a ({new_AGEMA_signal_10192, new_AGEMA_signal_10191, new_AGEMA_signal_10190, subc_out[13]}), .c ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_11374, new_AGEMA_signal_11373, new_AGEMA_signal_11372, subc_out[30]}), .a ({new_AGEMA_signal_8338, new_AGEMA_signal_8337, new_AGEMA_signal_8336, subc_out[14]}), .c ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_14272, new_AGEMA_signal_14271, new_AGEMA_signal_14270, subc_out[31]}), .a ({new_AGEMA_signal_9370, new_AGEMA_signal_9369, new_AGEMA_signal_9368, subc_out[15]}), .c ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10201, new_AGEMA_signal_10200, new_AGEMA_signal_10199, subc_out[1]}), .a ({new_AGEMA_signal_10189, new_AGEMA_signal_10188, new_AGEMA_signal_10187, subc_out[17]}), .c ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8356, new_AGEMA_signal_8355, new_AGEMA_signal_8354, subc_out[2]}), .a ({new_AGEMA_signal_8332, new_AGEMA_signal_8331, new_AGEMA_signal_8330, subc_out[18]}), .c ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9388, new_AGEMA_signal_9387, new_AGEMA_signal_9386, subc_out[3]}), .a ({new_AGEMA_signal_9364, new_AGEMA_signal_9363, new_AGEMA_signal_9362, subc_out[19]}), .c ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10198, new_AGEMA_signal_10197, new_AGEMA_signal_10196, subc_out[5]}), .a ({new_AGEMA_signal_10186, new_AGEMA_signal_10185, new_AGEMA_signal_10184, subc_out[21]}), .c ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8350, new_AGEMA_signal_8349, new_AGEMA_signal_8348, subc_out[6]}), .a ({new_AGEMA_signal_8326, new_AGEMA_signal_8325, new_AGEMA_signal_8324, subc_out[22]}), .c ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9382, new_AGEMA_signal_9381, new_AGEMA_signal_9380, subc_out[7]}), .a ({new_AGEMA_signal_9358, new_AGEMA_signal_9357, new_AGEMA_signal_9356, subc_out[23]}), .c ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10195, new_AGEMA_signal_10194, new_AGEMA_signal_10193, subc_out[9]}), .a ({new_AGEMA_signal_10183, new_AGEMA_signal_10182, new_AGEMA_signal_10181, subc_out[25]}), .c ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8344, new_AGEMA_signal_8343, new_AGEMA_signal_8342, subc_out[10]}), .a ({new_AGEMA_signal_8320, new_AGEMA_signal_8319, new_AGEMA_signal_8318, subc_out[26]}), .c ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9376, new_AGEMA_signal_9375, new_AGEMA_signal_9374, subc_out[11]}), .a ({new_AGEMA_signal_9352, new_AGEMA_signal_9351, new_AGEMA_signal_9350, subc_out[27]}), .c ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10192, new_AGEMA_signal_10191, new_AGEMA_signal_10190, subc_out[13]}), .a ({new_AGEMA_signal_15691, new_AGEMA_signal_15690, new_AGEMA_signal_15689, subc_out[29]}), .c ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8338, new_AGEMA_signal_8337, new_AGEMA_signal_8336, subc_out[14]}), .a ({new_AGEMA_signal_11374, new_AGEMA_signal_11373, new_AGEMA_signal_11372, subc_out[30]}), .c ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9370, new_AGEMA_signal_9369, new_AGEMA_signal_9368, subc_out[15]}), .a ({new_AGEMA_signal_14272, new_AGEMA_signal_14271, new_AGEMA_signal_14270, subc_out[31]}), .c ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_10189, new_AGEMA_signal_10188, new_AGEMA_signal_10187, subc_out[17]}), .a ({new_AGEMA_signal_10201, new_AGEMA_signal_10200, new_AGEMA_signal_10199, subc_out[1]}), .c ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_8332, new_AGEMA_signal_8331, new_AGEMA_signal_8330, subc_out[18]}), .a ({new_AGEMA_signal_8356, new_AGEMA_signal_8355, new_AGEMA_signal_8354, subc_out[2]}), .c ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) shiftr1_3_MUX_inst_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_9364, new_AGEMA_signal_9363, new_AGEMA_signal_9362, subc_out[19]}), .a ({new_AGEMA_signal_9388, new_AGEMA_signal_9387, new_AGEMA_signal_9386, subc_out[3]}), .c ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U44 ( .a ({new_AGEMA_signal_10513, new_AGEMA_signal_10512, new_AGEMA_signal_10511, mcs1_mcs_mat1_0_mcs_out[90]}), .b ({new_AGEMA_signal_17425, new_AGEMA_signal_17424, new_AGEMA_signal_17423, mcs1_mcs_mat1_0_mcs_out[94]}), .c ({new_AGEMA_signal_18127, new_AGEMA_signal_18126, new_AGEMA_signal_18125, mcs1_mcs_mat1_0_n93}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .c ({new_AGEMA_signal_16678, new_AGEMA_signal_16677, new_AGEMA_signal_16676, mcs1_mcs_mat1_0_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .b ({new_AGEMA_signal_8638, new_AGEMA_signal_8637, new_AGEMA_signal_8636, mcs1_mcs_mat1_0_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_9394, new_AGEMA_signal_9393, new_AGEMA_signal_9392, mcs1_mcs_mat1_0_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_8638, new_AGEMA_signal_8637, new_AGEMA_signal_8636, mcs1_mcs_mat1_0_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_10480, new_AGEMA_signal_10479, new_AGEMA_signal_10478, mcs1_mcs_mat1_0_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_11410, new_AGEMA_signal_11409, new_AGEMA_signal_11408, mcs1_mcs_mat1_0_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_8641, new_AGEMA_signal_8640, new_AGEMA_signal_8639, mcs1_mcs_mat1_0_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_10480, new_AGEMA_signal_10479, new_AGEMA_signal_10478, mcs1_mcs_mat1_0_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_8641, new_AGEMA_signal_8640, new_AGEMA_signal_8639, mcs1_mcs_mat1_0_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_8644, new_AGEMA_signal_8643, new_AGEMA_signal_8642, mcs1_mcs_mat1_0_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_11422, new_AGEMA_signal_11421, new_AGEMA_signal_11420, mcs1_mcs_mat1_0_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_12856, new_AGEMA_signal_12855, new_AGEMA_signal_12854, mcs1_mcs_mat1_0_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_9403, new_AGEMA_signal_9402, new_AGEMA_signal_9401, mcs1_mcs_mat1_0_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_10489, new_AGEMA_signal_10488, new_AGEMA_signal_10487, mcs1_mcs_mat1_0_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .c ({new_AGEMA_signal_9403, new_AGEMA_signal_9402, new_AGEMA_signal_9401, mcs1_mcs_mat1_0_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .b ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_11422, new_AGEMA_signal_11421, new_AGEMA_signal_11420, mcs1_mcs_mat1_0_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_8644, new_AGEMA_signal_8643, new_AGEMA_signal_8642, mcs1_mcs_mat1_0_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_17416, new_AGEMA_signal_17415, new_AGEMA_signal_17414, mcs1_mcs_mat1_0_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_18142, new_AGEMA_signal_18141, new_AGEMA_signal_18140, mcs1_mcs_mat1_0_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_12865, new_AGEMA_signal_12864, new_AGEMA_signal_12863, mcs1_mcs_mat1_0_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_17416, new_AGEMA_signal_17415, new_AGEMA_signal_17414, mcs1_mcs_mat1_0_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_12865, new_AGEMA_signal_12864, new_AGEMA_signal_12863, mcs1_mcs_mat1_0_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_8647, new_AGEMA_signal_8646, new_AGEMA_signal_8645, mcs1_mcs_mat1_0_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({new_AGEMA_signal_10501, new_AGEMA_signal_10500, new_AGEMA_signal_10499, mcs1_mcs_mat1_0_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_11434, new_AGEMA_signal_11433, new_AGEMA_signal_11432, mcs1_mcs_mat1_0_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_8650, new_AGEMA_signal_8649, new_AGEMA_signal_8648, mcs1_mcs_mat1_0_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_10501, new_AGEMA_signal_10500, new_AGEMA_signal_10499, mcs1_mcs_mat1_0_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .b ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .c ({new_AGEMA_signal_11437, new_AGEMA_signal_11436, new_AGEMA_signal_11435, mcs1_mcs_mat1_0_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_8650, new_AGEMA_signal_8649, new_AGEMA_signal_8648, mcs1_mcs_mat1_0_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_8653, new_AGEMA_signal_8652, new_AGEMA_signal_8651, mcs1_mcs_mat1_0_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_10507, new_AGEMA_signal_10506, new_AGEMA_signal_10505, mcs1_mcs_mat1_0_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_8653, new_AGEMA_signal_8652, new_AGEMA_signal_8651, mcs1_mcs_mat1_0_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .c ({new_AGEMA_signal_9415, new_AGEMA_signal_9414, new_AGEMA_signal_9413, mcs1_mcs_mat1_0_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_8653, new_AGEMA_signal_8652, new_AGEMA_signal_8651, mcs1_mcs_mat1_0_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_16687, new_AGEMA_signal_16686, new_AGEMA_signal_16685, mcs1_mcs_mat1_0_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .c ({new_AGEMA_signal_17425, new_AGEMA_signal_17424, new_AGEMA_signal_17423, mcs1_mcs_mat1_0_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_12886, new_AGEMA_signal_12885, new_AGEMA_signal_12884, mcs1_mcs_mat1_0_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_16687, new_AGEMA_signal_16686, new_AGEMA_signal_16685, mcs1_mcs_mat1_0_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_16690, new_AGEMA_signal_16689, new_AGEMA_signal_16688, mcs1_mcs_mat1_0_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_12886, new_AGEMA_signal_12885, new_AGEMA_signal_12884, mcs1_mcs_mat1_0_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .b ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .c ({new_AGEMA_signal_10513, new_AGEMA_signal_10512, new_AGEMA_signal_10511, mcs1_mcs_mat1_0_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .b ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_10516, new_AGEMA_signal_10515, new_AGEMA_signal_10514, mcs1_mcs_mat1_0_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({new_AGEMA_signal_11449, new_AGEMA_signal_11448, new_AGEMA_signal_11447, mcs1_mcs_mat1_0_mcs_out[87]}), .c ({new_AGEMA_signal_12889, new_AGEMA_signal_12888, new_AGEMA_signal_12887, mcs1_mcs_mat1_0_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .c ({new_AGEMA_signal_11449, new_AGEMA_signal_11448, new_AGEMA_signal_11447, mcs1_mcs_mat1_0_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .c ({new_AGEMA_signal_11458, new_AGEMA_signal_11457, new_AGEMA_signal_11456, mcs1_mcs_mat1_0_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_8656, new_AGEMA_signal_8655, new_AGEMA_signal_8654, mcs1_mcs_mat1_0_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_12904, new_AGEMA_signal_12903, new_AGEMA_signal_12902, mcs1_mcs_mat1_0_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_14356, new_AGEMA_signal_14355, new_AGEMA_signal_14354, mcs1_mcs_mat1_0_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_12904, new_AGEMA_signal_12903, new_AGEMA_signal_12902, mcs1_mcs_mat1_0_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_8659, new_AGEMA_signal_8658, new_AGEMA_signal_8657, mcs1_mcs_mat1_0_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_9424, new_AGEMA_signal_9423, new_AGEMA_signal_9422, mcs1_mcs_mat1_0_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_8659, new_AGEMA_signal_8658, new_AGEMA_signal_8657, mcs1_mcs_mat1_0_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_8662, new_AGEMA_signal_8661, new_AGEMA_signal_8660, mcs1_mcs_mat1_0_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_8665, new_AGEMA_signal_8664, new_AGEMA_signal_8663, mcs1_mcs_mat1_0_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .c ({new_AGEMA_signal_11482, new_AGEMA_signal_11481, new_AGEMA_signal_11480, mcs1_mcs_mat1_0_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_8665, new_AGEMA_signal_8664, new_AGEMA_signal_8663, mcs1_mcs_mat1_0_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_18790, new_AGEMA_signal_18789, new_AGEMA_signal_18788, mcs1_mcs_mat1_0_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_12922, new_AGEMA_signal_12921, new_AGEMA_signal_12920, mcs1_mcs_mat1_0_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_19522, new_AGEMA_signal_19521, new_AGEMA_signal_19520, mcs1_mcs_mat1_0_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_18160, new_AGEMA_signal_18159, new_AGEMA_signal_18158, mcs1_mcs_mat1_0_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_18790, new_AGEMA_signal_18789, new_AGEMA_signal_18788, mcs1_mcs_mat1_0_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_17440, new_AGEMA_signal_17439, new_AGEMA_signal_17438, mcs1_mcs_mat1_0_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_18160, new_AGEMA_signal_18159, new_AGEMA_signal_18158, mcs1_mcs_mat1_0_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_17440, new_AGEMA_signal_17439, new_AGEMA_signal_17438, mcs1_mcs_mat1_0_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_12922, new_AGEMA_signal_12921, new_AGEMA_signal_12920, mcs1_mcs_mat1_0_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_11491, new_AGEMA_signal_11490, new_AGEMA_signal_11489, mcs1_mcs_mat1_0_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_9436, new_AGEMA_signal_9435, new_AGEMA_signal_9434, mcs1_mcs_mat1_0_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_12925, new_AGEMA_signal_12924, new_AGEMA_signal_12923, mcs1_mcs_mat1_0_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_8668, new_AGEMA_signal_8667, new_AGEMA_signal_8666, mcs1_mcs_mat1_0_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .c ({new_AGEMA_signal_9436, new_AGEMA_signal_9435, new_AGEMA_signal_9434, mcs1_mcs_mat1_0_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .c ({new_AGEMA_signal_9439, new_AGEMA_signal_9438, new_AGEMA_signal_9437, mcs1_mcs_mat1_0_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .c ({new_AGEMA_signal_11491, new_AGEMA_signal_11490, new_AGEMA_signal_11489, mcs1_mcs_mat1_0_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_8668, new_AGEMA_signal_8667, new_AGEMA_signal_8666, mcs1_mcs_mat1_0_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_11494, new_AGEMA_signal_11493, new_AGEMA_signal_11492, mcs1_mcs_mat1_0_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_8668, new_AGEMA_signal_8667, new_AGEMA_signal_8666, mcs1_mcs_mat1_0_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .b ({new_AGEMA_signal_8671, new_AGEMA_signal_8670, new_AGEMA_signal_8669, mcs1_mcs_mat1_0_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_11506, new_AGEMA_signal_11505, new_AGEMA_signal_11504, mcs1_mcs_mat1_0_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_8671, new_AGEMA_signal_8670, new_AGEMA_signal_8669, mcs1_mcs_mat1_0_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({new_AGEMA_signal_11512, new_AGEMA_signal_11511, new_AGEMA_signal_11510, mcs1_mcs_mat1_0_mcs_out[51]}), .c ({new_AGEMA_signal_12940, new_AGEMA_signal_12939, new_AGEMA_signal_12938, mcs1_mcs_mat1_0_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .c ({new_AGEMA_signal_11512, new_AGEMA_signal_11511, new_AGEMA_signal_11510, mcs1_mcs_mat1_0_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_12943, new_AGEMA_signal_12942, new_AGEMA_signal_12941, mcs1_mcs_mat1_0_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_16705, new_AGEMA_signal_16704, new_AGEMA_signal_16703, mcs1_mcs_mat1_0_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_12943, new_AGEMA_signal_12942, new_AGEMA_signal_12941, mcs1_mcs_mat1_0_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_11515, new_AGEMA_signal_11514, new_AGEMA_signal_11513, mcs1_mcs_mat1_0_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_12949, new_AGEMA_signal_12948, new_AGEMA_signal_12947, mcs1_mcs_mat1_0_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .b ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_11515, new_AGEMA_signal_11514, new_AGEMA_signal_11513, mcs1_mcs_mat1_0_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_10540, new_AGEMA_signal_10539, new_AGEMA_signal_10538, mcs1_mcs_mat1_0_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_11518, new_AGEMA_signal_11517, new_AGEMA_signal_11516, mcs1_mcs_mat1_0_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .c ({new_AGEMA_signal_10540, new_AGEMA_signal_10539, new_AGEMA_signal_10538, mcs1_mcs_mat1_0_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_8674, new_AGEMA_signal_8673, new_AGEMA_signal_8672, mcs1_mcs_mat1_0_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({new_AGEMA_signal_8677, new_AGEMA_signal_8676, new_AGEMA_signal_8675, mcs1_mcs_mat1_0_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_10546, new_AGEMA_signal_10545, new_AGEMA_signal_10544, mcs1_mcs_mat1_0_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .b ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_11527, new_AGEMA_signal_11526, new_AGEMA_signal_11525, mcs1_mcs_mat1_0_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_8677, new_AGEMA_signal_8676, new_AGEMA_signal_8675, mcs1_mcs_mat1_0_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_14413, new_AGEMA_signal_14412, new_AGEMA_signal_14411, mcs1_mcs_mat1_0_mcs_out[35]}), .b ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_15793, new_AGEMA_signal_15792, new_AGEMA_signal_15791, mcs1_mcs_mat1_0_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_12967, new_AGEMA_signal_12966, new_AGEMA_signal_12965, mcs1_mcs_mat1_0_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_8680, new_AGEMA_signal_8679, new_AGEMA_signal_8678, mcs1_mcs_mat1_0_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_14413, new_AGEMA_signal_14412, new_AGEMA_signal_14411, mcs1_mcs_mat1_0_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_11533, new_AGEMA_signal_11532, new_AGEMA_signal_11531, mcs1_mcs_mat1_0_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .c ({new_AGEMA_signal_12967, new_AGEMA_signal_12966, new_AGEMA_signal_12965, mcs1_mcs_mat1_0_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .c ({new_AGEMA_signal_11533, new_AGEMA_signal_11532, new_AGEMA_signal_11531, mcs1_mcs_mat1_0_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_8680, new_AGEMA_signal_8679, new_AGEMA_signal_8678, mcs1_mcs_mat1_0_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_12970, new_AGEMA_signal_12969, new_AGEMA_signal_12968, mcs1_mcs_mat1_0_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_14416, new_AGEMA_signal_14415, new_AGEMA_signal_14414, mcs1_mcs_mat1_0_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({new_AGEMA_signal_17452, new_AGEMA_signal_17451, new_AGEMA_signal_17450, mcs1_mcs_mat1_0_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_18169, new_AGEMA_signal_18168, new_AGEMA_signal_18167, mcs1_mcs_mat1_0_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_12970, new_AGEMA_signal_12969, new_AGEMA_signal_12968, mcs1_mcs_mat1_0_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_17452, new_AGEMA_signal_17451, new_AGEMA_signal_17450, mcs1_mcs_mat1_0_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_12970, new_AGEMA_signal_12969, new_AGEMA_signal_12968, mcs1_mcs_mat1_0_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_8683, new_AGEMA_signal_8682, new_AGEMA_signal_8681, mcs1_mcs_mat1_0_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_8686, new_AGEMA_signal_8685, new_AGEMA_signal_8684, mcs1_mcs_mat1_0_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_10564, new_AGEMA_signal_10563, new_AGEMA_signal_10562, mcs1_mcs_mat1_0_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_11557, new_AGEMA_signal_11556, new_AGEMA_signal_11555, mcs1_mcs_mat1_0_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_10564, new_AGEMA_signal_10563, new_AGEMA_signal_10562, mcs1_mcs_mat1_0_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .c ({new_AGEMA_signal_11563, new_AGEMA_signal_11562, new_AGEMA_signal_11561, mcs1_mcs_mat1_0_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_8689, new_AGEMA_signal_8688, new_AGEMA_signal_8687, mcs1_mcs_mat1_0_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_13000, new_AGEMA_signal_12999, new_AGEMA_signal_12998, mcs1_mcs_mat1_0_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_8692, new_AGEMA_signal_8691, new_AGEMA_signal_8690, mcs1_mcs_mat1_0_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_8695, new_AGEMA_signal_8694, new_AGEMA_signal_8693, mcs1_mcs_mat1_0_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_10576, new_AGEMA_signal_10575, new_AGEMA_signal_10574, mcs1_mcs_mat1_0_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_8695, new_AGEMA_signal_8694, new_AGEMA_signal_8693, mcs1_mcs_mat1_0_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_9469, new_AGEMA_signal_9468, new_AGEMA_signal_9467, mcs1_mcs_mat1_0_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_8695, new_AGEMA_signal_8694, new_AGEMA_signal_8693, mcs1_mcs_mat1_0_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_11581, new_AGEMA_signal_11580, new_AGEMA_signal_11579, mcs1_mcs_mat1_0_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8698, new_AGEMA_signal_8697, new_AGEMA_signal_8696, mcs1_mcs_mat1_0_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_13012, new_AGEMA_signal_13011, new_AGEMA_signal_13010, mcs1_mcs_mat1_0_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_11581, new_AGEMA_signal_11580, new_AGEMA_signal_11579, mcs1_mcs_mat1_0_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .c ({new_AGEMA_signal_13018, new_AGEMA_signal_13017, new_AGEMA_signal_13016, mcs1_mcs_mat1_0_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_10582, new_AGEMA_signal_10581, new_AGEMA_signal_10580, mcs1_mcs_mat1_0_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_11581, new_AGEMA_signal_11580, new_AGEMA_signal_11579, mcs1_mcs_mat1_0_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_10582, new_AGEMA_signal_10581, new_AGEMA_signal_10580, mcs1_mcs_mat1_0_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .c ({new_AGEMA_signal_11584, new_AGEMA_signal_11583, new_AGEMA_signal_11582, mcs1_mcs_mat1_0_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_8698, new_AGEMA_signal_8697, new_AGEMA_signal_8696, mcs1_mcs_mat1_0_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U44 ( .a ({new_AGEMA_signal_10630, new_AGEMA_signal_10629, new_AGEMA_signal_10628, mcs1_mcs_mat1_1_mcs_out[90]}), .b ({new_AGEMA_signal_11629, new_AGEMA_signal_11628, new_AGEMA_signal_11627, mcs1_mcs_mat1_1_mcs_out[94]}), .c ({new_AGEMA_signal_13027, new_AGEMA_signal_13026, new_AGEMA_signal_13025, mcs1_mcs_mat1_1_n93}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .c ({new_AGEMA_signal_10588, new_AGEMA_signal_10587, new_AGEMA_signal_10586, mcs1_mcs_mat1_1_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .b ({new_AGEMA_signal_8701, new_AGEMA_signal_8700, new_AGEMA_signal_8699, mcs1_mcs_mat1_1_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_9478, new_AGEMA_signal_9477, new_AGEMA_signal_9476, mcs1_mcs_mat1_1_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_8701, new_AGEMA_signal_8700, new_AGEMA_signal_8699, mcs1_mcs_mat1_1_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_10597, new_AGEMA_signal_10596, new_AGEMA_signal_10595, mcs1_mcs_mat1_1_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_11596, new_AGEMA_signal_11595, new_AGEMA_signal_11594, mcs1_mcs_mat1_1_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_8704, new_AGEMA_signal_8703, new_AGEMA_signal_8702, mcs1_mcs_mat1_1_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_10597, new_AGEMA_signal_10596, new_AGEMA_signal_10595, mcs1_mcs_mat1_1_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_8704, new_AGEMA_signal_8703, new_AGEMA_signal_8702, mcs1_mcs_mat1_1_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_13045, new_AGEMA_signal_13044, new_AGEMA_signal_13043, mcs1_mcs_mat1_1_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_17488, new_AGEMA_signal_17487, new_AGEMA_signal_17486, mcs1_mcs_mat1_1_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_18199, new_AGEMA_signal_18198, new_AGEMA_signal_18197, mcs1_mcs_mat1_1_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_14488, new_AGEMA_signal_14487, new_AGEMA_signal_14486, mcs1_mcs_mat1_1_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_16765, new_AGEMA_signal_16764, new_AGEMA_signal_16763, mcs1_mcs_mat1_1_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .c ({new_AGEMA_signal_14488, new_AGEMA_signal_14487, new_AGEMA_signal_14486, mcs1_mcs_mat1_1_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .b ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_17488, new_AGEMA_signal_17487, new_AGEMA_signal_17486, mcs1_mcs_mat1_1_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_13045, new_AGEMA_signal_13044, new_AGEMA_signal_13043, mcs1_mcs_mat1_1_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_11605, new_AGEMA_signal_11604, new_AGEMA_signal_11603, mcs1_mcs_mat1_1_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_13048, new_AGEMA_signal_13047, new_AGEMA_signal_13046, mcs1_mcs_mat1_1_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_8707, new_AGEMA_signal_8706, new_AGEMA_signal_8705, mcs1_mcs_mat1_1_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_11605, new_AGEMA_signal_11604, new_AGEMA_signal_11603, mcs1_mcs_mat1_1_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_8707, new_AGEMA_signal_8706, new_AGEMA_signal_8705, mcs1_mcs_mat1_1_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_8710, new_AGEMA_signal_8709, new_AGEMA_signal_8708, mcs1_mcs_mat1_1_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({new_AGEMA_signal_10615, new_AGEMA_signal_10614, new_AGEMA_signal_10613, mcs1_mcs_mat1_1_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_11617, new_AGEMA_signal_11616, new_AGEMA_signal_11615, mcs1_mcs_mat1_1_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, new_AGEMA_signal_8711, mcs1_mcs_mat1_1_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_10615, new_AGEMA_signal_10614, new_AGEMA_signal_10613, mcs1_mcs_mat1_1_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .b ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .c ({new_AGEMA_signal_11620, new_AGEMA_signal_11619, new_AGEMA_signal_11618, mcs1_mcs_mat1_1_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, new_AGEMA_signal_8711, mcs1_mcs_mat1_1_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_13069, new_AGEMA_signal_13068, new_AGEMA_signal_13067, mcs1_mcs_mat1_1_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_16771, new_AGEMA_signal_16770, new_AGEMA_signal_16769, mcs1_mcs_mat1_1_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_13069, new_AGEMA_signal_13068, new_AGEMA_signal_13067, mcs1_mcs_mat1_1_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .c ({new_AGEMA_signal_14518, new_AGEMA_signal_14517, new_AGEMA_signal_14516, mcs1_mcs_mat1_1_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_13069, new_AGEMA_signal_13068, new_AGEMA_signal_13067, mcs1_mcs_mat1_1_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_10621, new_AGEMA_signal_10620, new_AGEMA_signal_10619, mcs1_mcs_mat1_1_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .c ({new_AGEMA_signal_11629, new_AGEMA_signal_11628, new_AGEMA_signal_11627, mcs1_mcs_mat1_1_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_8716, new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_1_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_10621, new_AGEMA_signal_10620, new_AGEMA_signal_10619, mcs1_mcs_mat1_1_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_10624, new_AGEMA_signal_10623, new_AGEMA_signal_10622, mcs1_mcs_mat1_1_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({new_AGEMA_signal_8716, new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_1_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .b ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .c ({new_AGEMA_signal_10630, new_AGEMA_signal_10629, new_AGEMA_signal_10628, mcs1_mcs_mat1_1_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .b ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_10633, new_AGEMA_signal_10632, new_AGEMA_signal_10631, mcs1_mcs_mat1_1_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({new_AGEMA_signal_11638, new_AGEMA_signal_11637, new_AGEMA_signal_11636, mcs1_mcs_mat1_1_mcs_out[87]}), .c ({new_AGEMA_signal_13075, new_AGEMA_signal_13074, new_AGEMA_signal_13073, mcs1_mcs_mat1_1_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .c ({new_AGEMA_signal_11638, new_AGEMA_signal_11637, new_AGEMA_signal_11636, mcs1_mcs_mat1_1_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .c ({new_AGEMA_signal_17503, new_AGEMA_signal_17502, new_AGEMA_signal_17501, mcs1_mcs_mat1_1_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_13078, new_AGEMA_signal_13077, new_AGEMA_signal_13076, mcs1_mcs_mat1_1_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, new_AGEMA_signal_8717, mcs1_mcs_mat1_1_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, new_AGEMA_signal_9497, mcs1_mcs_mat1_1_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, new_AGEMA_signal_8717, mcs1_mcs_mat1_1_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_8722, new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_1_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, new_AGEMA_signal_9503, mcs1_mcs_mat1_1_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_8722, new_AGEMA_signal_8721, new_AGEMA_signal_8720, mcs1_mcs_mat1_1_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, new_AGEMA_signal_8723, mcs1_mcs_mat1_1_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_13096, new_AGEMA_signal_13095, new_AGEMA_signal_13094, mcs1_mcs_mat1_1_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .c ({new_AGEMA_signal_17509, new_AGEMA_signal_17508, new_AGEMA_signal_17507, mcs1_mcs_mat1_1_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_13096, new_AGEMA_signal_13095, new_AGEMA_signal_13094, mcs1_mcs_mat1_1_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_14560, new_AGEMA_signal_14559, new_AGEMA_signal_14558, mcs1_mcs_mat1_1_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_8728, new_AGEMA_signal_8727, new_AGEMA_signal_8726, mcs1_mcs_mat1_1_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_15895, new_AGEMA_signal_15894, new_AGEMA_signal_15893, mcs1_mcs_mat1_1_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_13105, new_AGEMA_signal_13104, new_AGEMA_signal_13103, mcs1_mcs_mat1_1_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_14560, new_AGEMA_signal_14559, new_AGEMA_signal_14558, mcs1_mcs_mat1_1_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_11665, new_AGEMA_signal_11664, new_AGEMA_signal_11663, mcs1_mcs_mat1_1_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_13105, new_AGEMA_signal_13104, new_AGEMA_signal_13103, mcs1_mcs_mat1_1_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_11665, new_AGEMA_signal_11664, new_AGEMA_signal_11663, mcs1_mcs_mat1_1_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({new_AGEMA_signal_8728, new_AGEMA_signal_8727, new_AGEMA_signal_8726, mcs1_mcs_mat1_1_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_11674, new_AGEMA_signal_11673, new_AGEMA_signal_11672, mcs1_mcs_mat1_1_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_9517, new_AGEMA_signal_9516, new_AGEMA_signal_9515, mcs1_mcs_mat1_1_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_13108, new_AGEMA_signal_13107, new_AGEMA_signal_13106, mcs1_mcs_mat1_1_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, new_AGEMA_signal_8729, mcs1_mcs_mat1_1_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .c ({new_AGEMA_signal_9517, new_AGEMA_signal_9516, new_AGEMA_signal_9515, mcs1_mcs_mat1_1_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .c ({new_AGEMA_signal_9520, new_AGEMA_signal_9519, new_AGEMA_signal_9518, mcs1_mcs_mat1_1_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .c ({new_AGEMA_signal_11674, new_AGEMA_signal_11673, new_AGEMA_signal_11672, mcs1_mcs_mat1_1_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, new_AGEMA_signal_8729, mcs1_mcs_mat1_1_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_11677, new_AGEMA_signal_11676, new_AGEMA_signal_11675, mcs1_mcs_mat1_1_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_8731, new_AGEMA_signal_8730, new_AGEMA_signal_8729, mcs1_mcs_mat1_1_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .b ({new_AGEMA_signal_8734, new_AGEMA_signal_8733, new_AGEMA_signal_8732, mcs1_mcs_mat1_1_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_11689, new_AGEMA_signal_11688, new_AGEMA_signal_11687, mcs1_mcs_mat1_1_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({new_AGEMA_signal_8734, new_AGEMA_signal_8733, new_AGEMA_signal_8732, mcs1_mcs_mat1_1_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({new_AGEMA_signal_17515, new_AGEMA_signal_17514, new_AGEMA_signal_17513, mcs1_mcs_mat1_1_mcs_out[51]}), .c ({new_AGEMA_signal_18226, new_AGEMA_signal_18225, new_AGEMA_signal_18224, mcs1_mcs_mat1_1_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .c ({new_AGEMA_signal_17515, new_AGEMA_signal_17514, new_AGEMA_signal_17513, mcs1_mcs_mat1_1_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, new_AGEMA_signal_8735, mcs1_mcs_mat1_1_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_10657, new_AGEMA_signal_10656, new_AGEMA_signal_10655, mcs1_mcs_mat1_1_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, new_AGEMA_signal_8735, mcs1_mcs_mat1_1_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_11701, new_AGEMA_signal_11700, new_AGEMA_signal_11699, mcs1_mcs_mat1_1_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_13129, new_AGEMA_signal_13128, new_AGEMA_signal_13127, mcs1_mcs_mat1_1_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_11701, new_AGEMA_signal_11700, new_AGEMA_signal_11699, mcs1_mcs_mat1_1_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_10663, new_AGEMA_signal_10662, new_AGEMA_signal_10661, mcs1_mcs_mat1_1_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_11704, new_AGEMA_signal_11703, new_AGEMA_signal_11702, mcs1_mcs_mat1_1_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .c ({new_AGEMA_signal_10663, new_AGEMA_signal_10662, new_AGEMA_signal_10661, mcs1_mcs_mat1_1_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({new_AGEMA_signal_8740, new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_1_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, new_AGEMA_signal_8741, mcs1_mcs_mat1_1_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_10669, new_AGEMA_signal_10668, new_AGEMA_signal_10667, mcs1_mcs_mat1_1_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_11713, new_AGEMA_signal_11712, new_AGEMA_signal_11711, mcs1_mcs_mat1_1_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, new_AGEMA_signal_8741, mcs1_mcs_mat1_1_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_18874, new_AGEMA_signal_18873, new_AGEMA_signal_18872, mcs1_mcs_mat1_1_mcs_out[35]}), .b ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_19606, new_AGEMA_signal_19605, new_AGEMA_signal_19604, mcs1_mcs_mat1_1_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_18232, new_AGEMA_signal_18231, new_AGEMA_signal_18230, mcs1_mcs_mat1_1_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_13144, new_AGEMA_signal_13143, new_AGEMA_signal_13142, mcs1_mcs_mat1_1_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_18874, new_AGEMA_signal_18873, new_AGEMA_signal_18872, mcs1_mcs_mat1_1_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_17518, new_AGEMA_signal_17517, new_AGEMA_signal_17516, mcs1_mcs_mat1_1_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .c ({new_AGEMA_signal_18232, new_AGEMA_signal_18231, new_AGEMA_signal_18230, mcs1_mcs_mat1_1_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .c ({new_AGEMA_signal_17518, new_AGEMA_signal_17517, new_AGEMA_signal_17516, mcs1_mcs_mat1_1_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({new_AGEMA_signal_13144, new_AGEMA_signal_13143, new_AGEMA_signal_13142, mcs1_mcs_mat1_1_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_8746, new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_9538, new_AGEMA_signal_9537, new_AGEMA_signal_9536, mcs1_mcs_mat1_1_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({new_AGEMA_signal_11719, new_AGEMA_signal_11718, new_AGEMA_signal_11717, mcs1_mcs_mat1_1_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_13150, new_AGEMA_signal_13149, new_AGEMA_signal_13148, mcs1_mcs_mat1_1_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_8746, new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_11719, new_AGEMA_signal_11718, new_AGEMA_signal_11717, mcs1_mcs_mat1_1_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({new_AGEMA_signal_8746, new_AGEMA_signal_8745, new_AGEMA_signal_8744, mcs1_mcs_mat1_1_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, new_AGEMA_signal_8747, mcs1_mcs_mat1_1_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({new_AGEMA_signal_8752, new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_1_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_16789, new_AGEMA_signal_16788, new_AGEMA_signal_16787, mcs1_mcs_mat1_1_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_17524, new_AGEMA_signal_17523, new_AGEMA_signal_17522, mcs1_mcs_mat1_1_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_16789, new_AGEMA_signal_16788, new_AGEMA_signal_16787, mcs1_mcs_mat1_1_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .c ({new_AGEMA_signal_17530, new_AGEMA_signal_17529, new_AGEMA_signal_17528, mcs1_mcs_mat1_1_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({new_AGEMA_signal_13174, new_AGEMA_signal_13173, new_AGEMA_signal_13172, mcs1_mcs_mat1_1_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, new_AGEMA_signal_8753, mcs1_mcs_mat1_1_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({new_AGEMA_signal_8758, new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_1_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_8761, new_AGEMA_signal_8760, new_AGEMA_signal_8759, mcs1_mcs_mat1_1_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_10696, new_AGEMA_signal_10695, new_AGEMA_signal_10694, mcs1_mcs_mat1_1_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_8761, new_AGEMA_signal_8760, new_AGEMA_signal_8759, mcs1_mcs_mat1_1_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_9556, new_AGEMA_signal_9555, new_AGEMA_signal_9554, mcs1_mcs_mat1_1_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({new_AGEMA_signal_8761, new_AGEMA_signal_8760, new_AGEMA_signal_8759, mcs1_mcs_mat1_1_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_17542, new_AGEMA_signal_17541, new_AGEMA_signal_17540, mcs1_mcs_mat1_1_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_13195, new_AGEMA_signal_13194, new_AGEMA_signal_13193, mcs1_mcs_mat1_1_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_18244, new_AGEMA_signal_18243, new_AGEMA_signal_18242, mcs1_mcs_mat1_1_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_17542, new_AGEMA_signal_17541, new_AGEMA_signal_17540, mcs1_mcs_mat1_1_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .c ({new_AGEMA_signal_18250, new_AGEMA_signal_18249, new_AGEMA_signal_18248, mcs1_mcs_mat1_1_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_16801, new_AGEMA_signal_16800, new_AGEMA_signal_16799, mcs1_mcs_mat1_1_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_17542, new_AGEMA_signal_17541, new_AGEMA_signal_17540, mcs1_mcs_mat1_1_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_16801, new_AGEMA_signal_16800, new_AGEMA_signal_16799, mcs1_mcs_mat1_1_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .c ({new_AGEMA_signal_17545, new_AGEMA_signal_17544, new_AGEMA_signal_17543, mcs1_mcs_mat1_1_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({new_AGEMA_signal_13195, new_AGEMA_signal_13194, new_AGEMA_signal_13193, mcs1_mcs_mat1_1_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U44 ( .a ({new_AGEMA_signal_10741, new_AGEMA_signal_10740, new_AGEMA_signal_10739, mcs1_mcs_mat1_2_mcs_out[90]}), .b ({new_AGEMA_signal_11791, new_AGEMA_signal_11790, new_AGEMA_signal_11789, mcs1_mcs_mat1_2_mcs_out[94]}), .c ({new_AGEMA_signal_13201, new_AGEMA_signal_13200, new_AGEMA_signal_13199, mcs1_mcs_mat1_2_n93}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .c ({new_AGEMA_signal_10702, new_AGEMA_signal_10701, new_AGEMA_signal_10700, mcs1_mcs_mat1_2_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .b ({new_AGEMA_signal_8764, new_AGEMA_signal_8763, new_AGEMA_signal_8762, mcs1_mcs_mat1_2_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_9562, new_AGEMA_signal_9561, new_AGEMA_signal_9560, mcs1_mcs_mat1_2_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({new_AGEMA_signal_8764, new_AGEMA_signal_8763, new_AGEMA_signal_8762, mcs1_mcs_mat1_2_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_16849, new_AGEMA_signal_16848, new_AGEMA_signal_16847, mcs1_mcs_mat1_2_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_17563, new_AGEMA_signal_17562, new_AGEMA_signal_17561, mcs1_mcs_mat1_2_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_13213, new_AGEMA_signal_13212, new_AGEMA_signal_13211, mcs1_mcs_mat1_2_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_16849, new_AGEMA_signal_16848, new_AGEMA_signal_16847, mcs1_mcs_mat1_2_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({new_AGEMA_signal_13213, new_AGEMA_signal_13212, new_AGEMA_signal_13211, mcs1_mcs_mat1_2_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_8767, new_AGEMA_signal_8766, new_AGEMA_signal_8765, mcs1_mcs_mat1_2_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_11770, new_AGEMA_signal_11769, new_AGEMA_signal_11768, mcs1_mcs_mat1_2_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_13216, new_AGEMA_signal_13215, new_AGEMA_signal_13214, mcs1_mcs_mat1_2_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_9568, new_AGEMA_signal_9567, new_AGEMA_signal_9566, mcs1_mcs_mat1_2_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_10711, new_AGEMA_signal_10710, new_AGEMA_signal_10709, mcs1_mcs_mat1_2_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .c ({new_AGEMA_signal_9568, new_AGEMA_signal_9567, new_AGEMA_signal_9566, mcs1_mcs_mat1_2_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_11770, new_AGEMA_signal_11769, new_AGEMA_signal_11768, mcs1_mcs_mat1_2_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({new_AGEMA_signal_8767, new_AGEMA_signal_8766, new_AGEMA_signal_8765, mcs1_mcs_mat1_2_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_11776, new_AGEMA_signal_11775, new_AGEMA_signal_11774, mcs1_mcs_mat1_2_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_13225, new_AGEMA_signal_13224, new_AGEMA_signal_13223, mcs1_mcs_mat1_2_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_8770, new_AGEMA_signal_8769, new_AGEMA_signal_8768, mcs1_mcs_mat1_2_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_11776, new_AGEMA_signal_11775, new_AGEMA_signal_11774, mcs1_mcs_mat1_2_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({new_AGEMA_signal_8770, new_AGEMA_signal_8769, new_AGEMA_signal_8768, mcs1_mcs_mat1_2_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({new_AGEMA_signal_8773, new_AGEMA_signal_8772, new_AGEMA_signal_8771, mcs1_mcs_mat1_2_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({new_AGEMA_signal_16858, new_AGEMA_signal_16857, new_AGEMA_signal_16856, mcs1_mcs_mat1_2_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_17572, new_AGEMA_signal_17571, new_AGEMA_signal_17570, mcs1_mcs_mat1_2_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_13237, new_AGEMA_signal_13236, new_AGEMA_signal_13235, mcs1_mcs_mat1_2_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_16858, new_AGEMA_signal_16857, new_AGEMA_signal_16856, mcs1_mcs_mat1_2_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .b ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .c ({new_AGEMA_signal_17575, new_AGEMA_signal_17574, new_AGEMA_signal_17573, mcs1_mcs_mat1_2_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({new_AGEMA_signal_13237, new_AGEMA_signal_13236, new_AGEMA_signal_13235, mcs1_mcs_mat1_2_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_8776, new_AGEMA_signal_8775, new_AGEMA_signal_8774, mcs1_mcs_mat1_2_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_10726, new_AGEMA_signal_10725, new_AGEMA_signal_10724, mcs1_mcs_mat1_2_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_8776, new_AGEMA_signal_8775, new_AGEMA_signal_8774, mcs1_mcs_mat1_2_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .c ({new_AGEMA_signal_9580, new_AGEMA_signal_9579, new_AGEMA_signal_9578, mcs1_mcs_mat1_2_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({new_AGEMA_signal_8776, new_AGEMA_signal_8775, new_AGEMA_signal_8774, mcs1_mcs_mat1_2_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_10732, new_AGEMA_signal_10731, new_AGEMA_signal_10730, mcs1_mcs_mat1_2_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .c ({new_AGEMA_signal_11791, new_AGEMA_signal_11790, new_AGEMA_signal_11789, mcs1_mcs_mat1_2_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_8779, new_AGEMA_signal_8778, new_AGEMA_signal_8777, mcs1_mcs_mat1_2_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_10732, new_AGEMA_signal_10731, new_AGEMA_signal_10730, mcs1_mcs_mat1_2_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_10735, new_AGEMA_signal_10734, new_AGEMA_signal_10733, mcs1_mcs_mat1_2_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({new_AGEMA_signal_8779, new_AGEMA_signal_8778, new_AGEMA_signal_8777, mcs1_mcs_mat1_2_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .b ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .c ({new_AGEMA_signal_10741, new_AGEMA_signal_10740, new_AGEMA_signal_10739, mcs1_mcs_mat1_2_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .b ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_10744, new_AGEMA_signal_10743, new_AGEMA_signal_10742, mcs1_mcs_mat1_2_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({new_AGEMA_signal_17587, new_AGEMA_signal_17586, new_AGEMA_signal_17585, mcs1_mcs_mat1_2_mcs_out[87]}), .c ({new_AGEMA_signal_18286, new_AGEMA_signal_18285, new_AGEMA_signal_18284, mcs1_mcs_mat1_2_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .c ({new_AGEMA_signal_17587, new_AGEMA_signal_17586, new_AGEMA_signal_17585, mcs1_mcs_mat1_2_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .c ({new_AGEMA_signal_11806, new_AGEMA_signal_11805, new_AGEMA_signal_11804, mcs1_mcs_mat1_2_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({new_AGEMA_signal_8782, new_AGEMA_signal_8781, new_AGEMA_signal_8780, mcs1_mcs_mat1_2_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_8785, new_AGEMA_signal_8784, new_AGEMA_signal_8783, mcs1_mcs_mat1_2_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_9592, new_AGEMA_signal_9591, new_AGEMA_signal_9590, mcs1_mcs_mat1_2_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({new_AGEMA_signal_8785, new_AGEMA_signal_8784, new_AGEMA_signal_8783, mcs1_mcs_mat1_2_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_8788, new_AGEMA_signal_8787, new_AGEMA_signal_8786, mcs1_mcs_mat1_2_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_9598, new_AGEMA_signal_9597, new_AGEMA_signal_9596, mcs1_mcs_mat1_2_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({new_AGEMA_signal_8788, new_AGEMA_signal_8787, new_AGEMA_signal_8786, mcs1_mcs_mat1_2_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({new_AGEMA_signal_13267, new_AGEMA_signal_13266, new_AGEMA_signal_13265, mcs1_mcs_mat1_2_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_8791, new_AGEMA_signal_8790, new_AGEMA_signal_8789, mcs1_mcs_mat1_2_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .c ({new_AGEMA_signal_11827, new_AGEMA_signal_11826, new_AGEMA_signal_11825, mcs1_mcs_mat1_2_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({new_AGEMA_signal_8791, new_AGEMA_signal_8790, new_AGEMA_signal_8789, mcs1_mcs_mat1_2_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_14725, new_AGEMA_signal_14724, new_AGEMA_signal_14723, mcs1_mcs_mat1_2_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_8794, new_AGEMA_signal_8793, new_AGEMA_signal_8792, mcs1_mcs_mat1_2_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_16018, new_AGEMA_signal_16017, new_AGEMA_signal_16016, mcs1_mcs_mat1_2_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_13279, new_AGEMA_signal_13278, new_AGEMA_signal_13277, mcs1_mcs_mat1_2_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_14725, new_AGEMA_signal_14724, new_AGEMA_signal_14723, mcs1_mcs_mat1_2_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_11833, new_AGEMA_signal_11832, new_AGEMA_signal_11831, mcs1_mcs_mat1_2_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_13279, new_AGEMA_signal_13278, new_AGEMA_signal_13277, mcs1_mcs_mat1_2_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_11833, new_AGEMA_signal_11832, new_AGEMA_signal_11831, mcs1_mcs_mat1_2_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({new_AGEMA_signal_8794, new_AGEMA_signal_8793, new_AGEMA_signal_8792, mcs1_mcs_mat1_2_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_11842, new_AGEMA_signal_11841, new_AGEMA_signal_11840, mcs1_mcs_mat1_2_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_9610, new_AGEMA_signal_9609, new_AGEMA_signal_9608, mcs1_mcs_mat1_2_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_13282, new_AGEMA_signal_13281, new_AGEMA_signal_13280, mcs1_mcs_mat1_2_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_8797, new_AGEMA_signal_8796, new_AGEMA_signal_8795, mcs1_mcs_mat1_2_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .c ({new_AGEMA_signal_9610, new_AGEMA_signal_9609, new_AGEMA_signal_9608, mcs1_mcs_mat1_2_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .c ({new_AGEMA_signal_9613, new_AGEMA_signal_9612, new_AGEMA_signal_9611, mcs1_mcs_mat1_2_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .c ({new_AGEMA_signal_11842, new_AGEMA_signal_11841, new_AGEMA_signal_11840, mcs1_mcs_mat1_2_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_8797, new_AGEMA_signal_8796, new_AGEMA_signal_8795, mcs1_mcs_mat1_2_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_11845, new_AGEMA_signal_11844, new_AGEMA_signal_11843, mcs1_mcs_mat1_2_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({new_AGEMA_signal_8797, new_AGEMA_signal_8796, new_AGEMA_signal_8795, mcs1_mcs_mat1_2_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .b ({new_AGEMA_signal_13291, new_AGEMA_signal_13290, new_AGEMA_signal_13289, mcs1_mcs_mat1_2_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_17605, new_AGEMA_signal_17604, new_AGEMA_signal_17603, mcs1_mcs_mat1_2_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({new_AGEMA_signal_13291, new_AGEMA_signal_13290, new_AGEMA_signal_13289, mcs1_mcs_mat1_2_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({new_AGEMA_signal_11851, new_AGEMA_signal_11850, new_AGEMA_signal_11849, mcs1_mcs_mat1_2_mcs_out[51]}), .c ({new_AGEMA_signal_13294, new_AGEMA_signal_13293, new_AGEMA_signal_13292, mcs1_mcs_mat1_2_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .c ({new_AGEMA_signal_11851, new_AGEMA_signal_11850, new_AGEMA_signal_11849, mcs1_mcs_mat1_2_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_8800, new_AGEMA_signal_8799, new_AGEMA_signal_8798, mcs1_mcs_mat1_2_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_10765, new_AGEMA_signal_10764, new_AGEMA_signal_10763, mcs1_mcs_mat1_2_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({new_AGEMA_signal_8800, new_AGEMA_signal_8799, new_AGEMA_signal_8798, mcs1_mcs_mat1_2_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_11860, new_AGEMA_signal_11859, new_AGEMA_signal_11858, mcs1_mcs_mat1_2_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_13303, new_AGEMA_signal_13302, new_AGEMA_signal_13301, mcs1_mcs_mat1_2_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .b ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_11860, new_AGEMA_signal_11859, new_AGEMA_signal_11858, mcs1_mcs_mat1_2_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_10771, new_AGEMA_signal_10770, new_AGEMA_signal_10769, mcs1_mcs_mat1_2_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_11863, new_AGEMA_signal_11862, new_AGEMA_signal_11861, mcs1_mcs_mat1_2_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .c ({new_AGEMA_signal_10771, new_AGEMA_signal_10770, new_AGEMA_signal_10769, mcs1_mcs_mat1_2_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({new_AGEMA_signal_8803, new_AGEMA_signal_8802, new_AGEMA_signal_8801, mcs1_mcs_mat1_2_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({new_AGEMA_signal_13312, new_AGEMA_signal_13311, new_AGEMA_signal_13310, mcs1_mcs_mat1_2_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_16882, new_AGEMA_signal_16881, new_AGEMA_signal_16880, mcs1_mcs_mat1_2_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .b ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_17614, new_AGEMA_signal_17613, new_AGEMA_signal_17612, mcs1_mcs_mat1_2_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({new_AGEMA_signal_13312, new_AGEMA_signal_13311, new_AGEMA_signal_13310, mcs1_mcs_mat1_2_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_14749, new_AGEMA_signal_14748, new_AGEMA_signal_14747, mcs1_mcs_mat1_2_mcs_out[35]}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_16027, new_AGEMA_signal_16026, new_AGEMA_signal_16025, mcs1_mcs_mat1_2_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_13318, new_AGEMA_signal_13317, new_AGEMA_signal_13316, mcs1_mcs_mat1_2_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_8806, new_AGEMA_signal_8805, new_AGEMA_signal_8804, mcs1_mcs_mat1_2_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_14749, new_AGEMA_signal_14748, new_AGEMA_signal_14747, mcs1_mcs_mat1_2_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_11869, new_AGEMA_signal_11868, new_AGEMA_signal_11867, mcs1_mcs_mat1_2_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .c ({new_AGEMA_signal_13318, new_AGEMA_signal_13317, new_AGEMA_signal_13316, mcs1_mcs_mat1_2_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .c ({new_AGEMA_signal_11869, new_AGEMA_signal_11868, new_AGEMA_signal_11867, mcs1_mcs_mat1_2_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({new_AGEMA_signal_8806, new_AGEMA_signal_8805, new_AGEMA_signal_8804, mcs1_mcs_mat1_2_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_8809, new_AGEMA_signal_8808, new_AGEMA_signal_8807, mcs1_mcs_mat1_2_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_9628, new_AGEMA_signal_9627, new_AGEMA_signal_9626, mcs1_mcs_mat1_2_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({new_AGEMA_signal_11875, new_AGEMA_signal_11874, new_AGEMA_signal_11873, mcs1_mcs_mat1_2_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_13324, new_AGEMA_signal_13323, new_AGEMA_signal_13322, mcs1_mcs_mat1_2_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_8809, new_AGEMA_signal_8808, new_AGEMA_signal_8807, mcs1_mcs_mat1_2_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_11875, new_AGEMA_signal_11874, new_AGEMA_signal_11873, mcs1_mcs_mat1_2_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({new_AGEMA_signal_8809, new_AGEMA_signal_8808, new_AGEMA_signal_8807, mcs1_mcs_mat1_2_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({new_AGEMA_signal_8812, new_AGEMA_signal_8811, new_AGEMA_signal_8810, mcs1_mcs_mat1_2_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({new_AGEMA_signal_13339, new_AGEMA_signal_13338, new_AGEMA_signal_13337, mcs1_mcs_mat1_2_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_10786, new_AGEMA_signal_10785, new_AGEMA_signal_10784, mcs1_mcs_mat1_2_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_11893, new_AGEMA_signal_11892, new_AGEMA_signal_11891, mcs1_mcs_mat1_2_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_10786, new_AGEMA_signal_10785, new_AGEMA_signal_10784, mcs1_mcs_mat1_2_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .c ({new_AGEMA_signal_11899, new_AGEMA_signal_11898, new_AGEMA_signal_11897, mcs1_mcs_mat1_2_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({new_AGEMA_signal_8815, new_AGEMA_signal_8814, new_AGEMA_signal_8813, mcs1_mcs_mat1_2_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({new_AGEMA_signal_8818, new_AGEMA_signal_8817, new_AGEMA_signal_8816, mcs1_mcs_mat1_2_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({new_AGEMA_signal_8821, new_AGEMA_signal_8820, new_AGEMA_signal_8819, mcs1_mcs_mat1_2_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_13366, new_AGEMA_signal_13365, new_AGEMA_signal_13364, mcs1_mcs_mat1_2_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_16900, new_AGEMA_signal_16899, new_AGEMA_signal_16898, mcs1_mcs_mat1_2_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_13366, new_AGEMA_signal_13365, new_AGEMA_signal_13364, mcs1_mcs_mat1_2_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_14791, new_AGEMA_signal_14790, new_AGEMA_signal_14789, mcs1_mcs_mat1_2_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({new_AGEMA_signal_13366, new_AGEMA_signal_13365, new_AGEMA_signal_13364, mcs1_mcs_mat1_2_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_11920, new_AGEMA_signal_11919, new_AGEMA_signal_11918, mcs1_mcs_mat1_2_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8824, new_AGEMA_signal_8823, new_AGEMA_signal_8822, mcs1_mcs_mat1_2_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_13369, new_AGEMA_signal_13368, new_AGEMA_signal_13367, mcs1_mcs_mat1_2_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_11920, new_AGEMA_signal_11919, new_AGEMA_signal_11918, mcs1_mcs_mat1_2_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .c ({new_AGEMA_signal_13375, new_AGEMA_signal_13374, new_AGEMA_signal_13373, mcs1_mcs_mat1_2_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_10801, new_AGEMA_signal_10800, new_AGEMA_signal_10799, mcs1_mcs_mat1_2_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_11920, new_AGEMA_signal_11919, new_AGEMA_signal_11918, mcs1_mcs_mat1_2_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_10801, new_AGEMA_signal_10800, new_AGEMA_signal_10799, mcs1_mcs_mat1_2_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .c ({new_AGEMA_signal_11923, new_AGEMA_signal_11922, new_AGEMA_signal_11921, mcs1_mcs_mat1_2_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({new_AGEMA_signal_8824, new_AGEMA_signal_8823, new_AGEMA_signal_8822, mcs1_mcs_mat1_2_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U44 ( .a ({new_AGEMA_signal_16969, new_AGEMA_signal_16968, new_AGEMA_signal_16967, mcs1_mcs_mat1_3_mcs_out[90]}), .b ({new_AGEMA_signal_11968, new_AGEMA_signal_11967, new_AGEMA_signal_11966, mcs1_mcs_mat1_3_mcs_out[94]}), .c ({new_AGEMA_signal_17641, new_AGEMA_signal_17640, new_AGEMA_signal_17639, mcs1_mcs_mat1_3_n93}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .c ({new_AGEMA_signal_10807, new_AGEMA_signal_10806, new_AGEMA_signal_10805, mcs1_mcs_mat1_3_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .b ({new_AGEMA_signal_13381, new_AGEMA_signal_13380, new_AGEMA_signal_13379, mcs1_mcs_mat1_3_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_14824, new_AGEMA_signal_14823, new_AGEMA_signal_14822, mcs1_mcs_mat1_3_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({new_AGEMA_signal_13381, new_AGEMA_signal_13380, new_AGEMA_signal_13379, mcs1_mcs_mat1_3_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_10810, new_AGEMA_signal_10809, new_AGEMA_signal_10808, mcs1_mcs_mat1_3_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_11929, new_AGEMA_signal_11928, new_AGEMA_signal_11927, mcs1_mcs_mat1_3_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_8827, new_AGEMA_signal_8826, new_AGEMA_signal_8825, mcs1_mcs_mat1_3_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_10810, new_AGEMA_signal_10809, new_AGEMA_signal_10808, mcs1_mcs_mat1_3_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({new_AGEMA_signal_8827, new_AGEMA_signal_8826, new_AGEMA_signal_8825, mcs1_mcs_mat1_3_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_8830, new_AGEMA_signal_8829, new_AGEMA_signal_8828, mcs1_mcs_mat1_3_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_11941, new_AGEMA_signal_11940, new_AGEMA_signal_11939, mcs1_mcs_mat1_3_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_13390, new_AGEMA_signal_13389, new_AGEMA_signal_13388, mcs1_mcs_mat1_3_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_9652, new_AGEMA_signal_9651, new_AGEMA_signal_9650, mcs1_mcs_mat1_3_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_10819, new_AGEMA_signal_10818, new_AGEMA_signal_10817, mcs1_mcs_mat1_3_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .c ({new_AGEMA_signal_9652, new_AGEMA_signal_9651, new_AGEMA_signal_9650, mcs1_mcs_mat1_3_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .b ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_11941, new_AGEMA_signal_11940, new_AGEMA_signal_11939, mcs1_mcs_mat1_3_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({new_AGEMA_signal_8830, new_AGEMA_signal_8829, new_AGEMA_signal_8828, mcs1_mcs_mat1_3_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_11947, new_AGEMA_signal_11946, new_AGEMA_signal_11945, mcs1_mcs_mat1_3_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_13399, new_AGEMA_signal_13398, new_AGEMA_signal_13397, mcs1_mcs_mat1_3_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_8833, new_AGEMA_signal_8832, new_AGEMA_signal_8831, mcs1_mcs_mat1_3_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_11947, new_AGEMA_signal_11946, new_AGEMA_signal_11945, mcs1_mcs_mat1_3_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({new_AGEMA_signal_8833, new_AGEMA_signal_8832, new_AGEMA_signal_8831, mcs1_mcs_mat1_3_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({new_AGEMA_signal_13405, new_AGEMA_signal_13404, new_AGEMA_signal_13403, mcs1_mcs_mat1_3_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({new_AGEMA_signal_10828, new_AGEMA_signal_10827, new_AGEMA_signal_10826, mcs1_mcs_mat1_3_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_11953, new_AGEMA_signal_11952, new_AGEMA_signal_11951, mcs1_mcs_mat1_3_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_8836, new_AGEMA_signal_8835, new_AGEMA_signal_8834, mcs1_mcs_mat1_3_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_10828, new_AGEMA_signal_10827, new_AGEMA_signal_10826, mcs1_mcs_mat1_3_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .b ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .c ({new_AGEMA_signal_11956, new_AGEMA_signal_11955, new_AGEMA_signal_11954, mcs1_mcs_mat1_3_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({new_AGEMA_signal_8836, new_AGEMA_signal_8835, new_AGEMA_signal_8834, mcs1_mcs_mat1_3_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_8839, new_AGEMA_signal_8838, new_AGEMA_signal_8837, mcs1_mcs_mat1_3_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_10834, new_AGEMA_signal_10833, new_AGEMA_signal_10832, mcs1_mcs_mat1_3_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_8839, new_AGEMA_signal_8838, new_AGEMA_signal_8837, mcs1_mcs_mat1_3_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .c ({new_AGEMA_signal_9664, new_AGEMA_signal_9663, new_AGEMA_signal_9662, mcs1_mcs_mat1_3_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({new_AGEMA_signal_8839, new_AGEMA_signal_8838, new_AGEMA_signal_8837, mcs1_mcs_mat1_3_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_10840, new_AGEMA_signal_10839, new_AGEMA_signal_10838, mcs1_mcs_mat1_3_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .c ({new_AGEMA_signal_11968, new_AGEMA_signal_11967, new_AGEMA_signal_11966, mcs1_mcs_mat1_3_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_8842, new_AGEMA_signal_8841, new_AGEMA_signal_8840, mcs1_mcs_mat1_3_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_10840, new_AGEMA_signal_10839, new_AGEMA_signal_10838, mcs1_mcs_mat1_3_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_10843, new_AGEMA_signal_10842, new_AGEMA_signal_10841, mcs1_mcs_mat1_3_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({new_AGEMA_signal_8842, new_AGEMA_signal_8841, new_AGEMA_signal_8840, mcs1_mcs_mat1_3_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .b ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .c ({new_AGEMA_signal_16969, new_AGEMA_signal_16968, new_AGEMA_signal_16967, mcs1_mcs_mat1_3_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .b ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_16972, new_AGEMA_signal_16971, new_AGEMA_signal_16970, mcs1_mcs_mat1_3_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({new_AGEMA_signal_11977, new_AGEMA_signal_11976, new_AGEMA_signal_11975, mcs1_mcs_mat1_3_mcs_out[87]}), .c ({new_AGEMA_signal_13423, new_AGEMA_signal_13422, new_AGEMA_signal_13421, mcs1_mcs_mat1_3_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .c ({new_AGEMA_signal_11977, new_AGEMA_signal_11976, new_AGEMA_signal_11975, mcs1_mcs_mat1_3_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .c ({new_AGEMA_signal_11986, new_AGEMA_signal_11985, new_AGEMA_signal_11984, mcs1_mcs_mat1_3_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, new_AGEMA_signal_8843, mcs1_mcs_mat1_3_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_8848, new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_3_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_9676, new_AGEMA_signal_9675, new_AGEMA_signal_9674, mcs1_mcs_mat1_3_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({new_AGEMA_signal_8848, new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_3_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_13441, new_AGEMA_signal_13440, new_AGEMA_signal_13439, mcs1_mcs_mat1_3_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_14878, new_AGEMA_signal_14877, new_AGEMA_signal_14876, mcs1_mcs_mat1_3_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({new_AGEMA_signal_13441, new_AGEMA_signal_13440, new_AGEMA_signal_13439, mcs1_mcs_mat1_3_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, new_AGEMA_signal_8849, mcs1_mcs_mat1_3_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_8854, new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_3_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .c ({new_AGEMA_signal_12007, new_AGEMA_signal_12006, new_AGEMA_signal_12005, mcs1_mcs_mat1_3_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({new_AGEMA_signal_8854, new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_3_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_14902, new_AGEMA_signal_14901, new_AGEMA_signal_14900, mcs1_mcs_mat1_3_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, new_AGEMA_signal_8855, mcs1_mcs_mat1_3_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_16114, new_AGEMA_signal_16113, new_AGEMA_signal_16112, mcs1_mcs_mat1_3_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_13459, new_AGEMA_signal_13458, new_AGEMA_signal_13457, mcs1_mcs_mat1_3_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_14902, new_AGEMA_signal_14901, new_AGEMA_signal_14900, mcs1_mcs_mat1_3_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_12013, new_AGEMA_signal_12012, new_AGEMA_signal_12011, mcs1_mcs_mat1_3_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_13459, new_AGEMA_signal_13458, new_AGEMA_signal_13457, mcs1_mcs_mat1_3_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_12013, new_AGEMA_signal_12012, new_AGEMA_signal_12011, mcs1_mcs_mat1_3_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({new_AGEMA_signal_8857, new_AGEMA_signal_8856, new_AGEMA_signal_8855, mcs1_mcs_mat1_3_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_17683, new_AGEMA_signal_17682, new_AGEMA_signal_17681, mcs1_mcs_mat1_3_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_14905, new_AGEMA_signal_14904, new_AGEMA_signal_14903, mcs1_mcs_mat1_3_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_18361, new_AGEMA_signal_18360, new_AGEMA_signal_18359, mcs1_mcs_mat1_3_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_13462, new_AGEMA_signal_13461, new_AGEMA_signal_13460, mcs1_mcs_mat1_3_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .c ({new_AGEMA_signal_14905, new_AGEMA_signal_14904, new_AGEMA_signal_14903, mcs1_mcs_mat1_3_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .c ({new_AGEMA_signal_14908, new_AGEMA_signal_14907, new_AGEMA_signal_14906, mcs1_mcs_mat1_3_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .c ({new_AGEMA_signal_17683, new_AGEMA_signal_17682, new_AGEMA_signal_17681, mcs1_mcs_mat1_3_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_13462, new_AGEMA_signal_13461, new_AGEMA_signal_13460, mcs1_mcs_mat1_3_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_17686, new_AGEMA_signal_17685, new_AGEMA_signal_17684, mcs1_mcs_mat1_3_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({new_AGEMA_signal_13462, new_AGEMA_signal_13461, new_AGEMA_signal_13460, mcs1_mcs_mat1_3_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .b ({new_AGEMA_signal_8860, new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_3_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_12025, new_AGEMA_signal_12024, new_AGEMA_signal_12023, mcs1_mcs_mat1_3_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({new_AGEMA_signal_8860, new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_3_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({new_AGEMA_signal_12031, new_AGEMA_signal_12030, new_AGEMA_signal_12029, mcs1_mcs_mat1_3_mcs_out[51]}), .c ({new_AGEMA_signal_13471, new_AGEMA_signal_13470, new_AGEMA_signal_13469, mcs1_mcs_mat1_3_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .c ({new_AGEMA_signal_12031, new_AGEMA_signal_12030, new_AGEMA_signal_12029, mcs1_mcs_mat1_3_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, new_AGEMA_signal_8861, mcs1_mcs_mat1_3_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_10870, new_AGEMA_signal_10869, new_AGEMA_signal_10868, mcs1_mcs_mat1_3_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, new_AGEMA_signal_8861, mcs1_mcs_mat1_3_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_17692, new_AGEMA_signal_17691, new_AGEMA_signal_17690, mcs1_mcs_mat1_3_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_18373, new_AGEMA_signal_18372, new_AGEMA_signal_18371, mcs1_mcs_mat1_3_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .b ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_17692, new_AGEMA_signal_17691, new_AGEMA_signal_17690, mcs1_mcs_mat1_3_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_16987, new_AGEMA_signal_16986, new_AGEMA_signal_16985, mcs1_mcs_mat1_3_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_17695, new_AGEMA_signal_17694, new_AGEMA_signal_17693, mcs1_mcs_mat1_3_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .c ({new_AGEMA_signal_16987, new_AGEMA_signal_16986, new_AGEMA_signal_16985, mcs1_mcs_mat1_3_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({new_AGEMA_signal_13477, new_AGEMA_signal_13476, new_AGEMA_signal_13475, mcs1_mcs_mat1_3_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({new_AGEMA_signal_8866, new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_3_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_10876, new_AGEMA_signal_10875, new_AGEMA_signal_10874, mcs1_mcs_mat1_3_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .b ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_12043, new_AGEMA_signal_12042, new_AGEMA_signal_12041, mcs1_mcs_mat1_3_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({new_AGEMA_signal_8866, new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_3_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_14932, new_AGEMA_signal_14931, new_AGEMA_signal_14930, mcs1_mcs_mat1_3_mcs_out[35]}), .b ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_16132, new_AGEMA_signal_16131, new_AGEMA_signal_16130, mcs1_mcs_mat1_3_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_13489, new_AGEMA_signal_13488, new_AGEMA_signal_13487, mcs1_mcs_mat1_3_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, new_AGEMA_signal_8867, mcs1_mcs_mat1_3_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_14932, new_AGEMA_signal_14931, new_AGEMA_signal_14930, mcs1_mcs_mat1_3_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_12049, new_AGEMA_signal_12048, new_AGEMA_signal_12047, mcs1_mcs_mat1_3_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .c ({new_AGEMA_signal_13489, new_AGEMA_signal_13488, new_AGEMA_signal_13487, mcs1_mcs_mat1_3_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .c ({new_AGEMA_signal_12049, new_AGEMA_signal_12048, new_AGEMA_signal_12047, mcs1_mcs_mat1_3_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({new_AGEMA_signal_8869, new_AGEMA_signal_8868, new_AGEMA_signal_8867, mcs1_mcs_mat1_3_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_8872, new_AGEMA_signal_8871, new_AGEMA_signal_8870, mcs1_mcs_mat1_3_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_9703, new_AGEMA_signal_9702, new_AGEMA_signal_9701, mcs1_mcs_mat1_3_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({new_AGEMA_signal_12055, new_AGEMA_signal_12054, new_AGEMA_signal_12053, mcs1_mcs_mat1_3_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_13495, new_AGEMA_signal_13494, new_AGEMA_signal_13493, mcs1_mcs_mat1_3_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_8872, new_AGEMA_signal_8871, new_AGEMA_signal_8870, mcs1_mcs_mat1_3_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_12055, new_AGEMA_signal_12054, new_AGEMA_signal_12053, mcs1_mcs_mat1_3_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({new_AGEMA_signal_8872, new_AGEMA_signal_8871, new_AGEMA_signal_8870, mcs1_mcs_mat1_3_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({new_AGEMA_signal_13501, new_AGEMA_signal_13500, new_AGEMA_signal_13499, mcs1_mcs_mat1_3_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, new_AGEMA_signal_8873, mcs1_mcs_mat1_3_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_10894, new_AGEMA_signal_10893, new_AGEMA_signal_10892, mcs1_mcs_mat1_3_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_12073, new_AGEMA_signal_12072, new_AGEMA_signal_12071, mcs1_mcs_mat1_3_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_10894, new_AGEMA_signal_10893, new_AGEMA_signal_10892, mcs1_mcs_mat1_3_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .c ({new_AGEMA_signal_12079, new_AGEMA_signal_12078, new_AGEMA_signal_12077, mcs1_mcs_mat1_3_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({new_AGEMA_signal_8878, new_AGEMA_signal_8877, new_AGEMA_signal_8876, mcs1_mcs_mat1_3_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, new_AGEMA_signal_8879, mcs1_mcs_mat1_3_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({new_AGEMA_signal_13531, new_AGEMA_signal_13530, new_AGEMA_signal_13529, mcs1_mcs_mat1_3_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_8884, new_AGEMA_signal_8883, new_AGEMA_signal_8882, mcs1_mcs_mat1_3_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_10903, new_AGEMA_signal_10902, new_AGEMA_signal_10901, mcs1_mcs_mat1_3_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_8884, new_AGEMA_signal_8883, new_AGEMA_signal_8882, mcs1_mcs_mat1_3_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_9718, new_AGEMA_signal_9717, new_AGEMA_signal_9716, mcs1_mcs_mat1_3_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({new_AGEMA_signal_8884, new_AGEMA_signal_8883, new_AGEMA_signal_8882, mcs1_mcs_mat1_3_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_12097, new_AGEMA_signal_12096, new_AGEMA_signal_12095, mcs1_mcs_mat1_3_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, new_AGEMA_signal_8885, mcs1_mcs_mat1_3_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_13537, new_AGEMA_signal_13536, new_AGEMA_signal_13535, mcs1_mcs_mat1_3_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_12097, new_AGEMA_signal_12096, new_AGEMA_signal_12095, mcs1_mcs_mat1_3_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .c ({new_AGEMA_signal_13543, new_AGEMA_signal_13542, new_AGEMA_signal_13541, mcs1_mcs_mat1_3_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_10909, new_AGEMA_signal_10908, new_AGEMA_signal_10907, mcs1_mcs_mat1_3_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_12097, new_AGEMA_signal_12096, new_AGEMA_signal_12095, mcs1_mcs_mat1_3_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_10909, new_AGEMA_signal_10908, new_AGEMA_signal_10907, mcs1_mcs_mat1_3_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .c ({new_AGEMA_signal_12100, new_AGEMA_signal_12099, new_AGEMA_signal_12098, mcs1_mcs_mat1_3_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, new_AGEMA_signal_8885, mcs1_mcs_mat1_3_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U44 ( .a ({new_AGEMA_signal_10954, new_AGEMA_signal_10953, new_AGEMA_signal_10952, mcs1_mcs_mat1_4_mcs_out[90]}), .b ({new_AGEMA_signal_17752, new_AGEMA_signal_17751, new_AGEMA_signal_17750, mcs1_mcs_mat1_4_mcs_out[94]}), .c ({new_AGEMA_signal_18406, new_AGEMA_signal_18405, new_AGEMA_signal_18404, mcs1_mcs_mat1_4_n93}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .c ({new_AGEMA_signal_17059, new_AGEMA_signal_17058, new_AGEMA_signal_17057, mcs1_mcs_mat1_4_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .b ({new_AGEMA_signal_8890, new_AGEMA_signal_8889, new_AGEMA_signal_8888, mcs1_mcs_mat1_4_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_9727, new_AGEMA_signal_9726, new_AGEMA_signal_9725, mcs1_mcs_mat1_4_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({new_AGEMA_signal_8890, new_AGEMA_signal_8889, new_AGEMA_signal_8888, mcs1_mcs_mat1_4_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_10921, new_AGEMA_signal_10920, new_AGEMA_signal_10919, mcs1_mcs_mat1_4_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_12112, new_AGEMA_signal_12111, new_AGEMA_signal_12110, mcs1_mcs_mat1_4_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_8893, new_AGEMA_signal_8892, new_AGEMA_signal_8891, mcs1_mcs_mat1_4_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_10921, new_AGEMA_signal_10920, new_AGEMA_signal_10919, mcs1_mcs_mat1_4_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({new_AGEMA_signal_8893, new_AGEMA_signal_8892, new_AGEMA_signal_8891, mcs1_mcs_mat1_4_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_8896, new_AGEMA_signal_8895, new_AGEMA_signal_8894, mcs1_mcs_mat1_4_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_12124, new_AGEMA_signal_12123, new_AGEMA_signal_12122, mcs1_mcs_mat1_4_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_13561, new_AGEMA_signal_13560, new_AGEMA_signal_13559, mcs1_mcs_mat1_4_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_9736, new_AGEMA_signal_9735, new_AGEMA_signal_9734, mcs1_mcs_mat1_4_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_10930, new_AGEMA_signal_10929, new_AGEMA_signal_10928, mcs1_mcs_mat1_4_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .c ({new_AGEMA_signal_9736, new_AGEMA_signal_9735, new_AGEMA_signal_9734, mcs1_mcs_mat1_4_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_12124, new_AGEMA_signal_12123, new_AGEMA_signal_12122, mcs1_mcs_mat1_4_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({new_AGEMA_signal_8896, new_AGEMA_signal_8895, new_AGEMA_signal_8894, mcs1_mcs_mat1_4_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_17743, new_AGEMA_signal_17742, new_AGEMA_signal_17741, mcs1_mcs_mat1_4_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_18421, new_AGEMA_signal_18420, new_AGEMA_signal_18419, mcs1_mcs_mat1_4_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_13570, new_AGEMA_signal_13569, new_AGEMA_signal_13568, mcs1_mcs_mat1_4_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_17743, new_AGEMA_signal_17742, new_AGEMA_signal_17741, mcs1_mcs_mat1_4_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({new_AGEMA_signal_13570, new_AGEMA_signal_13569, new_AGEMA_signal_13568, mcs1_mcs_mat1_4_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({new_AGEMA_signal_8899, new_AGEMA_signal_8898, new_AGEMA_signal_8897, mcs1_mcs_mat1_4_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({new_AGEMA_signal_10942, new_AGEMA_signal_10941, new_AGEMA_signal_10940, mcs1_mcs_mat1_4_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_12136, new_AGEMA_signal_12135, new_AGEMA_signal_12134, mcs1_mcs_mat1_4_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_8902, new_AGEMA_signal_8901, new_AGEMA_signal_8900, mcs1_mcs_mat1_4_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_10942, new_AGEMA_signal_10941, new_AGEMA_signal_10940, mcs1_mcs_mat1_4_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .b ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .c ({new_AGEMA_signal_12139, new_AGEMA_signal_12138, new_AGEMA_signal_12137, mcs1_mcs_mat1_4_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({new_AGEMA_signal_8902, new_AGEMA_signal_8901, new_AGEMA_signal_8900, mcs1_mcs_mat1_4_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_8905, new_AGEMA_signal_8904, new_AGEMA_signal_8903, mcs1_mcs_mat1_4_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_10948, new_AGEMA_signal_10947, new_AGEMA_signal_10946, mcs1_mcs_mat1_4_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_8905, new_AGEMA_signal_8904, new_AGEMA_signal_8903, mcs1_mcs_mat1_4_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .c ({new_AGEMA_signal_9748, new_AGEMA_signal_9747, new_AGEMA_signal_9746, mcs1_mcs_mat1_4_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({new_AGEMA_signal_8905, new_AGEMA_signal_8904, new_AGEMA_signal_8903, mcs1_mcs_mat1_4_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_17068, new_AGEMA_signal_17067, new_AGEMA_signal_17066, mcs1_mcs_mat1_4_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .c ({new_AGEMA_signal_17752, new_AGEMA_signal_17751, new_AGEMA_signal_17750, mcs1_mcs_mat1_4_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_13591, new_AGEMA_signal_13590, new_AGEMA_signal_13589, mcs1_mcs_mat1_4_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_17068, new_AGEMA_signal_17067, new_AGEMA_signal_17066, mcs1_mcs_mat1_4_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_17071, new_AGEMA_signal_17070, new_AGEMA_signal_17069, mcs1_mcs_mat1_4_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({new_AGEMA_signal_13591, new_AGEMA_signal_13590, new_AGEMA_signal_13589, mcs1_mcs_mat1_4_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .b ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .c ({new_AGEMA_signal_10954, new_AGEMA_signal_10953, new_AGEMA_signal_10952, mcs1_mcs_mat1_4_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .b ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_10957, new_AGEMA_signal_10956, new_AGEMA_signal_10955, mcs1_mcs_mat1_4_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({new_AGEMA_signal_12151, new_AGEMA_signal_12150, new_AGEMA_signal_12149, mcs1_mcs_mat1_4_mcs_out[87]}), .c ({new_AGEMA_signal_13594, new_AGEMA_signal_13593, new_AGEMA_signal_13592, mcs1_mcs_mat1_4_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .c ({new_AGEMA_signal_12151, new_AGEMA_signal_12150, new_AGEMA_signal_12149, mcs1_mcs_mat1_4_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .c ({new_AGEMA_signal_12160, new_AGEMA_signal_12159, new_AGEMA_signal_12158, mcs1_mcs_mat1_4_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({new_AGEMA_signal_8908, new_AGEMA_signal_8907, new_AGEMA_signal_8906, mcs1_mcs_mat1_4_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_13609, new_AGEMA_signal_13608, new_AGEMA_signal_13607, mcs1_mcs_mat1_4_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_15058, new_AGEMA_signal_15057, new_AGEMA_signal_15056, mcs1_mcs_mat1_4_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({new_AGEMA_signal_13609, new_AGEMA_signal_13608, new_AGEMA_signal_13607, mcs1_mcs_mat1_4_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_8911, new_AGEMA_signal_8910, new_AGEMA_signal_8909, mcs1_mcs_mat1_4_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_9757, new_AGEMA_signal_9756, new_AGEMA_signal_9755, mcs1_mcs_mat1_4_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({new_AGEMA_signal_8911, new_AGEMA_signal_8910, new_AGEMA_signal_8909, mcs1_mcs_mat1_4_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({new_AGEMA_signal_8914, new_AGEMA_signal_8913, new_AGEMA_signal_8912, mcs1_mcs_mat1_4_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_8917, new_AGEMA_signal_8916, new_AGEMA_signal_8915, mcs1_mcs_mat1_4_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .c ({new_AGEMA_signal_12184, new_AGEMA_signal_12183, new_AGEMA_signal_12182, mcs1_mcs_mat1_4_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({new_AGEMA_signal_8917, new_AGEMA_signal_8916, new_AGEMA_signal_8915, mcs1_mcs_mat1_4_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_19087, new_AGEMA_signal_19086, new_AGEMA_signal_19085, mcs1_mcs_mat1_4_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_13627, new_AGEMA_signal_13626, new_AGEMA_signal_13625, mcs1_mcs_mat1_4_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_19807, new_AGEMA_signal_19806, new_AGEMA_signal_19805, mcs1_mcs_mat1_4_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_18439, new_AGEMA_signal_18438, new_AGEMA_signal_18437, mcs1_mcs_mat1_4_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_19087, new_AGEMA_signal_19086, new_AGEMA_signal_19085, mcs1_mcs_mat1_4_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_17767, new_AGEMA_signal_17766, new_AGEMA_signal_17765, mcs1_mcs_mat1_4_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_18439, new_AGEMA_signal_18438, new_AGEMA_signal_18437, mcs1_mcs_mat1_4_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_17767, new_AGEMA_signal_17766, new_AGEMA_signal_17765, mcs1_mcs_mat1_4_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({new_AGEMA_signal_13627, new_AGEMA_signal_13626, new_AGEMA_signal_13625, mcs1_mcs_mat1_4_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_12193, new_AGEMA_signal_12192, new_AGEMA_signal_12191, mcs1_mcs_mat1_4_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_9769, new_AGEMA_signal_9768, new_AGEMA_signal_9767, mcs1_mcs_mat1_4_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_13630, new_AGEMA_signal_13629, new_AGEMA_signal_13628, mcs1_mcs_mat1_4_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_8920, new_AGEMA_signal_8919, new_AGEMA_signal_8918, mcs1_mcs_mat1_4_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .c ({new_AGEMA_signal_9769, new_AGEMA_signal_9768, new_AGEMA_signal_9767, mcs1_mcs_mat1_4_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .c ({new_AGEMA_signal_9772, new_AGEMA_signal_9771, new_AGEMA_signal_9770, mcs1_mcs_mat1_4_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .c ({new_AGEMA_signal_12193, new_AGEMA_signal_12192, new_AGEMA_signal_12191, mcs1_mcs_mat1_4_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_8920, new_AGEMA_signal_8919, new_AGEMA_signal_8918, mcs1_mcs_mat1_4_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_12196, new_AGEMA_signal_12195, new_AGEMA_signal_12194, mcs1_mcs_mat1_4_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({new_AGEMA_signal_8920, new_AGEMA_signal_8919, new_AGEMA_signal_8918, mcs1_mcs_mat1_4_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .b ({new_AGEMA_signal_8923, new_AGEMA_signal_8922, new_AGEMA_signal_8921, mcs1_mcs_mat1_4_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_12208, new_AGEMA_signal_12207, new_AGEMA_signal_12206, mcs1_mcs_mat1_4_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({new_AGEMA_signal_8923, new_AGEMA_signal_8922, new_AGEMA_signal_8921, mcs1_mcs_mat1_4_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({new_AGEMA_signal_12214, new_AGEMA_signal_12213, new_AGEMA_signal_12212, mcs1_mcs_mat1_4_mcs_out[51]}), .c ({new_AGEMA_signal_13645, new_AGEMA_signal_13644, new_AGEMA_signal_13643, mcs1_mcs_mat1_4_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .c ({new_AGEMA_signal_12214, new_AGEMA_signal_12213, new_AGEMA_signal_12212, mcs1_mcs_mat1_4_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_13648, new_AGEMA_signal_13647, new_AGEMA_signal_13646, mcs1_mcs_mat1_4_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_17086, new_AGEMA_signal_17085, new_AGEMA_signal_17084, mcs1_mcs_mat1_4_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({new_AGEMA_signal_13648, new_AGEMA_signal_13647, new_AGEMA_signal_13646, mcs1_mcs_mat1_4_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_12217, new_AGEMA_signal_12216, new_AGEMA_signal_12215, mcs1_mcs_mat1_4_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_13654, new_AGEMA_signal_13653, new_AGEMA_signal_13652, mcs1_mcs_mat1_4_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_12217, new_AGEMA_signal_12216, new_AGEMA_signal_12215, mcs1_mcs_mat1_4_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_10981, new_AGEMA_signal_10980, new_AGEMA_signal_10979, mcs1_mcs_mat1_4_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_12220, new_AGEMA_signal_12219, new_AGEMA_signal_12218, mcs1_mcs_mat1_4_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .c ({new_AGEMA_signal_10981, new_AGEMA_signal_10980, new_AGEMA_signal_10979, mcs1_mcs_mat1_4_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({new_AGEMA_signal_8926, new_AGEMA_signal_8925, new_AGEMA_signal_8924, mcs1_mcs_mat1_4_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({new_AGEMA_signal_8929, new_AGEMA_signal_8928, new_AGEMA_signal_8927, mcs1_mcs_mat1_4_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_10987, new_AGEMA_signal_10986, new_AGEMA_signal_10985, mcs1_mcs_mat1_4_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_12229, new_AGEMA_signal_12228, new_AGEMA_signal_12227, mcs1_mcs_mat1_4_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({new_AGEMA_signal_8929, new_AGEMA_signal_8928, new_AGEMA_signal_8927, mcs1_mcs_mat1_4_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_15115, new_AGEMA_signal_15114, new_AGEMA_signal_15113, mcs1_mcs_mat1_4_mcs_out[35]}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_16234, new_AGEMA_signal_16233, new_AGEMA_signal_16232, mcs1_mcs_mat1_4_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_13672, new_AGEMA_signal_13671, new_AGEMA_signal_13670, mcs1_mcs_mat1_4_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_8932, new_AGEMA_signal_8931, new_AGEMA_signal_8930, mcs1_mcs_mat1_4_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_15115, new_AGEMA_signal_15114, new_AGEMA_signal_15113, mcs1_mcs_mat1_4_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_12235, new_AGEMA_signal_12234, new_AGEMA_signal_12233, mcs1_mcs_mat1_4_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .c ({new_AGEMA_signal_13672, new_AGEMA_signal_13671, new_AGEMA_signal_13670, mcs1_mcs_mat1_4_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .c ({new_AGEMA_signal_12235, new_AGEMA_signal_12234, new_AGEMA_signal_12233, mcs1_mcs_mat1_4_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({new_AGEMA_signal_8932, new_AGEMA_signal_8931, new_AGEMA_signal_8930, mcs1_mcs_mat1_4_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_13675, new_AGEMA_signal_13674, new_AGEMA_signal_13673, mcs1_mcs_mat1_4_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_15118, new_AGEMA_signal_15117, new_AGEMA_signal_15116, mcs1_mcs_mat1_4_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({new_AGEMA_signal_17779, new_AGEMA_signal_17778, new_AGEMA_signal_17777, mcs1_mcs_mat1_4_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_18448, new_AGEMA_signal_18447, new_AGEMA_signal_18446, mcs1_mcs_mat1_4_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_13675, new_AGEMA_signal_13674, new_AGEMA_signal_13673, mcs1_mcs_mat1_4_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_17779, new_AGEMA_signal_17778, new_AGEMA_signal_17777, mcs1_mcs_mat1_4_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({new_AGEMA_signal_13675, new_AGEMA_signal_13674, new_AGEMA_signal_13673, mcs1_mcs_mat1_4_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({new_AGEMA_signal_8935, new_AGEMA_signal_8934, new_AGEMA_signal_8933, mcs1_mcs_mat1_4_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({new_AGEMA_signal_8938, new_AGEMA_signal_8937, new_AGEMA_signal_8936, mcs1_mcs_mat1_4_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_11005, new_AGEMA_signal_11004, new_AGEMA_signal_11003, mcs1_mcs_mat1_4_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_12259, new_AGEMA_signal_12258, new_AGEMA_signal_12257, mcs1_mcs_mat1_4_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_11005, new_AGEMA_signal_11004, new_AGEMA_signal_11003, mcs1_mcs_mat1_4_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .c ({new_AGEMA_signal_12265, new_AGEMA_signal_12264, new_AGEMA_signal_12263, mcs1_mcs_mat1_4_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({new_AGEMA_signal_8941, new_AGEMA_signal_8940, new_AGEMA_signal_8939, mcs1_mcs_mat1_4_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({new_AGEMA_signal_13705, new_AGEMA_signal_13704, new_AGEMA_signal_13703, mcs1_mcs_mat1_4_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({new_AGEMA_signal_8944, new_AGEMA_signal_8943, new_AGEMA_signal_8942, mcs1_mcs_mat1_4_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_8947, new_AGEMA_signal_8946, new_AGEMA_signal_8945, mcs1_mcs_mat1_4_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_11017, new_AGEMA_signal_11016, new_AGEMA_signal_11015, mcs1_mcs_mat1_4_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_8947, new_AGEMA_signal_8946, new_AGEMA_signal_8945, mcs1_mcs_mat1_4_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_9802, new_AGEMA_signal_9801, new_AGEMA_signal_9800, mcs1_mcs_mat1_4_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({new_AGEMA_signal_8947, new_AGEMA_signal_8946, new_AGEMA_signal_8945, mcs1_mcs_mat1_4_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_12283, new_AGEMA_signal_12282, new_AGEMA_signal_12281, mcs1_mcs_mat1_4_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_8950, new_AGEMA_signal_8949, new_AGEMA_signal_8948, mcs1_mcs_mat1_4_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_13717, new_AGEMA_signal_13716, new_AGEMA_signal_13715, mcs1_mcs_mat1_4_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_12283, new_AGEMA_signal_12282, new_AGEMA_signal_12281, mcs1_mcs_mat1_4_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .c ({new_AGEMA_signal_13723, new_AGEMA_signal_13722, new_AGEMA_signal_13721, mcs1_mcs_mat1_4_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_11023, new_AGEMA_signal_11022, new_AGEMA_signal_11021, mcs1_mcs_mat1_4_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_12283, new_AGEMA_signal_12282, new_AGEMA_signal_12281, mcs1_mcs_mat1_4_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_11023, new_AGEMA_signal_11022, new_AGEMA_signal_11021, mcs1_mcs_mat1_4_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .c ({new_AGEMA_signal_12286, new_AGEMA_signal_12285, new_AGEMA_signal_12284, mcs1_mcs_mat1_4_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({new_AGEMA_signal_8950, new_AGEMA_signal_8949, new_AGEMA_signal_8948, mcs1_mcs_mat1_4_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U44 ( .a ({new_AGEMA_signal_11071, new_AGEMA_signal_11070, new_AGEMA_signal_11069, mcs1_mcs_mat1_5_mcs_out[90]}), .b ({new_AGEMA_signal_12331, new_AGEMA_signal_12330, new_AGEMA_signal_12329, mcs1_mcs_mat1_5_mcs_out[94]}), .c ({new_AGEMA_signal_13732, new_AGEMA_signal_13731, new_AGEMA_signal_13730, mcs1_mcs_mat1_5_n93}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .c ({new_AGEMA_signal_11029, new_AGEMA_signal_11028, new_AGEMA_signal_11027, mcs1_mcs_mat1_5_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .b ({new_AGEMA_signal_8953, new_AGEMA_signal_8952, new_AGEMA_signal_8951, mcs1_mcs_mat1_5_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_9811, new_AGEMA_signal_9810, new_AGEMA_signal_9809, mcs1_mcs_mat1_5_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({new_AGEMA_signal_8953, new_AGEMA_signal_8952, new_AGEMA_signal_8951, mcs1_mcs_mat1_5_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_11038, new_AGEMA_signal_11037, new_AGEMA_signal_11036, mcs1_mcs_mat1_5_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_12298, new_AGEMA_signal_12297, new_AGEMA_signal_12296, mcs1_mcs_mat1_5_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_8956, new_AGEMA_signal_8955, new_AGEMA_signal_8954, mcs1_mcs_mat1_5_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_11038, new_AGEMA_signal_11037, new_AGEMA_signal_11036, mcs1_mcs_mat1_5_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({new_AGEMA_signal_8956, new_AGEMA_signal_8955, new_AGEMA_signal_8954, mcs1_mcs_mat1_5_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_13750, new_AGEMA_signal_13749, new_AGEMA_signal_13748, mcs1_mcs_mat1_5_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_17815, new_AGEMA_signal_17814, new_AGEMA_signal_17813, mcs1_mcs_mat1_5_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_18478, new_AGEMA_signal_18477, new_AGEMA_signal_18476, mcs1_mcs_mat1_5_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_15190, new_AGEMA_signal_15189, new_AGEMA_signal_15188, mcs1_mcs_mat1_5_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_17146, new_AGEMA_signal_17145, new_AGEMA_signal_17144, mcs1_mcs_mat1_5_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .c ({new_AGEMA_signal_15190, new_AGEMA_signal_15189, new_AGEMA_signal_15188, mcs1_mcs_mat1_5_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .b ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_17815, new_AGEMA_signal_17814, new_AGEMA_signal_17813, mcs1_mcs_mat1_5_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({new_AGEMA_signal_13750, new_AGEMA_signal_13749, new_AGEMA_signal_13748, mcs1_mcs_mat1_5_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_12307, new_AGEMA_signal_12306, new_AGEMA_signal_12305, mcs1_mcs_mat1_5_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_13753, new_AGEMA_signal_13752, new_AGEMA_signal_13751, mcs1_mcs_mat1_5_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_8959, new_AGEMA_signal_8958, new_AGEMA_signal_8957, mcs1_mcs_mat1_5_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_12307, new_AGEMA_signal_12306, new_AGEMA_signal_12305, mcs1_mcs_mat1_5_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({new_AGEMA_signal_8959, new_AGEMA_signal_8958, new_AGEMA_signal_8957, mcs1_mcs_mat1_5_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({new_AGEMA_signal_8962, new_AGEMA_signal_8961, new_AGEMA_signal_8960, mcs1_mcs_mat1_5_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({new_AGEMA_signal_11056, new_AGEMA_signal_11055, new_AGEMA_signal_11054, mcs1_mcs_mat1_5_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_12319, new_AGEMA_signal_12318, new_AGEMA_signal_12317, mcs1_mcs_mat1_5_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_8965, new_AGEMA_signal_8964, new_AGEMA_signal_8963, mcs1_mcs_mat1_5_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_11056, new_AGEMA_signal_11055, new_AGEMA_signal_11054, mcs1_mcs_mat1_5_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .b ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .c ({new_AGEMA_signal_12322, new_AGEMA_signal_12321, new_AGEMA_signal_12320, mcs1_mcs_mat1_5_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({new_AGEMA_signal_8965, new_AGEMA_signal_8964, new_AGEMA_signal_8963, mcs1_mcs_mat1_5_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_13774, new_AGEMA_signal_13773, new_AGEMA_signal_13772, mcs1_mcs_mat1_5_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_17152, new_AGEMA_signal_17151, new_AGEMA_signal_17150, mcs1_mcs_mat1_5_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_13774, new_AGEMA_signal_13773, new_AGEMA_signal_13772, mcs1_mcs_mat1_5_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .c ({new_AGEMA_signal_15220, new_AGEMA_signal_15219, new_AGEMA_signal_15218, mcs1_mcs_mat1_5_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({new_AGEMA_signal_13774, new_AGEMA_signal_13773, new_AGEMA_signal_13772, mcs1_mcs_mat1_5_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_11062, new_AGEMA_signal_11061, new_AGEMA_signal_11060, mcs1_mcs_mat1_5_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .c ({new_AGEMA_signal_12331, new_AGEMA_signal_12330, new_AGEMA_signal_12329, mcs1_mcs_mat1_5_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_8968, new_AGEMA_signal_8967, new_AGEMA_signal_8966, mcs1_mcs_mat1_5_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_11062, new_AGEMA_signal_11061, new_AGEMA_signal_11060, mcs1_mcs_mat1_5_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_11065, new_AGEMA_signal_11064, new_AGEMA_signal_11063, mcs1_mcs_mat1_5_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({new_AGEMA_signal_8968, new_AGEMA_signal_8967, new_AGEMA_signal_8966, mcs1_mcs_mat1_5_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .b ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .c ({new_AGEMA_signal_11071, new_AGEMA_signal_11070, new_AGEMA_signal_11069, mcs1_mcs_mat1_5_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .b ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_11074, new_AGEMA_signal_11073, new_AGEMA_signal_11072, mcs1_mcs_mat1_5_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({new_AGEMA_signal_12340, new_AGEMA_signal_12339, new_AGEMA_signal_12338, mcs1_mcs_mat1_5_mcs_out[87]}), .c ({new_AGEMA_signal_13780, new_AGEMA_signal_13779, new_AGEMA_signal_13778, mcs1_mcs_mat1_5_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .c ({new_AGEMA_signal_12340, new_AGEMA_signal_12339, new_AGEMA_signal_12338, mcs1_mcs_mat1_5_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .c ({new_AGEMA_signal_17830, new_AGEMA_signal_17829, new_AGEMA_signal_17828, mcs1_mcs_mat1_5_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({new_AGEMA_signal_13783, new_AGEMA_signal_13782, new_AGEMA_signal_13781, mcs1_mcs_mat1_5_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_8971, new_AGEMA_signal_8970, new_AGEMA_signal_8969, mcs1_mcs_mat1_5_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_9832, new_AGEMA_signal_9831, new_AGEMA_signal_9830, mcs1_mcs_mat1_5_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({new_AGEMA_signal_8971, new_AGEMA_signal_8970, new_AGEMA_signal_8969, mcs1_mcs_mat1_5_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_8974, new_AGEMA_signal_8973, new_AGEMA_signal_8972, mcs1_mcs_mat1_5_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_9838, new_AGEMA_signal_9837, new_AGEMA_signal_9836, mcs1_mcs_mat1_5_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({new_AGEMA_signal_8974, new_AGEMA_signal_8973, new_AGEMA_signal_8972, mcs1_mcs_mat1_5_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({new_AGEMA_signal_8977, new_AGEMA_signal_8976, new_AGEMA_signal_8975, mcs1_mcs_mat1_5_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_13801, new_AGEMA_signal_13800, new_AGEMA_signal_13799, mcs1_mcs_mat1_5_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .c ({new_AGEMA_signal_17836, new_AGEMA_signal_17835, new_AGEMA_signal_17834, mcs1_mcs_mat1_5_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({new_AGEMA_signal_13801, new_AGEMA_signal_13800, new_AGEMA_signal_13799, mcs1_mcs_mat1_5_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_15262, new_AGEMA_signal_15261, new_AGEMA_signal_15260, mcs1_mcs_mat1_5_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_8980, new_AGEMA_signal_8979, new_AGEMA_signal_8978, mcs1_mcs_mat1_5_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_16336, new_AGEMA_signal_16335, new_AGEMA_signal_16334, mcs1_mcs_mat1_5_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_13810, new_AGEMA_signal_13809, new_AGEMA_signal_13808, mcs1_mcs_mat1_5_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_15262, new_AGEMA_signal_15261, new_AGEMA_signal_15260, mcs1_mcs_mat1_5_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_12367, new_AGEMA_signal_12366, new_AGEMA_signal_12365, mcs1_mcs_mat1_5_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_13810, new_AGEMA_signal_13809, new_AGEMA_signal_13808, mcs1_mcs_mat1_5_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_12367, new_AGEMA_signal_12366, new_AGEMA_signal_12365, mcs1_mcs_mat1_5_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({new_AGEMA_signal_8980, new_AGEMA_signal_8979, new_AGEMA_signal_8978, mcs1_mcs_mat1_5_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_12376, new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_5_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_9850, new_AGEMA_signal_9849, new_AGEMA_signal_9848, mcs1_mcs_mat1_5_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_13813, new_AGEMA_signal_13812, new_AGEMA_signal_13811, mcs1_mcs_mat1_5_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_8983, new_AGEMA_signal_8982, new_AGEMA_signal_8981, mcs1_mcs_mat1_5_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .c ({new_AGEMA_signal_9850, new_AGEMA_signal_9849, new_AGEMA_signal_9848, mcs1_mcs_mat1_5_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .c ({new_AGEMA_signal_9853, new_AGEMA_signal_9852, new_AGEMA_signal_9851, mcs1_mcs_mat1_5_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .c ({new_AGEMA_signal_12376, new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_5_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_8983, new_AGEMA_signal_8982, new_AGEMA_signal_8981, mcs1_mcs_mat1_5_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, new_AGEMA_signal_12377, mcs1_mcs_mat1_5_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({new_AGEMA_signal_8983, new_AGEMA_signal_8982, new_AGEMA_signal_8981, mcs1_mcs_mat1_5_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .b ({new_AGEMA_signal_8986, new_AGEMA_signal_8985, new_AGEMA_signal_8984, mcs1_mcs_mat1_5_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_12391, new_AGEMA_signal_12390, new_AGEMA_signal_12389, mcs1_mcs_mat1_5_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({new_AGEMA_signal_8986, new_AGEMA_signal_8985, new_AGEMA_signal_8984, mcs1_mcs_mat1_5_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({new_AGEMA_signal_17842, new_AGEMA_signal_17841, new_AGEMA_signal_17840, mcs1_mcs_mat1_5_mcs_out[51]}), .c ({new_AGEMA_signal_18505, new_AGEMA_signal_18504, new_AGEMA_signal_18503, mcs1_mcs_mat1_5_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .c ({new_AGEMA_signal_17842, new_AGEMA_signal_17841, new_AGEMA_signal_17840, mcs1_mcs_mat1_5_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_8989, new_AGEMA_signal_8988, new_AGEMA_signal_8987, mcs1_mcs_mat1_5_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_11098, new_AGEMA_signal_11097, new_AGEMA_signal_11096, mcs1_mcs_mat1_5_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({new_AGEMA_signal_8989, new_AGEMA_signal_8988, new_AGEMA_signal_8987, mcs1_mcs_mat1_5_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_12403, new_AGEMA_signal_12402, new_AGEMA_signal_12401, mcs1_mcs_mat1_5_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_13834, new_AGEMA_signal_13833, new_AGEMA_signal_13832, mcs1_mcs_mat1_5_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .b ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_12403, new_AGEMA_signal_12402, new_AGEMA_signal_12401, mcs1_mcs_mat1_5_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_11104, new_AGEMA_signal_11103, new_AGEMA_signal_11102, mcs1_mcs_mat1_5_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_12406, new_AGEMA_signal_12405, new_AGEMA_signal_12404, mcs1_mcs_mat1_5_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .c ({new_AGEMA_signal_11104, new_AGEMA_signal_11103, new_AGEMA_signal_11102, mcs1_mcs_mat1_5_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({new_AGEMA_signal_8992, new_AGEMA_signal_8991, new_AGEMA_signal_8990, mcs1_mcs_mat1_5_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({new_AGEMA_signal_8995, new_AGEMA_signal_8994, new_AGEMA_signal_8993, mcs1_mcs_mat1_5_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_11110, new_AGEMA_signal_11109, new_AGEMA_signal_11108, mcs1_mcs_mat1_5_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .b ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_12415, new_AGEMA_signal_12414, new_AGEMA_signal_12413, mcs1_mcs_mat1_5_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({new_AGEMA_signal_8995, new_AGEMA_signal_8994, new_AGEMA_signal_8993, mcs1_mcs_mat1_5_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_19171, new_AGEMA_signal_19170, new_AGEMA_signal_19169, mcs1_mcs_mat1_5_mcs_out[35]}), .b ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_19891, new_AGEMA_signal_19890, new_AGEMA_signal_19889, mcs1_mcs_mat1_5_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_18511, new_AGEMA_signal_18510, new_AGEMA_signal_18509, mcs1_mcs_mat1_5_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_13849, new_AGEMA_signal_13848, new_AGEMA_signal_13847, mcs1_mcs_mat1_5_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_19171, new_AGEMA_signal_19170, new_AGEMA_signal_19169, mcs1_mcs_mat1_5_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_17845, new_AGEMA_signal_17844, new_AGEMA_signal_17843, mcs1_mcs_mat1_5_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .c ({new_AGEMA_signal_18511, new_AGEMA_signal_18510, new_AGEMA_signal_18509, mcs1_mcs_mat1_5_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .c ({new_AGEMA_signal_17845, new_AGEMA_signal_17844, new_AGEMA_signal_17843, mcs1_mcs_mat1_5_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({new_AGEMA_signal_13849, new_AGEMA_signal_13848, new_AGEMA_signal_13847, mcs1_mcs_mat1_5_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_8998, new_AGEMA_signal_8997, new_AGEMA_signal_8996, mcs1_mcs_mat1_5_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_9871, new_AGEMA_signal_9870, new_AGEMA_signal_9869, mcs1_mcs_mat1_5_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({new_AGEMA_signal_12421, new_AGEMA_signal_12420, new_AGEMA_signal_12419, mcs1_mcs_mat1_5_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_13855, new_AGEMA_signal_13854, new_AGEMA_signal_13853, mcs1_mcs_mat1_5_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_8998, new_AGEMA_signal_8997, new_AGEMA_signal_8996, mcs1_mcs_mat1_5_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_12421, new_AGEMA_signal_12420, new_AGEMA_signal_12419, mcs1_mcs_mat1_5_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({new_AGEMA_signal_8998, new_AGEMA_signal_8997, new_AGEMA_signal_8996, mcs1_mcs_mat1_5_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({new_AGEMA_signal_9001, new_AGEMA_signal_9000, new_AGEMA_signal_8999, mcs1_mcs_mat1_5_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({new_AGEMA_signal_9004, new_AGEMA_signal_9003, new_AGEMA_signal_9002, mcs1_mcs_mat1_5_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_17170, new_AGEMA_signal_17169, new_AGEMA_signal_17168, mcs1_mcs_mat1_5_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_17851, new_AGEMA_signal_17850, new_AGEMA_signal_17849, mcs1_mcs_mat1_5_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_17170, new_AGEMA_signal_17169, new_AGEMA_signal_17168, mcs1_mcs_mat1_5_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .c ({new_AGEMA_signal_17857, new_AGEMA_signal_17856, new_AGEMA_signal_17855, mcs1_mcs_mat1_5_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({new_AGEMA_signal_13879, new_AGEMA_signal_13878, new_AGEMA_signal_13877, mcs1_mcs_mat1_5_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({new_AGEMA_signal_9007, new_AGEMA_signal_9006, new_AGEMA_signal_9005, mcs1_mcs_mat1_5_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({new_AGEMA_signal_9010, new_AGEMA_signal_9009, new_AGEMA_signal_9008, mcs1_mcs_mat1_5_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_9013, new_AGEMA_signal_9012, new_AGEMA_signal_9011, mcs1_mcs_mat1_5_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_11137, new_AGEMA_signal_11136, new_AGEMA_signal_11135, mcs1_mcs_mat1_5_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_9013, new_AGEMA_signal_9012, new_AGEMA_signal_9011, mcs1_mcs_mat1_5_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_9889, new_AGEMA_signal_9888, new_AGEMA_signal_9887, mcs1_mcs_mat1_5_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({new_AGEMA_signal_9013, new_AGEMA_signal_9012, new_AGEMA_signal_9011, mcs1_mcs_mat1_5_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_17869, new_AGEMA_signal_17868, new_AGEMA_signal_17867, mcs1_mcs_mat1_5_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_13900, new_AGEMA_signal_13899, new_AGEMA_signal_13898, mcs1_mcs_mat1_5_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_18523, new_AGEMA_signal_18522, new_AGEMA_signal_18521, mcs1_mcs_mat1_5_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_17869, new_AGEMA_signal_17868, new_AGEMA_signal_17867, mcs1_mcs_mat1_5_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .c ({new_AGEMA_signal_18529, new_AGEMA_signal_18528, new_AGEMA_signal_18527, mcs1_mcs_mat1_5_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_17182, new_AGEMA_signal_17181, new_AGEMA_signal_17180, mcs1_mcs_mat1_5_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_17869, new_AGEMA_signal_17868, new_AGEMA_signal_17867, mcs1_mcs_mat1_5_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_17182, new_AGEMA_signal_17181, new_AGEMA_signal_17180, mcs1_mcs_mat1_5_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .c ({new_AGEMA_signal_17872, new_AGEMA_signal_17871, new_AGEMA_signal_17870, mcs1_mcs_mat1_5_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({new_AGEMA_signal_13900, new_AGEMA_signal_13899, new_AGEMA_signal_13898, mcs1_mcs_mat1_5_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U44 ( .a ({new_AGEMA_signal_11182, new_AGEMA_signal_11181, new_AGEMA_signal_11180, mcs1_mcs_mat1_6_mcs_out[90]}), .b ({new_AGEMA_signal_12493, new_AGEMA_signal_12492, new_AGEMA_signal_12491, mcs1_mcs_mat1_6_mcs_out[94]}), .c ({new_AGEMA_signal_13906, new_AGEMA_signal_13905, new_AGEMA_signal_13904, mcs1_mcs_mat1_6_n93}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .c ({new_AGEMA_signal_11143, new_AGEMA_signal_11142, new_AGEMA_signal_11141, mcs1_mcs_mat1_6_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .b ({new_AGEMA_signal_9016, new_AGEMA_signal_9015, new_AGEMA_signal_9014, mcs1_mcs_mat1_6_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_9895, new_AGEMA_signal_9894, new_AGEMA_signal_9893, mcs1_mcs_mat1_6_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({new_AGEMA_signal_9016, new_AGEMA_signal_9015, new_AGEMA_signal_9014, mcs1_mcs_mat1_6_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_17230, new_AGEMA_signal_17229, new_AGEMA_signal_17228, mcs1_mcs_mat1_6_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_17890, new_AGEMA_signal_17889, new_AGEMA_signal_17888, mcs1_mcs_mat1_6_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_13918, new_AGEMA_signal_13917, new_AGEMA_signal_13916, mcs1_mcs_mat1_6_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_17230, new_AGEMA_signal_17229, new_AGEMA_signal_17228, mcs1_mcs_mat1_6_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({new_AGEMA_signal_13918, new_AGEMA_signal_13917, new_AGEMA_signal_13916, mcs1_mcs_mat1_6_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_9019, new_AGEMA_signal_9018, new_AGEMA_signal_9017, mcs1_mcs_mat1_6_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_12472, new_AGEMA_signal_12471, new_AGEMA_signal_12470, mcs1_mcs_mat1_6_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_13921, new_AGEMA_signal_13920, new_AGEMA_signal_13919, mcs1_mcs_mat1_6_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_9901, new_AGEMA_signal_9900, new_AGEMA_signal_9899, mcs1_mcs_mat1_6_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_11152, new_AGEMA_signal_11151, new_AGEMA_signal_11150, mcs1_mcs_mat1_6_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .c ({new_AGEMA_signal_9901, new_AGEMA_signal_9900, new_AGEMA_signal_9899, mcs1_mcs_mat1_6_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .b ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_12472, new_AGEMA_signal_12471, new_AGEMA_signal_12470, mcs1_mcs_mat1_6_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({new_AGEMA_signal_9019, new_AGEMA_signal_9018, new_AGEMA_signal_9017, mcs1_mcs_mat1_6_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_12478, new_AGEMA_signal_12477, new_AGEMA_signal_12476, mcs1_mcs_mat1_6_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_13930, new_AGEMA_signal_13929, new_AGEMA_signal_13928, mcs1_mcs_mat1_6_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_9022, new_AGEMA_signal_9021, new_AGEMA_signal_9020, mcs1_mcs_mat1_6_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_12478, new_AGEMA_signal_12477, new_AGEMA_signal_12476, mcs1_mcs_mat1_6_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({new_AGEMA_signal_9022, new_AGEMA_signal_9021, new_AGEMA_signal_9020, mcs1_mcs_mat1_6_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({new_AGEMA_signal_9025, new_AGEMA_signal_9024, new_AGEMA_signal_9023, mcs1_mcs_mat1_6_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({new_AGEMA_signal_17239, new_AGEMA_signal_17238, new_AGEMA_signal_17237, mcs1_mcs_mat1_6_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_17899, new_AGEMA_signal_17898, new_AGEMA_signal_17897, mcs1_mcs_mat1_6_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_13942, new_AGEMA_signal_13941, new_AGEMA_signal_13940, mcs1_mcs_mat1_6_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_17239, new_AGEMA_signal_17238, new_AGEMA_signal_17237, mcs1_mcs_mat1_6_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .b ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .c ({new_AGEMA_signal_17902, new_AGEMA_signal_17901, new_AGEMA_signal_17900, mcs1_mcs_mat1_6_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({new_AGEMA_signal_13942, new_AGEMA_signal_13941, new_AGEMA_signal_13940, mcs1_mcs_mat1_6_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_9028, new_AGEMA_signal_9027, new_AGEMA_signal_9026, mcs1_mcs_mat1_6_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_11167, new_AGEMA_signal_11166, new_AGEMA_signal_11165, mcs1_mcs_mat1_6_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_9028, new_AGEMA_signal_9027, new_AGEMA_signal_9026, mcs1_mcs_mat1_6_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .c ({new_AGEMA_signal_9913, new_AGEMA_signal_9912, new_AGEMA_signal_9911, mcs1_mcs_mat1_6_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({new_AGEMA_signal_9028, new_AGEMA_signal_9027, new_AGEMA_signal_9026, mcs1_mcs_mat1_6_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_11173, new_AGEMA_signal_11172, new_AGEMA_signal_11171, mcs1_mcs_mat1_6_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .c ({new_AGEMA_signal_12493, new_AGEMA_signal_12492, new_AGEMA_signal_12491, mcs1_mcs_mat1_6_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_9031, new_AGEMA_signal_9030, new_AGEMA_signal_9029, mcs1_mcs_mat1_6_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_11173, new_AGEMA_signal_11172, new_AGEMA_signal_11171, mcs1_mcs_mat1_6_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_11176, new_AGEMA_signal_11175, new_AGEMA_signal_11174, mcs1_mcs_mat1_6_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({new_AGEMA_signal_9031, new_AGEMA_signal_9030, new_AGEMA_signal_9029, mcs1_mcs_mat1_6_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .b ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .c ({new_AGEMA_signal_11182, new_AGEMA_signal_11181, new_AGEMA_signal_11180, mcs1_mcs_mat1_6_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .b ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_11185, new_AGEMA_signal_11184, new_AGEMA_signal_11183, mcs1_mcs_mat1_6_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({new_AGEMA_signal_17914, new_AGEMA_signal_17913, new_AGEMA_signal_17912, mcs1_mcs_mat1_6_mcs_out[87]}), .c ({new_AGEMA_signal_18565, new_AGEMA_signal_18564, new_AGEMA_signal_18563, mcs1_mcs_mat1_6_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .c ({new_AGEMA_signal_17914, new_AGEMA_signal_17913, new_AGEMA_signal_17912, mcs1_mcs_mat1_6_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .c ({new_AGEMA_signal_12508, new_AGEMA_signal_12507, new_AGEMA_signal_12506, mcs1_mcs_mat1_6_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({new_AGEMA_signal_9034, new_AGEMA_signal_9033, new_AGEMA_signal_9032, mcs1_mcs_mat1_6_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_9037, new_AGEMA_signal_9036, new_AGEMA_signal_9035, mcs1_mcs_mat1_6_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_9925, new_AGEMA_signal_9924, new_AGEMA_signal_9923, mcs1_mcs_mat1_6_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({new_AGEMA_signal_9037, new_AGEMA_signal_9036, new_AGEMA_signal_9035, mcs1_mcs_mat1_6_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_9040, new_AGEMA_signal_9039, new_AGEMA_signal_9038, mcs1_mcs_mat1_6_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_9931, new_AGEMA_signal_9930, new_AGEMA_signal_9929, mcs1_mcs_mat1_6_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({new_AGEMA_signal_9040, new_AGEMA_signal_9039, new_AGEMA_signal_9038, mcs1_mcs_mat1_6_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({new_AGEMA_signal_13972, new_AGEMA_signal_13971, new_AGEMA_signal_13970, mcs1_mcs_mat1_6_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_9043, new_AGEMA_signal_9042, new_AGEMA_signal_9041, mcs1_mcs_mat1_6_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .c ({new_AGEMA_signal_12529, new_AGEMA_signal_12528, new_AGEMA_signal_12527, mcs1_mcs_mat1_6_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({new_AGEMA_signal_9043, new_AGEMA_signal_9042, new_AGEMA_signal_9041, mcs1_mcs_mat1_6_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_15427, new_AGEMA_signal_15426, new_AGEMA_signal_15425, mcs1_mcs_mat1_6_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_9046, new_AGEMA_signal_9045, new_AGEMA_signal_9044, mcs1_mcs_mat1_6_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_16459, new_AGEMA_signal_16458, new_AGEMA_signal_16457, mcs1_mcs_mat1_6_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_13984, new_AGEMA_signal_13983, new_AGEMA_signal_13982, mcs1_mcs_mat1_6_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_15427, new_AGEMA_signal_15426, new_AGEMA_signal_15425, mcs1_mcs_mat1_6_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_12535, new_AGEMA_signal_12534, new_AGEMA_signal_12533, mcs1_mcs_mat1_6_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_13984, new_AGEMA_signal_13983, new_AGEMA_signal_13982, mcs1_mcs_mat1_6_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_12535, new_AGEMA_signal_12534, new_AGEMA_signal_12533, mcs1_mcs_mat1_6_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({new_AGEMA_signal_9046, new_AGEMA_signal_9045, new_AGEMA_signal_9044, mcs1_mcs_mat1_6_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_12544, new_AGEMA_signal_12543, new_AGEMA_signal_12542, mcs1_mcs_mat1_6_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_9943, new_AGEMA_signal_9942, new_AGEMA_signal_9941, mcs1_mcs_mat1_6_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_13987, new_AGEMA_signal_13986, new_AGEMA_signal_13985, mcs1_mcs_mat1_6_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_9049, new_AGEMA_signal_9048, new_AGEMA_signal_9047, mcs1_mcs_mat1_6_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .c ({new_AGEMA_signal_9943, new_AGEMA_signal_9942, new_AGEMA_signal_9941, mcs1_mcs_mat1_6_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .c ({new_AGEMA_signal_9946, new_AGEMA_signal_9945, new_AGEMA_signal_9944, mcs1_mcs_mat1_6_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .c ({new_AGEMA_signal_12544, new_AGEMA_signal_12543, new_AGEMA_signal_12542, mcs1_mcs_mat1_6_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_9049, new_AGEMA_signal_9048, new_AGEMA_signal_9047, mcs1_mcs_mat1_6_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_12547, new_AGEMA_signal_12546, new_AGEMA_signal_12545, mcs1_mcs_mat1_6_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({new_AGEMA_signal_9049, new_AGEMA_signal_9048, new_AGEMA_signal_9047, mcs1_mcs_mat1_6_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .b ({new_AGEMA_signal_13996, new_AGEMA_signal_13995, new_AGEMA_signal_13994, mcs1_mcs_mat1_6_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_17932, new_AGEMA_signal_17931, new_AGEMA_signal_17930, mcs1_mcs_mat1_6_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({new_AGEMA_signal_13996, new_AGEMA_signal_13995, new_AGEMA_signal_13994, mcs1_mcs_mat1_6_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({new_AGEMA_signal_12553, new_AGEMA_signal_12552, new_AGEMA_signal_12551, mcs1_mcs_mat1_6_mcs_out[51]}), .c ({new_AGEMA_signal_13999, new_AGEMA_signal_13998, new_AGEMA_signal_13997, mcs1_mcs_mat1_6_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .c ({new_AGEMA_signal_12553, new_AGEMA_signal_12552, new_AGEMA_signal_12551, mcs1_mcs_mat1_6_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_9052, new_AGEMA_signal_9051, new_AGEMA_signal_9050, mcs1_mcs_mat1_6_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_11206, new_AGEMA_signal_11205, new_AGEMA_signal_11204, mcs1_mcs_mat1_6_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({new_AGEMA_signal_9052, new_AGEMA_signal_9051, new_AGEMA_signal_9050, mcs1_mcs_mat1_6_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_12562, new_AGEMA_signal_12561, new_AGEMA_signal_12560, mcs1_mcs_mat1_6_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_14008, new_AGEMA_signal_14007, new_AGEMA_signal_14006, mcs1_mcs_mat1_6_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_12562, new_AGEMA_signal_12561, new_AGEMA_signal_12560, mcs1_mcs_mat1_6_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_11212, new_AGEMA_signal_11211, new_AGEMA_signal_11210, mcs1_mcs_mat1_6_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_12565, new_AGEMA_signal_12564, new_AGEMA_signal_12563, mcs1_mcs_mat1_6_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .c ({new_AGEMA_signal_11212, new_AGEMA_signal_11211, new_AGEMA_signal_11210, mcs1_mcs_mat1_6_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({new_AGEMA_signal_9055, new_AGEMA_signal_9054, new_AGEMA_signal_9053, mcs1_mcs_mat1_6_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({new_AGEMA_signal_14017, new_AGEMA_signal_14016, new_AGEMA_signal_14015, mcs1_mcs_mat1_6_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_17263, new_AGEMA_signal_17262, new_AGEMA_signal_17261, mcs1_mcs_mat1_6_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .b ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_17941, new_AGEMA_signal_17940, new_AGEMA_signal_17939, mcs1_mcs_mat1_6_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({new_AGEMA_signal_14017, new_AGEMA_signal_14016, new_AGEMA_signal_14015, mcs1_mcs_mat1_6_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_15451, new_AGEMA_signal_15450, new_AGEMA_signal_15449, mcs1_mcs_mat1_6_mcs_out[35]}), .b ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_16468, new_AGEMA_signal_16467, new_AGEMA_signal_16466, mcs1_mcs_mat1_6_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_14023, new_AGEMA_signal_14022, new_AGEMA_signal_14021, mcs1_mcs_mat1_6_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_9058, new_AGEMA_signal_9057, new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_15451, new_AGEMA_signal_15450, new_AGEMA_signal_15449, mcs1_mcs_mat1_6_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_12571, new_AGEMA_signal_12570, new_AGEMA_signal_12569, mcs1_mcs_mat1_6_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .c ({new_AGEMA_signal_14023, new_AGEMA_signal_14022, new_AGEMA_signal_14021, mcs1_mcs_mat1_6_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .c ({new_AGEMA_signal_12571, new_AGEMA_signal_12570, new_AGEMA_signal_12569, mcs1_mcs_mat1_6_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466]}), .c ({new_AGEMA_signal_9058, new_AGEMA_signal_9057, new_AGEMA_signal_9056, mcs1_mcs_mat1_6_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_9061, new_AGEMA_signal_9060, new_AGEMA_signal_9059, mcs1_mcs_mat1_6_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_9961, new_AGEMA_signal_9960, new_AGEMA_signal_9959, mcs1_mcs_mat1_6_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({new_AGEMA_signal_12577, new_AGEMA_signal_12576, new_AGEMA_signal_12575, mcs1_mcs_mat1_6_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_14029, new_AGEMA_signal_14028, new_AGEMA_signal_14027, mcs1_mcs_mat1_6_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_9061, new_AGEMA_signal_9060, new_AGEMA_signal_9059, mcs1_mcs_mat1_6_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_12577, new_AGEMA_signal_12576, new_AGEMA_signal_12575, mcs1_mcs_mat1_6_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({new_AGEMA_signal_9061, new_AGEMA_signal_9060, new_AGEMA_signal_9059, mcs1_mcs_mat1_6_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478]}), .c ({new_AGEMA_signal_9064, new_AGEMA_signal_9063, new_AGEMA_signal_9062, mcs1_mcs_mat1_6_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({new_AGEMA_signal_14044, new_AGEMA_signal_14043, new_AGEMA_signal_14042, mcs1_mcs_mat1_6_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_11227, new_AGEMA_signal_11226, new_AGEMA_signal_11225, mcs1_mcs_mat1_6_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_12595, new_AGEMA_signal_12594, new_AGEMA_signal_12593, mcs1_mcs_mat1_6_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_11227, new_AGEMA_signal_11226, new_AGEMA_signal_11225, mcs1_mcs_mat1_6_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .c ({new_AGEMA_signal_12601, new_AGEMA_signal_12600, new_AGEMA_signal_12599, mcs1_mcs_mat1_6_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({new_AGEMA_signal_9067, new_AGEMA_signal_9066, new_AGEMA_signal_9065, mcs1_mcs_mat1_6_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({new_AGEMA_signal_9070, new_AGEMA_signal_9069, new_AGEMA_signal_9068, mcs1_mcs_mat1_6_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502]}), .c ({new_AGEMA_signal_9073, new_AGEMA_signal_9072, new_AGEMA_signal_9071, mcs1_mcs_mat1_6_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_14071, new_AGEMA_signal_14070, new_AGEMA_signal_14069, mcs1_mcs_mat1_6_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_17281, new_AGEMA_signal_17280, new_AGEMA_signal_17279, mcs1_mcs_mat1_6_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_14071, new_AGEMA_signal_14070, new_AGEMA_signal_14069, mcs1_mcs_mat1_6_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_15493, new_AGEMA_signal_15492, new_AGEMA_signal_15491, mcs1_mcs_mat1_6_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({new_AGEMA_signal_14071, new_AGEMA_signal_14070, new_AGEMA_signal_14069, mcs1_mcs_mat1_6_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_12622, new_AGEMA_signal_12621, new_AGEMA_signal_12620, mcs1_mcs_mat1_6_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_9076, new_AGEMA_signal_9075, new_AGEMA_signal_9074, mcs1_mcs_mat1_6_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_14074, new_AGEMA_signal_14073, new_AGEMA_signal_14072, mcs1_mcs_mat1_6_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_12622, new_AGEMA_signal_12621, new_AGEMA_signal_12620, mcs1_mcs_mat1_6_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .c ({new_AGEMA_signal_14080, new_AGEMA_signal_14079, new_AGEMA_signal_14078, mcs1_mcs_mat1_6_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_11242, new_AGEMA_signal_11241, new_AGEMA_signal_11240, mcs1_mcs_mat1_6_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_12622, new_AGEMA_signal_12621, new_AGEMA_signal_12620, mcs1_mcs_mat1_6_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_11242, new_AGEMA_signal_11241, new_AGEMA_signal_11240, mcs1_mcs_mat1_6_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .c ({new_AGEMA_signal_12625, new_AGEMA_signal_12624, new_AGEMA_signal_12623, mcs1_mcs_mat1_6_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514]}), .c ({new_AGEMA_signal_9076, new_AGEMA_signal_9075, new_AGEMA_signal_9074, mcs1_mcs_mat1_6_mcs_rom0_31_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U44 ( .a ({new_AGEMA_signal_17350, new_AGEMA_signal_17349, new_AGEMA_signal_17348, mcs1_mcs_mat1_7_mcs_out[90]}), .b ({new_AGEMA_signal_12670, new_AGEMA_signal_12669, new_AGEMA_signal_12668, mcs1_mcs_mat1_7_mcs_out[94]}), .c ({new_AGEMA_signal_17968, new_AGEMA_signal_17967, new_AGEMA_signal_17966, mcs1_mcs_mat1_7_n93}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_0_U1 ( .a ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .c ({new_AGEMA_signal_11248, new_AGEMA_signal_11247, new_AGEMA_signal_11246, mcs1_mcs_mat1_7_mcs_out[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U6 ( .a ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .b ({new_AGEMA_signal_14086, new_AGEMA_signal_14085, new_AGEMA_signal_14084, mcs1_mcs_mat1_7_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_15526, new_AGEMA_signal_15525, new_AGEMA_signal_15524, mcs1_mcs_mat1_7_mcs_rom0_1_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({new_AGEMA_signal_14086, new_AGEMA_signal_14085, new_AGEMA_signal_14084, mcs1_mcs_mat1_7_mcs_rom0_1_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U6 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_11251, new_AGEMA_signal_11250, new_AGEMA_signal_11249, mcs1_mcs_mat1_7_mcs_rom0_2_n9}), .c ({new_AGEMA_signal_12631, new_AGEMA_signal_12630, new_AGEMA_signal_12629, mcs1_mcs_mat1_7_mcs_rom0_2_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U5 ( .a ({new_AGEMA_signal_9079, new_AGEMA_signal_9078, new_AGEMA_signal_9077, mcs1_mcs_mat1_7_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_11251, new_AGEMA_signal_11250, new_AGEMA_signal_11249, mcs1_mcs_mat1_7_mcs_rom0_2_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526]}), .c ({new_AGEMA_signal_9079, new_AGEMA_signal_9078, new_AGEMA_signal_9077, mcs1_mcs_mat1_7_mcs_rom0_2_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U9 ( .a ({new_AGEMA_signal_9082, new_AGEMA_signal_9081, new_AGEMA_signal_9080, mcs1_mcs_mat1_7_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_12643, new_AGEMA_signal_12642, new_AGEMA_signal_12641, mcs1_mcs_mat1_7_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_14095, new_AGEMA_signal_14094, new_AGEMA_signal_14093, mcs1_mcs_mat1_7_mcs_out[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U7 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_9985, new_AGEMA_signal_9984, new_AGEMA_signal_9983, mcs1_mcs_mat1_7_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_11260, new_AGEMA_signal_11259, new_AGEMA_signal_11258, mcs1_mcs_mat1_7_mcs_rom0_3_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U6 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .c ({new_AGEMA_signal_9985, new_AGEMA_signal_9984, new_AGEMA_signal_9983, mcs1_mcs_mat1_7_mcs_rom0_3_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U1 ( .a ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_12643, new_AGEMA_signal_12642, new_AGEMA_signal_12641, mcs1_mcs_mat1_7_mcs_rom0_3_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({new_AGEMA_signal_9082, new_AGEMA_signal_9081, new_AGEMA_signal_9080, mcs1_mcs_mat1_7_mcs_rom0_3_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U5 ( .a ({new_AGEMA_signal_12649, new_AGEMA_signal_12648, new_AGEMA_signal_12647, mcs1_mcs_mat1_7_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_14104, new_AGEMA_signal_14103, new_AGEMA_signal_14102, mcs1_mcs_mat1_7_mcs_rom0_4_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U1 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_9085, new_AGEMA_signal_9084, new_AGEMA_signal_9083, mcs1_mcs_mat1_7_mcs_rom0_4_x0x4}), .c ({new_AGEMA_signal_12649, new_AGEMA_signal_12648, new_AGEMA_signal_12647, mcs1_mcs_mat1_7_mcs_rom0_4_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538]}), .c ({new_AGEMA_signal_9085, new_AGEMA_signal_9084, new_AGEMA_signal_9083, mcs1_mcs_mat1_7_mcs_rom0_4_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({new_AGEMA_signal_14110, new_AGEMA_signal_14109, new_AGEMA_signal_14108, mcs1_mcs_mat1_7_mcs_rom0_5_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U7 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({new_AGEMA_signal_11269, new_AGEMA_signal_11268, new_AGEMA_signal_11267, mcs1_mcs_mat1_7_mcs_rom0_6_n10}), .c ({new_AGEMA_signal_12655, new_AGEMA_signal_12654, new_AGEMA_signal_12653, mcs1_mcs_mat1_7_mcs_out[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U6 ( .a ({new_AGEMA_signal_9088, new_AGEMA_signal_9087, new_AGEMA_signal_9086, mcs1_mcs_mat1_7_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_11269, new_AGEMA_signal_11268, new_AGEMA_signal_11267, mcs1_mcs_mat1_7_mcs_rom0_6_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U4 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .b ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .c ({new_AGEMA_signal_12658, new_AGEMA_signal_12657, new_AGEMA_signal_12656, mcs1_mcs_mat1_7_mcs_rom0_6_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({new_AGEMA_signal_9088, new_AGEMA_signal_9087, new_AGEMA_signal_9086, mcs1_mcs_mat1_7_mcs_rom0_6_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U7 ( .a ({new_AGEMA_signal_9091, new_AGEMA_signal_9090, new_AGEMA_signal_9089, mcs1_mcs_mat1_7_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_11275, new_AGEMA_signal_11274, new_AGEMA_signal_11273, mcs1_mcs_mat1_7_mcs_out[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U1 ( .a ({new_AGEMA_signal_9091, new_AGEMA_signal_9090, new_AGEMA_signal_9089, mcs1_mcs_mat1_7_mcs_rom0_7_x0x4}), .b ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .c ({new_AGEMA_signal_9997, new_AGEMA_signal_9996, new_AGEMA_signal_9995, mcs1_mcs_mat1_7_mcs_rom0_7_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({new_AGEMA_signal_9091, new_AGEMA_signal_9090, new_AGEMA_signal_9089, mcs1_mcs_mat1_7_mcs_rom0_7_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U7 ( .a ({new_AGEMA_signal_11281, new_AGEMA_signal_11280, new_AGEMA_signal_11279, mcs1_mcs_mat1_7_mcs_rom0_8_n7}), .b ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .c ({new_AGEMA_signal_12670, new_AGEMA_signal_12669, new_AGEMA_signal_12668, mcs1_mcs_mat1_7_mcs_out[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U6 ( .a ({new_AGEMA_signal_9094, new_AGEMA_signal_9093, new_AGEMA_signal_9092, mcs1_mcs_mat1_7_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_11281, new_AGEMA_signal_11280, new_AGEMA_signal_11279, mcs1_mcs_mat1_7_mcs_rom0_8_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U4 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_11284, new_AGEMA_signal_11283, new_AGEMA_signal_11282, mcs1_mcs_mat1_7_mcs_rom0_8_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562]}), .c ({new_AGEMA_signal_9094, new_AGEMA_signal_9093, new_AGEMA_signal_9092, mcs1_mcs_mat1_7_mcs_rom0_8_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_9_U2 ( .a ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .c ({new_AGEMA_signal_17350, new_AGEMA_signal_17349, new_AGEMA_signal_17348, mcs1_mcs_mat1_7_mcs_out[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_9_U1 ( .a ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .b ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_17353, new_AGEMA_signal_17352, new_AGEMA_signal_17351, mcs1_mcs_mat1_7_mcs_out[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_10_U2 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({new_AGEMA_signal_12679, new_AGEMA_signal_12678, new_AGEMA_signal_12677, mcs1_mcs_mat1_7_mcs_out[87]}), .c ({new_AGEMA_signal_14128, new_AGEMA_signal_14127, new_AGEMA_signal_14126, mcs1_mcs_mat1_7_mcs_out[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_10_U1 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .c ({new_AGEMA_signal_12679, new_AGEMA_signal_12678, new_AGEMA_signal_12677, mcs1_mcs_mat1_7_mcs_out[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .c ({new_AGEMA_signal_12688, new_AGEMA_signal_12687, new_AGEMA_signal_12686, mcs1_mcs_mat1_7_mcs_rom0_11_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({new_AGEMA_signal_9097, new_AGEMA_signal_9096, new_AGEMA_signal_9095, mcs1_mcs_mat1_7_mcs_rom0_11_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U5 ( .a ({new_AGEMA_signal_9100, new_AGEMA_signal_9099, new_AGEMA_signal_9098, mcs1_mcs_mat1_7_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_10009, new_AGEMA_signal_10008, new_AGEMA_signal_10007, mcs1_mcs_mat1_7_mcs_out[78]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574]}), .c ({new_AGEMA_signal_9100, new_AGEMA_signal_9099, new_AGEMA_signal_9098, mcs1_mcs_mat1_7_mcs_rom0_12_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U3 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_14146, new_AGEMA_signal_14145, new_AGEMA_signal_14144, mcs1_mcs_mat1_7_mcs_rom0_13_x0x4}), .c ({new_AGEMA_signal_15580, new_AGEMA_signal_15579, new_AGEMA_signal_15578, mcs1_mcs_mat1_7_mcs_rom0_13_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({new_AGEMA_signal_14146, new_AGEMA_signal_14145, new_AGEMA_signal_14144, mcs1_mcs_mat1_7_mcs_rom0_13_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586]}), .c ({new_AGEMA_signal_9103, new_AGEMA_signal_9102, new_AGEMA_signal_9101, mcs1_mcs_mat1_7_mcs_rom0_14_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U5 ( .a ({new_AGEMA_signal_9106, new_AGEMA_signal_9105, new_AGEMA_signal_9104, mcs1_mcs_mat1_7_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .c ({new_AGEMA_signal_12709, new_AGEMA_signal_12708, new_AGEMA_signal_12707, mcs1_mcs_mat1_7_mcs_out[65]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({new_AGEMA_signal_9106, new_AGEMA_signal_9105, new_AGEMA_signal_9104, mcs1_mcs_mat1_7_mcs_rom0_15_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U4 ( .a ({new_AGEMA_signal_15604, new_AGEMA_signal_15603, new_AGEMA_signal_15602, mcs1_mcs_mat1_7_mcs_rom0_16_n4}), .b ({new_AGEMA_signal_9109, new_AGEMA_signal_9108, new_AGEMA_signal_9107, mcs1_mcs_mat1_7_mcs_rom0_16_x0x4}), .c ({new_AGEMA_signal_16555, new_AGEMA_signal_16554, new_AGEMA_signal_16553, mcs1_mcs_mat1_7_mcs_out[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U3 ( .a ({new_AGEMA_signal_14164, new_AGEMA_signal_14163, new_AGEMA_signal_14162, mcs1_mcs_mat1_7_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_15604, new_AGEMA_signal_15603, new_AGEMA_signal_15602, mcs1_mcs_mat1_7_mcs_rom0_16_n4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U2 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_12715, new_AGEMA_signal_12714, new_AGEMA_signal_12713, mcs1_mcs_mat1_7_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_14164, new_AGEMA_signal_14163, new_AGEMA_signal_14162, mcs1_mcs_mat1_7_mcs_rom0_16_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_12715, new_AGEMA_signal_12714, new_AGEMA_signal_12713, mcs1_mcs_mat1_7_mcs_rom0_16_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598]}), .c ({new_AGEMA_signal_9109, new_AGEMA_signal_9108, new_AGEMA_signal_9107, mcs1_mcs_mat1_7_mcs_rom0_16_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U9 ( .a ({new_AGEMA_signal_18010, new_AGEMA_signal_18009, new_AGEMA_signal_18008, mcs1_mcs_mat1_7_mcs_rom0_17_n10}), .b ({new_AGEMA_signal_15607, new_AGEMA_signal_15606, new_AGEMA_signal_15605, mcs1_mcs_mat1_7_mcs_rom0_17_n9}), .c ({new_AGEMA_signal_18640, new_AGEMA_signal_18639, new_AGEMA_signal_18638, mcs1_mcs_mat1_7_mcs_out[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U8 ( .a ({new_AGEMA_signal_14167, new_AGEMA_signal_14166, new_AGEMA_signal_14165, mcs1_mcs_mat1_7_mcs_rom0_17_x0x4}), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .c ({new_AGEMA_signal_15607, new_AGEMA_signal_15606, new_AGEMA_signal_15605, mcs1_mcs_mat1_7_mcs_rom0_17_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U6 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .c ({new_AGEMA_signal_15610, new_AGEMA_signal_15609, new_AGEMA_signal_15608, mcs1_mcs_mat1_7_mcs_rom0_17_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U4 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .c ({new_AGEMA_signal_18010, new_AGEMA_signal_18009, new_AGEMA_signal_18008, mcs1_mcs_mat1_7_mcs_rom0_17_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U2 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_14167, new_AGEMA_signal_14166, new_AGEMA_signal_14165, mcs1_mcs_mat1_7_mcs_rom0_17_x0x4}), .c ({new_AGEMA_signal_18013, new_AGEMA_signal_18012, new_AGEMA_signal_18011, mcs1_mcs_mat1_7_mcs_rom0_17_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({new_AGEMA_signal_14167, new_AGEMA_signal_14166, new_AGEMA_signal_14165, mcs1_mcs_mat1_7_mcs_rom0_17_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U1 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .b ({new_AGEMA_signal_9112, new_AGEMA_signal_9111, new_AGEMA_signal_9110, mcs1_mcs_mat1_7_mcs_rom0_18_x0x4}), .c ({new_AGEMA_signal_12727, new_AGEMA_signal_12726, new_AGEMA_signal_12725, mcs1_mcs_mat1_7_mcs_rom0_18_n9}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({new_AGEMA_signal_9112, new_AGEMA_signal_9111, new_AGEMA_signal_9110, mcs1_mcs_mat1_7_mcs_rom0_18_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_19_U2 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({new_AGEMA_signal_12733, new_AGEMA_signal_12732, new_AGEMA_signal_12731, mcs1_mcs_mat1_7_mcs_out[51]}), .c ({new_AGEMA_signal_14176, new_AGEMA_signal_14175, new_AGEMA_signal_14174, mcs1_mcs_mat1_7_mcs_out[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_19_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .c ({new_AGEMA_signal_12733, new_AGEMA_signal_12732, new_AGEMA_signal_12731, mcs1_mcs_mat1_7_mcs_out[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U6 ( .a ({new_AGEMA_signal_9115, new_AGEMA_signal_9114, new_AGEMA_signal_9113, mcs1_mcs_mat1_7_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_11311, new_AGEMA_signal_11310, new_AGEMA_signal_11309, mcs1_mcs_mat1_7_mcs_out[46]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({new_AGEMA_signal_9115, new_AGEMA_signal_9114, new_AGEMA_signal_9113, mcs1_mcs_mat1_7_mcs_rom0_20_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U7 ( .a ({new_AGEMA_signal_18019, new_AGEMA_signal_18018, new_AGEMA_signal_18017, mcs1_mcs_mat1_7_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_18652, new_AGEMA_signal_18651, new_AGEMA_signal_18650, mcs1_mcs_mat1_7_mcs_rom0_21_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U4 ( .a ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .b ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_18019, new_AGEMA_signal_18018, new_AGEMA_signal_18017, mcs1_mcs_mat1_7_mcs_rom0_21_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U2 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_17368, new_AGEMA_signal_17367, new_AGEMA_signal_17366, mcs1_mcs_mat1_7_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_18022, new_AGEMA_signal_18021, new_AGEMA_signal_18020, mcs1_mcs_mat1_7_mcs_rom0_21_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U1 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .c ({new_AGEMA_signal_17368, new_AGEMA_signal_17367, new_AGEMA_signal_17366, mcs1_mcs_mat1_7_mcs_rom0_21_n11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622]}), .c ({new_AGEMA_signal_14182, new_AGEMA_signal_14181, new_AGEMA_signal_14180, mcs1_mcs_mat1_7_mcs_rom0_21_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U8 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({new_AGEMA_signal_9118, new_AGEMA_signal_9117, new_AGEMA_signal_9116, mcs1_mcs_mat1_7_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_11317, new_AGEMA_signal_11316, new_AGEMA_signal_11315, mcs1_mcs_mat1_7_mcs_rom0_22_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U4 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_12745, new_AGEMA_signal_12744, new_AGEMA_signal_12743, mcs1_mcs_mat1_7_mcs_rom0_22_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({new_AGEMA_signal_9118, new_AGEMA_signal_9117, new_AGEMA_signal_9116, mcs1_mcs_mat1_7_mcs_rom0_22_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U4 ( .a ({new_AGEMA_signal_15634, new_AGEMA_signal_15633, new_AGEMA_signal_15632, mcs1_mcs_mat1_7_mcs_out[35]}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_16573, new_AGEMA_signal_16572, new_AGEMA_signal_16571, mcs1_mcs_mat1_7_mcs_rom0_23_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U3 ( .a ({new_AGEMA_signal_14194, new_AGEMA_signal_14193, new_AGEMA_signal_14192, mcs1_mcs_mat1_7_mcs_rom0_23_n4}), .b ({new_AGEMA_signal_9121, new_AGEMA_signal_9120, new_AGEMA_signal_9119, mcs1_mcs_mat1_7_mcs_rom0_23_x0x4}), .c ({new_AGEMA_signal_15634, new_AGEMA_signal_15633, new_AGEMA_signal_15632, mcs1_mcs_mat1_7_mcs_out[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U2 ( .a ({new_AGEMA_signal_12751, new_AGEMA_signal_12750, new_AGEMA_signal_12749, mcs1_mcs_mat1_7_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .c ({new_AGEMA_signal_14194, new_AGEMA_signal_14193, new_AGEMA_signal_14192, mcs1_mcs_mat1_7_mcs_rom0_23_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .c ({new_AGEMA_signal_12751, new_AGEMA_signal_12750, new_AGEMA_signal_12749, mcs1_mcs_mat1_7_mcs_rom0_23_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634]}), .c ({new_AGEMA_signal_9121, new_AGEMA_signal_9120, new_AGEMA_signal_9119, mcs1_mcs_mat1_7_mcs_rom0_23_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U7 ( .a ({new_AGEMA_signal_9124, new_AGEMA_signal_9123, new_AGEMA_signal_9122, mcs1_mcs_mat1_7_mcs_rom0_24_x0x4}), .b ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_10036, new_AGEMA_signal_10035, new_AGEMA_signal_10034, mcs1_mcs_mat1_7_mcs_rom0_24_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U6 ( .a ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({new_AGEMA_signal_12757, new_AGEMA_signal_12756, new_AGEMA_signal_12755, mcs1_mcs_mat1_7_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_14200, new_AGEMA_signal_14199, new_AGEMA_signal_14198, mcs1_mcs_mat1_7_mcs_out[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U4 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_9124, new_AGEMA_signal_9123, new_AGEMA_signal_9122, mcs1_mcs_mat1_7_mcs_rom0_24_x0x4}), .c ({new_AGEMA_signal_12757, new_AGEMA_signal_12756, new_AGEMA_signal_12755, mcs1_mcs_mat1_7_mcs_rom0_24_n12}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({new_AGEMA_signal_9124, new_AGEMA_signal_9123, new_AGEMA_signal_9122, mcs1_mcs_mat1_7_mcs_rom0_24_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646]}), .c ({new_AGEMA_signal_14206, new_AGEMA_signal_14205, new_AGEMA_signal_14204, mcs1_mcs_mat1_7_mcs_rom0_25_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652]}), .c ({new_AGEMA_signal_9127, new_AGEMA_signal_9126, new_AGEMA_signal_9125, mcs1_mcs_mat1_7_mcs_rom0_26_x0x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U9 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_11335, new_AGEMA_signal_11334, new_AGEMA_signal_11333, mcs1_mcs_mat1_7_mcs_rom0_27_n11}), .c ({new_AGEMA_signal_12775, new_AGEMA_signal_12774, new_AGEMA_signal_12773, mcs1_mcs_mat1_7_mcs_rom0_27_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U3 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_11335, new_AGEMA_signal_11334, new_AGEMA_signal_11333, mcs1_mcs_mat1_7_mcs_rom0_27_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U1 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .c ({new_AGEMA_signal_12781, new_AGEMA_signal_12780, new_AGEMA_signal_12779, mcs1_mcs_mat1_7_mcs_rom0_27_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658]}), .c ({new_AGEMA_signal_9130, new_AGEMA_signal_9129, new_AGEMA_signal_9128, mcs1_mcs_mat1_7_mcs_rom0_27_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664]}), .c ({new_AGEMA_signal_9133, new_AGEMA_signal_9132, new_AGEMA_signal_9131, mcs1_mcs_mat1_7_mcs_rom0_28_x0x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x0x4_AND_U1 ( .a ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({new_AGEMA_signal_14236, new_AGEMA_signal_14235, new_AGEMA_signal_14234, mcs1_mcs_mat1_7_mcs_rom0_29_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U7 ( .a ({new_AGEMA_signal_9136, new_AGEMA_signal_9135, new_AGEMA_signal_9134, mcs1_mcs_mat1_7_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_11344, new_AGEMA_signal_11343, new_AGEMA_signal_11342, mcs1_mcs_mat1_7_mcs_out[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U1 ( .a ({new_AGEMA_signal_9136, new_AGEMA_signal_9135, new_AGEMA_signal_9134, mcs1_mcs_mat1_7_mcs_rom0_30_x0x4}), .b ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_10051, new_AGEMA_signal_10050, new_AGEMA_signal_10049, mcs1_mcs_mat1_7_mcs_rom0_30_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676]}), .c ({new_AGEMA_signal_9136, new_AGEMA_signal_9135, new_AGEMA_signal_9134, mcs1_mcs_mat1_7_mcs_rom0_30_x0x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U10 ( .a ({new_AGEMA_signal_12799, new_AGEMA_signal_12798, new_AGEMA_signal_12797, mcs1_mcs_mat1_7_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_9139, new_AGEMA_signal_9138, new_AGEMA_signal_9137, mcs1_mcs_mat1_7_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_14242, new_AGEMA_signal_14241, new_AGEMA_signal_14240, mcs1_mcs_mat1_7_mcs_out[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U6 ( .a ({new_AGEMA_signal_12799, new_AGEMA_signal_12798, new_AGEMA_signal_12797, mcs1_mcs_mat1_7_mcs_rom0_31_n12}), .b ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .c ({new_AGEMA_signal_14248, new_AGEMA_signal_14247, new_AGEMA_signal_14246, mcs1_mcs_mat1_7_mcs_rom0_31_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U5 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_11350, new_AGEMA_signal_11349, new_AGEMA_signal_11348, mcs1_mcs_mat1_7_mcs_rom0_31_n11}), .c ({new_AGEMA_signal_12799, new_AGEMA_signal_12798, new_AGEMA_signal_12797, mcs1_mcs_mat1_7_mcs_rom0_31_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U4 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_11350, new_AGEMA_signal_11349, new_AGEMA_signal_11348, mcs1_mcs_mat1_7_mcs_rom0_31_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U2 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .c ({new_AGEMA_signal_12802, new_AGEMA_signal_12801, new_AGEMA_signal_12800, mcs1_mcs_mat1_7_mcs_rom0_31_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x0x4_AND_U1 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682]}), .c ({new_AGEMA_signal_9139, new_AGEMA_signal_9138, new_AGEMA_signal_9137, mcs1_mcs_mat1_7_mcs_rom0_31_x0x4}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(3), .pipeline(0)) U515 ( .a ({new_AGEMA_signal_21346, new_AGEMA_signal_21345, new_AGEMA_signal_21344, mcs_out[128]}), .b ({w0_s3[0], w0_s2[0], w0_s1[0], w0_s0[0]}), .c ({new_AGEMA_signal_21406, new_AGEMA_signal_21405, new_AGEMA_signal_21404, y0_1[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U516 ( .a ({new_AGEMA_signal_19915, new_AGEMA_signal_19914, new_AGEMA_signal_19913, mcs_out[228]}), .b ({w0_s3[100], w0_s2[100], w0_s1[100], w0_s0[100]}), .c ({new_AGEMA_signal_20080, new_AGEMA_signal_20079, new_AGEMA_signal_20078, y0_1[100]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U517 ( .a ({new_AGEMA_signal_20686, new_AGEMA_signal_20685, new_AGEMA_signal_20684, mcs_out[229]}), .b ({w0_s3[101], w0_s2[101], w0_s1[101], w0_s0[101]}), .c ({new_AGEMA_signal_20830, new_AGEMA_signal_20829, new_AGEMA_signal_20828, y0_1[101]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U518 ( .a ({new_AGEMA_signal_21310, new_AGEMA_signal_21309, new_AGEMA_signal_21308, mcs_out[230]}), .b ({w0_s3[102], w0_s2[102], w0_s1[102], w0_s0[102]}), .c ({new_AGEMA_signal_21409, new_AGEMA_signal_21408, new_AGEMA_signal_21407, y0_1[102]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U519 ( .a ({new_AGEMA_signal_21307, new_AGEMA_signal_21306, new_AGEMA_signal_21305, mcs_out[231]}), .b ({w0_s3[103], w0_s2[103], w0_s1[103], w0_s0[103]}), .c ({new_AGEMA_signal_21412, new_AGEMA_signal_21411, new_AGEMA_signal_21410, y0_1[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U520 ( .a ({new_AGEMA_signal_21283, new_AGEMA_signal_21282, new_AGEMA_signal_21281, mcs_out[232]}), .b ({w0_s3[104], w0_s2[104], w0_s1[104], w0_s0[104]}), .c ({new_AGEMA_signal_21415, new_AGEMA_signal_21414, new_AGEMA_signal_21413, y0_1[104]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U521 ( .a ({new_AGEMA_signal_19126, new_AGEMA_signal_19125, new_AGEMA_signal_19124, mcs_out[233]}), .b ({w0_s3[105], w0_s2[105], w0_s1[105], w0_s0[105]}), .c ({new_AGEMA_signal_19372, new_AGEMA_signal_19371, new_AGEMA_signal_19370, y0_1[105]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U522 ( .a ({new_AGEMA_signal_19840, new_AGEMA_signal_19839, new_AGEMA_signal_19838, mcs_out[234]}), .b ({w0_s3[106], w0_s2[106], w0_s1[106], w0_s0[106]}), .c ({new_AGEMA_signal_20083, new_AGEMA_signal_20082, new_AGEMA_signal_20081, y0_1[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U523 ( .a ({new_AGEMA_signal_20632, new_AGEMA_signal_20631, new_AGEMA_signal_20630, mcs_out[235]}), .b ({w0_s3[107], w0_s2[107], w0_s1[107], w0_s0[107]}), .c ({new_AGEMA_signal_20833, new_AGEMA_signal_20832, new_AGEMA_signal_20831, y0_1[107]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U524 ( .a ({new_AGEMA_signal_17731, new_AGEMA_signal_17730, new_AGEMA_signal_17729, mcs_out[236]}), .b ({w0_s3[108], w0_s2[108], w0_s1[108], w0_s0[108]}), .c ({new_AGEMA_signal_18052, new_AGEMA_signal_18051, new_AGEMA_signal_18050, y0_1[108]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U525 ( .a ({new_AGEMA_signal_18403, new_AGEMA_signal_18402, new_AGEMA_signal_18401, mcs_out[237]}), .b ({w0_s3[109], w0_s2[109], w0_s1[109], w0_s0[109]}), .c ({new_AGEMA_signal_18676, new_AGEMA_signal_18675, new_AGEMA_signal_18674, y0_1[109]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U526 ( .a ({new_AGEMA_signal_20650, new_AGEMA_signal_20649, new_AGEMA_signal_20648, mcs_out[138]}), .b ({w0_s3[10], w0_s2[10], w0_s1[10], w0_s0[10]}), .c ({new_AGEMA_signal_20836, new_AGEMA_signal_20835, new_AGEMA_signal_20834, y0_1[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U527 ( .a ({new_AGEMA_signal_18400, new_AGEMA_signal_18399, new_AGEMA_signal_18398, mcs_out[238]}), .b ({w0_s3[110], w0_s2[110], w0_s1[110], w0_s0[110]}), .c ({new_AGEMA_signal_18679, new_AGEMA_signal_18678, new_AGEMA_signal_18677, y0_1[110]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U528 ( .a ({new_AGEMA_signal_17722, new_AGEMA_signal_17721, new_AGEMA_signal_17720, mcs_out[239]}), .b ({w0_s3[111], w0_s2[111], w0_s1[111], w0_s0[111]}), .c ({new_AGEMA_signal_18055, new_AGEMA_signal_18054, new_AGEMA_signal_18053, y0_1[111]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U529 ( .a ({new_AGEMA_signal_20536, new_AGEMA_signal_20535, new_AGEMA_signal_20534, mcs_out[240]}), .b ({w0_s3[112], w0_s2[112], w0_s1[112], w0_s0[112]}), .c ({new_AGEMA_signal_20839, new_AGEMA_signal_20838, new_AGEMA_signal_20837, y0_1[112]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U530 ( .a ({new_AGEMA_signal_21226, new_AGEMA_signal_21225, new_AGEMA_signal_21224, mcs_out[241]}), .b ({w0_s3[113], w0_s2[113], w0_s1[113], w0_s0[113]}), .c ({new_AGEMA_signal_21418, new_AGEMA_signal_21417, new_AGEMA_signal_21416, y0_1[113]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U531 ( .a ({new_AGEMA_signal_18973, new_AGEMA_signal_18972, new_AGEMA_signal_18971, mcs_out[242]}), .b ({w0_s3[114], w0_s2[114], w0_s1[114], w0_s0[114]}), .c ({new_AGEMA_signal_19375, new_AGEMA_signal_19374, new_AGEMA_signal_19373, y0_1[114]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U532 ( .a ({new_AGEMA_signal_21223, new_AGEMA_signal_21222, new_AGEMA_signal_21221, mcs_out[243]}), .b ({w0_s3[115], w0_s2[115], w0_s1[115], w0_s0[115]}), .c ({new_AGEMA_signal_21421, new_AGEMA_signal_21420, new_AGEMA_signal_21419, y0_1[115]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U533 ( .a ({new_AGEMA_signal_19630, new_AGEMA_signal_19629, new_AGEMA_signal_19628, mcs_out[244]}), .b ({w0_s3[116], w0_s2[116], w0_s1[116], w0_s0[116]}), .c ({new_AGEMA_signal_20086, new_AGEMA_signal_20085, new_AGEMA_signal_20084, y0_1[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U534 ( .a ({new_AGEMA_signal_20479, new_AGEMA_signal_20478, new_AGEMA_signal_20477, mcs_out[245]}), .b ({w0_s3[117], w0_s2[117], w0_s1[117], w0_s0[117]}), .c ({new_AGEMA_signal_20842, new_AGEMA_signal_20841, new_AGEMA_signal_20840, y0_1[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U535 ( .a ({new_AGEMA_signal_21199, new_AGEMA_signal_21198, new_AGEMA_signal_21197, mcs_out[246]}), .b ({w0_s3[118], w0_s2[118], w0_s1[118], w0_s0[118]}), .c ({new_AGEMA_signal_21424, new_AGEMA_signal_21423, new_AGEMA_signal_21422, y0_1[118]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U536 ( .a ({new_AGEMA_signal_21196, new_AGEMA_signal_21195, new_AGEMA_signal_21194, mcs_out[247]}), .b ({w0_s3[119], w0_s2[119], w0_s1[119], w0_s0[119]}), .c ({new_AGEMA_signal_21427, new_AGEMA_signal_21426, new_AGEMA_signal_21425, y0_1[119]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U537 ( .a ({new_AGEMA_signal_21289, new_AGEMA_signal_21288, new_AGEMA_signal_21287, mcs_out[139]}), .b ({w0_s3[11], w0_s2[11], w0_s1[11], w0_s0[11]}), .c ({new_AGEMA_signal_21430, new_AGEMA_signal_21429, new_AGEMA_signal_21428, y0_1[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U538 ( .a ({new_AGEMA_signal_21172, new_AGEMA_signal_21171, new_AGEMA_signal_21170, mcs_out[248]}), .b ({w0_s3[120], w0_s2[120], w0_s1[120], w0_s0[120]}), .c ({new_AGEMA_signal_21433, new_AGEMA_signal_21432, new_AGEMA_signal_21431, y0_1[120]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U539 ( .a ({new_AGEMA_signal_18829, new_AGEMA_signal_18828, new_AGEMA_signal_18827, mcs_out[249]}), .b ({w0_s3[121], w0_s2[121], w0_s1[121], w0_s0[121]}), .c ({new_AGEMA_signal_19378, new_AGEMA_signal_19377, new_AGEMA_signal_19376, y0_1[121]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U540 ( .a ({new_AGEMA_signal_19555, new_AGEMA_signal_19554, new_AGEMA_signal_19553, mcs_out[250]}), .b ({w0_s3[122], w0_s2[122], w0_s1[122], w0_s0[122]}), .c ({new_AGEMA_signal_20089, new_AGEMA_signal_20088, new_AGEMA_signal_20087, y0_1[122]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U541 ( .a ({new_AGEMA_signal_20425, new_AGEMA_signal_20424, new_AGEMA_signal_20423, mcs_out[251]}), .b ({w0_s3[123], w0_s2[123], w0_s1[123], w0_s0[123]}), .c ({new_AGEMA_signal_20845, new_AGEMA_signal_20844, new_AGEMA_signal_20843, y0_1[123]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U542 ( .a ({new_AGEMA_signal_17404, new_AGEMA_signal_17403, new_AGEMA_signal_17402, mcs_out[252]}), .b ({w0_s3[124], w0_s2[124], w0_s1[124], w0_s0[124]}), .c ({new_AGEMA_signal_18058, new_AGEMA_signal_18057, new_AGEMA_signal_18056, y0_1[124]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U543 ( .a ({new_AGEMA_signal_18124, new_AGEMA_signal_18123, new_AGEMA_signal_18122, mcs_out[253]}), .b ({w0_s3[125], w0_s2[125], w0_s1[125], w0_s0[125]}), .c ({new_AGEMA_signal_18682, new_AGEMA_signal_18681, new_AGEMA_signal_18680, y0_1[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U544 ( .a ({new_AGEMA_signal_18121, new_AGEMA_signal_18120, new_AGEMA_signal_18119, mcs_out[254]}), .b ({w0_s3[126], w0_s2[126], w0_s1[126], w0_s0[126]}), .c ({new_AGEMA_signal_18685, new_AGEMA_signal_18684, new_AGEMA_signal_18683, y0_1[126]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U545 ( .a ({new_AGEMA_signal_17395, new_AGEMA_signal_17394, new_AGEMA_signal_17393, mcs_out[255]}), .b ({w0_s3[127], w0_s2[127], w0_s1[127], w0_s0[127]}), .c ({new_AGEMA_signal_18061, new_AGEMA_signal_18060, new_AGEMA_signal_18059, y0_1[127]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U546 ( .a ({new_AGEMA_signal_21268, new_AGEMA_signal_21267, new_AGEMA_signal_21266, mcs_out[140]}), .b ({w0_s3[12], w0_s2[12], w0_s1[12], w0_s0[12]}), .c ({new_AGEMA_signal_21436, new_AGEMA_signal_21435, new_AGEMA_signal_21434, y0_1[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U547 ( .a ({new_AGEMA_signal_19057, new_AGEMA_signal_19056, new_AGEMA_signal_19055, mcs_out[141]}), .b ({w0_s3[13], w0_s2[13], w0_s1[13], w0_s0[13]}), .c ({new_AGEMA_signal_19381, new_AGEMA_signal_19380, new_AGEMA_signal_19379, y0_1[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U548 ( .a ({new_AGEMA_signal_17734, new_AGEMA_signal_17733, new_AGEMA_signal_17732, mcs_out[142]}), .b ({w0_s3[14], w0_s2[14], w0_s1[14], w0_s0[14]}), .c ({new_AGEMA_signal_18064, new_AGEMA_signal_18063, new_AGEMA_signal_18062, y0_1[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U549 ( .a ({new_AGEMA_signal_20605, new_AGEMA_signal_20604, new_AGEMA_signal_20603, mcs_out[143]}), .b ({w0_s3[15], w0_s2[15], w0_s1[15], w0_s0[15]}), .c ({new_AGEMA_signal_20848, new_AGEMA_signal_20847, new_AGEMA_signal_20846, y0_1[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U550 ( .a ({new_AGEMA_signal_21235, new_AGEMA_signal_21234, new_AGEMA_signal_21233, mcs_out[144]}), .b ({w0_s3[16], w0_s2[16], w0_s1[16], w0_s0[16]}), .c ({new_AGEMA_signal_21439, new_AGEMA_signal_21438, new_AGEMA_signal_21437, y0_1[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U551 ( .a ({new_AGEMA_signal_19720, new_AGEMA_signal_19719, new_AGEMA_signal_19718, mcs_out[145]}), .b ({w0_s3[17], w0_s2[17], w0_s1[17], w0_s0[17]}), .c ({new_AGEMA_signal_20092, new_AGEMA_signal_20091, new_AGEMA_signal_20090, y0_1[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U552 ( .a ({new_AGEMA_signal_21232, new_AGEMA_signal_21231, new_AGEMA_signal_21230, mcs_out[146]}), .b ({w0_s3[18], w0_s2[18], w0_s1[18], w0_s0[18]}), .c ({new_AGEMA_signal_21442, new_AGEMA_signal_21441, new_AGEMA_signal_21440, y0_1[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U553 ( .a ({new_AGEMA_signal_18979, new_AGEMA_signal_18978, new_AGEMA_signal_18977, mcs_out[147]}), .b ({w0_s3[19], w0_s2[19], w0_s1[19], w0_s0[19]}), .c ({new_AGEMA_signal_19384, new_AGEMA_signal_19383, new_AGEMA_signal_19382, y0_1[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U554 ( .a ({new_AGEMA_signal_20005, new_AGEMA_signal_20004, new_AGEMA_signal_20003, mcs_out[129]}), .b ({w0_s3[1], w0_s2[1], w0_s1[1], w0_s0[1]}), .c ({new_AGEMA_signal_20095, new_AGEMA_signal_20094, new_AGEMA_signal_20093, y0_1[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U555 ( .a ({new_AGEMA_signal_20497, new_AGEMA_signal_20496, new_AGEMA_signal_20495, mcs_out[148]}), .b ({w0_s3[20], w0_s2[20], w0_s1[20], w0_s0[20]}), .c ({new_AGEMA_signal_20851, new_AGEMA_signal_20850, new_AGEMA_signal_20849, y0_1[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U556 ( .a ({new_AGEMA_signal_21205, new_AGEMA_signal_21204, new_AGEMA_signal_21203, mcs_out[149]}), .b ({w0_s3[21], w0_s2[21], w0_s1[21], w0_s0[21]}), .c ({new_AGEMA_signal_21445, new_AGEMA_signal_21444, new_AGEMA_signal_21443, y0_1[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U557 ( .a ({new_AGEMA_signal_21202, new_AGEMA_signal_21201, new_AGEMA_signal_21200, mcs_out[150]}), .b ({w0_s3[22], w0_s2[22], w0_s1[22], w0_s0[22]}), .c ({new_AGEMA_signal_21448, new_AGEMA_signal_21447, new_AGEMA_signal_21446, y0_1[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U558 ( .a ({new_AGEMA_signal_20488, new_AGEMA_signal_20487, new_AGEMA_signal_20486, mcs_out[151]}), .b ({w0_s3[23], w0_s2[23], w0_s1[23], w0_s0[23]}), .c ({new_AGEMA_signal_20854, new_AGEMA_signal_20853, new_AGEMA_signal_20852, y0_1[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U559 ( .a ({new_AGEMA_signal_21682, new_AGEMA_signal_21681, new_AGEMA_signal_21680, mcs_out[152]}), .b ({w0_s3[24], w0_s2[24], w0_s1[24], w0_s0[24]}), .c ({new_AGEMA_signal_21790, new_AGEMA_signal_21789, new_AGEMA_signal_21788, y0_1[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U560 ( .a ({new_AGEMA_signal_18844, new_AGEMA_signal_18843, new_AGEMA_signal_18842, mcs_out[153]}), .b ({w0_s3[25], w0_s2[25], w0_s1[25], w0_s0[25]}), .c ({new_AGEMA_signal_19387, new_AGEMA_signal_19386, new_AGEMA_signal_19385, y0_1[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U561 ( .a ({new_AGEMA_signal_20443, new_AGEMA_signal_20442, new_AGEMA_signal_20441, mcs_out[154]}), .b ({w0_s3[26], w0_s2[26], w0_s1[26], w0_s0[26]}), .c ({new_AGEMA_signal_20857, new_AGEMA_signal_20856, new_AGEMA_signal_20855, y0_1[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U562 ( .a ({new_AGEMA_signal_21178, new_AGEMA_signal_21177, new_AGEMA_signal_21176, mcs_out[155]}), .b ({w0_s3[27], w0_s2[27], w0_s1[27], w0_s0[27]}), .c ({new_AGEMA_signal_21451, new_AGEMA_signal_21450, new_AGEMA_signal_21449, y0_1[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U563 ( .a ({new_AGEMA_signal_21157, new_AGEMA_signal_21156, new_AGEMA_signal_21155, mcs_out[156]}), .b ({w0_s3[28], w0_s2[28], w0_s1[28], w0_s0[28]}), .c ({new_AGEMA_signal_21454, new_AGEMA_signal_21453, new_AGEMA_signal_21452, y0_1[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U564 ( .a ({new_AGEMA_signal_18760, new_AGEMA_signal_18759, new_AGEMA_signal_18758, mcs_out[157]}), .b ({w0_s3[29], w0_s2[29], w0_s1[29], w0_s0[29]}), .c ({new_AGEMA_signal_19390, new_AGEMA_signal_19389, new_AGEMA_signal_19388, y0_1[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U565 ( .a ({new_AGEMA_signal_21343, new_AGEMA_signal_21342, new_AGEMA_signal_21341, mcs_out[130]}), .b ({w0_s3[2], w0_s2[2], w0_s1[2], w0_s0[2]}), .c ({new_AGEMA_signal_21457, new_AGEMA_signal_21456, new_AGEMA_signal_21455, y0_1[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U566 ( .a ({new_AGEMA_signal_17407, new_AGEMA_signal_17406, new_AGEMA_signal_17405, mcs_out[158]}), .b ({w0_s3[30], w0_s2[30], w0_s1[30], w0_s0[30]}), .c ({new_AGEMA_signal_18067, new_AGEMA_signal_18066, new_AGEMA_signal_18065, y0_1[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U567 ( .a ({new_AGEMA_signal_20398, new_AGEMA_signal_20397, new_AGEMA_signal_20396, mcs_out[159]}), .b ({w0_s3[31], w0_s2[31], w0_s1[31], w0_s0[31]}), .c ({new_AGEMA_signal_20860, new_AGEMA_signal_20859, new_AGEMA_signal_20858, y0_1[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U568 ( .a ({new_AGEMA_signal_17974, new_AGEMA_signal_17973, new_AGEMA_signal_17972, mcs_out[160]}), .b ({w0_s3[32], w0_s2[32], w0_s1[32], w0_s0[32]}), .c ({new_AGEMA_signal_18070, new_AGEMA_signal_18069, new_AGEMA_signal_18068, y0_1[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U569 ( .a ({new_AGEMA_signal_18613, new_AGEMA_signal_18612, new_AGEMA_signal_18611, mcs_out[161]}), .b ({w0_s3[33], w0_s2[33], w0_s1[33], w0_s0[33]}), .c ({new_AGEMA_signal_18688, new_AGEMA_signal_18687, new_AGEMA_signal_18686, y0_1[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U570 ( .a ({new_AGEMA_signal_18610, new_AGEMA_signal_18609, new_AGEMA_signal_18608, mcs_out[162]}), .b ({w0_s3[34], w0_s2[34], w0_s1[34], w0_s0[34]}), .c ({new_AGEMA_signal_18691, new_AGEMA_signal_18690, new_AGEMA_signal_18689, y0_1[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U571 ( .a ({new_AGEMA_signal_18607, new_AGEMA_signal_18606, new_AGEMA_signal_18605, mcs_out[163]}), .b ({w0_s3[35], w0_s2[35], w0_s1[35], w0_s0[35]}), .c ({new_AGEMA_signal_18694, new_AGEMA_signal_18693, new_AGEMA_signal_18692, y0_1[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U572 ( .a ({new_AGEMA_signal_19927, new_AGEMA_signal_19926, new_AGEMA_signal_19925, mcs_out[164]}), .b ({w0_s3[36], w0_s2[36], w0_s1[36], w0_s0[36]}), .c ({new_AGEMA_signal_20098, new_AGEMA_signal_20097, new_AGEMA_signal_20096, y0_1[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U573 ( .a ({new_AGEMA_signal_17881, new_AGEMA_signal_17880, new_AGEMA_signal_17879, mcs_out[165]}), .b ({w0_s3[37], w0_s2[37], w0_s1[37], w0_s0[37]}), .c ({new_AGEMA_signal_18073, new_AGEMA_signal_18072, new_AGEMA_signal_18071, y0_1[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U574 ( .a ({new_AGEMA_signal_16396, new_AGEMA_signal_16395, new_AGEMA_signal_16394, mcs_out[166]}), .b ({w0_s3[38], w0_s2[38], w0_s1[38], w0_s0[38]}), .c ({new_AGEMA_signal_16600, new_AGEMA_signal_16599, new_AGEMA_signal_16598, y0_1[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U575 ( .a ({new_AGEMA_signal_19207, new_AGEMA_signal_19206, new_AGEMA_signal_19205, mcs_out[167]}), .b ({w0_s3[39], w0_s2[39], w0_s1[39], w0_s0[39]}), .c ({new_AGEMA_signal_19393, new_AGEMA_signal_19392, new_AGEMA_signal_19391, y0_1[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U576 ( .a ({new_AGEMA_signal_19276, new_AGEMA_signal_19275, new_AGEMA_signal_19274, mcs_out[131]}), .b ({w0_s3[3], w0_s2[3], w0_s1[3], w0_s0[3]}), .c ({new_AGEMA_signal_19396, new_AGEMA_signal_19395, new_AGEMA_signal_19394, y0_1[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U577 ( .a ({new_AGEMA_signal_20641, new_AGEMA_signal_20640, new_AGEMA_signal_20639, mcs_out[168]}), .b ({w0_s3[40], w0_s2[40], w0_s1[40], w0_s0[40]}), .c ({new_AGEMA_signal_20863, new_AGEMA_signal_20862, new_AGEMA_signal_20861, y0_1[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U578 ( .a ({new_AGEMA_signal_19855, new_AGEMA_signal_19854, new_AGEMA_signal_19853, mcs_out[169]}), .b ({w0_s3[41], w0_s2[41], w0_s1[41], w0_s0[41]}), .c ({new_AGEMA_signal_20101, new_AGEMA_signal_20100, new_AGEMA_signal_20099, y0_1[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U579 ( .a ({new_AGEMA_signal_19852, new_AGEMA_signal_19851, new_AGEMA_signal_19850, mcs_out[170]}), .b ({w0_s3[42], w0_s2[42], w0_s1[42], w0_s0[42]}), .c ({new_AGEMA_signal_20104, new_AGEMA_signal_20103, new_AGEMA_signal_20102, y0_1[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U580 ( .a ({new_AGEMA_signal_19849, new_AGEMA_signal_19848, new_AGEMA_signal_19847, mcs_out[171]}), .b ({w0_s3[43], w0_s2[43], w0_s1[43], w0_s0[43]}), .c ({new_AGEMA_signal_20107, new_AGEMA_signal_20106, new_AGEMA_signal_20105, y0_1[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U581 ( .a ({new_AGEMA_signal_21265, new_AGEMA_signal_21264, new_AGEMA_signal_21263, mcs_out[172]}), .b ({w0_s3[44], w0_s2[44], w0_s1[44], w0_s0[44]}), .c ({new_AGEMA_signal_21460, new_AGEMA_signal_21459, new_AGEMA_signal_21458, y0_1[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U582 ( .a ({new_AGEMA_signal_19054, new_AGEMA_signal_19053, new_AGEMA_signal_19052, mcs_out[173]}), .b ({w0_s3[45], w0_s2[45], w0_s1[45], w0_s0[45]}), .c ({new_AGEMA_signal_19399, new_AGEMA_signal_19398, new_AGEMA_signal_19397, y0_1[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U583 ( .a ({new_AGEMA_signal_19051, new_AGEMA_signal_19050, new_AGEMA_signal_19049, mcs_out[174]}), .b ({w0_s3[46], w0_s2[46], w0_s1[46], w0_s0[46]}), .c ({new_AGEMA_signal_19402, new_AGEMA_signal_19401, new_AGEMA_signal_19400, y0_1[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U584 ( .a ({new_AGEMA_signal_20596, new_AGEMA_signal_20595, new_AGEMA_signal_20594, mcs_out[175]}), .b ({w0_s3[47], w0_s2[47], w0_s1[47], w0_s0[47]}), .c ({new_AGEMA_signal_20866, new_AGEMA_signal_20865, new_AGEMA_signal_20864, y0_1[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U585 ( .a ({new_AGEMA_signal_17647, new_AGEMA_signal_17646, new_AGEMA_signal_17645, mcs_out[176]}), .b ({w0_s3[48], w0_s2[48], w0_s1[48], w0_s0[48]}), .c ({new_AGEMA_signal_18076, new_AGEMA_signal_18075, new_AGEMA_signal_18074, y0_1[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U586 ( .a ({new_AGEMA_signal_18334, new_AGEMA_signal_18333, new_AGEMA_signal_18332, mcs_out[177]}), .b ({w0_s3[49], w0_s2[49], w0_s1[49], w0_s0[49]}), .c ({new_AGEMA_signal_18697, new_AGEMA_signal_18696, new_AGEMA_signal_18695, y0_1[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U587 ( .a ({new_AGEMA_signal_20704, new_AGEMA_signal_20703, new_AGEMA_signal_20702, mcs_out[132]}), .b ({w0_s3[4], w0_s2[4], w0_s1[4], w0_s0[4]}), .c ({new_AGEMA_signal_20869, new_AGEMA_signal_20868, new_AGEMA_signal_20867, y0_1[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U588 ( .a ({new_AGEMA_signal_18331, new_AGEMA_signal_18330, new_AGEMA_signal_18329, mcs_out[178]}), .b ({w0_s3[50], w0_s2[50], w0_s1[50], w0_s0[50]}), .c ({new_AGEMA_signal_18700, new_AGEMA_signal_18699, new_AGEMA_signal_18698, y0_1[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U589 ( .a ({new_AGEMA_signal_18328, new_AGEMA_signal_18327, new_AGEMA_signal_18326, mcs_out[179]}), .b ({w0_s3[51], w0_s2[51], w0_s1[51], w0_s0[51]}), .c ({new_AGEMA_signal_18703, new_AGEMA_signal_18702, new_AGEMA_signal_18701, y0_1[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U590 ( .a ({new_AGEMA_signal_19642, new_AGEMA_signal_19641, new_AGEMA_signal_19640, mcs_out[180]}), .b ({w0_s3[52], w0_s2[52], w0_s1[52], w0_s0[52]}), .c ({new_AGEMA_signal_20110, new_AGEMA_signal_20109, new_AGEMA_signal_20108, y0_1[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U591 ( .a ({new_AGEMA_signal_17554, new_AGEMA_signal_17553, new_AGEMA_signal_17552, mcs_out[181]}), .b ({w0_s3[53], w0_s2[53], w0_s1[53], w0_s0[53]}), .c ({new_AGEMA_signal_18079, new_AGEMA_signal_18078, new_AGEMA_signal_18077, y0_1[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U592 ( .a ({new_AGEMA_signal_15955, new_AGEMA_signal_15954, new_AGEMA_signal_15953, mcs_out[182]}), .b ({w0_s3[54], w0_s2[54], w0_s1[54], w0_s0[54]}), .c ({new_AGEMA_signal_16603, new_AGEMA_signal_16602, new_AGEMA_signal_16601, y0_1[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U593 ( .a ({new_AGEMA_signal_18910, new_AGEMA_signal_18909, new_AGEMA_signal_18908, mcs_out[183]}), .b ({w0_s3[55], w0_s2[55], w0_s1[55], w0_s0[55]}), .c ({new_AGEMA_signal_19405, new_AGEMA_signal_19404, new_AGEMA_signal_19403, y0_1[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U594 ( .a ({new_AGEMA_signal_20434, new_AGEMA_signal_20433, new_AGEMA_signal_20432, mcs_out[184]}), .b ({w0_s3[56], w0_s2[56], w0_s1[56], w0_s0[56]}), .c ({new_AGEMA_signal_20872, new_AGEMA_signal_20871, new_AGEMA_signal_20870, y0_1[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U595 ( .a ({new_AGEMA_signal_19570, new_AGEMA_signal_19569, new_AGEMA_signal_19568, mcs_out[185]}), .b ({w0_s3[57], w0_s2[57], w0_s1[57], w0_s0[57]}), .c ({new_AGEMA_signal_20113, new_AGEMA_signal_20112, new_AGEMA_signal_20111, y0_1[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U596 ( .a ({new_AGEMA_signal_19567, new_AGEMA_signal_19566, new_AGEMA_signal_19565, mcs_out[186]}), .b ({w0_s3[58], w0_s2[58], w0_s1[58], w0_s0[58]}), .c ({new_AGEMA_signal_20116, new_AGEMA_signal_20115, new_AGEMA_signal_20114, y0_1[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U597 ( .a ({new_AGEMA_signal_19564, new_AGEMA_signal_19563, new_AGEMA_signal_19562, mcs_out[187]}), .b ({w0_s3[59], w0_s2[59], w0_s1[59], w0_s0[59]}), .c ({new_AGEMA_signal_20119, new_AGEMA_signal_20118, new_AGEMA_signal_20117, y0_1[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U598 ( .a ({new_AGEMA_signal_21316, new_AGEMA_signal_21315, new_AGEMA_signal_21314, mcs_out[133]}), .b ({w0_s3[5], w0_s2[5], w0_s1[5], w0_s0[5]}), .c ({new_AGEMA_signal_21463, new_AGEMA_signal_21462, new_AGEMA_signal_21461, y0_1[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U599 ( .a ({new_AGEMA_signal_21154, new_AGEMA_signal_21153, new_AGEMA_signal_21152, mcs_out[188]}), .b ({w0_s3[60], w0_s2[60], w0_s1[60], w0_s0[60]}), .c ({new_AGEMA_signal_21466, new_AGEMA_signal_21465, new_AGEMA_signal_21464, y0_1[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U600 ( .a ({new_AGEMA_signal_18757, new_AGEMA_signal_18756, new_AGEMA_signal_18755, mcs_out[189]}), .b ({w0_s3[61], w0_s2[61], w0_s1[61], w0_s0[61]}), .c ({new_AGEMA_signal_19408, new_AGEMA_signal_19407, new_AGEMA_signal_19406, y0_1[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U601 ( .a ({new_AGEMA_signal_18754, new_AGEMA_signal_18753, new_AGEMA_signal_18752, mcs_out[190]}), .b ({w0_s3[62], w0_s2[62], w0_s1[62], w0_s0[62]}), .c ({new_AGEMA_signal_19411, new_AGEMA_signal_19410, new_AGEMA_signal_19409, y0_1[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U602 ( .a ({new_AGEMA_signal_20389, new_AGEMA_signal_20388, new_AGEMA_signal_20387, mcs_out[191]}), .b ({w0_s3[63], w0_s2[63], w0_s1[63], w0_s0[63]}), .c ({new_AGEMA_signal_20875, new_AGEMA_signal_20874, new_AGEMA_signal_20873, y0_1[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U603 ( .a ({new_AGEMA_signal_21340, new_AGEMA_signal_21339, new_AGEMA_signal_21338, mcs_out[192]}), .b ({w0_s3[64], w0_s2[64], w0_s1[64], w0_s0[64]}), .c ({new_AGEMA_signal_21469, new_AGEMA_signal_21468, new_AGEMA_signal_21467, y0_1[64]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U604 ( .a ({new_AGEMA_signal_20752, new_AGEMA_signal_20751, new_AGEMA_signal_20750, mcs_out[193]}), .b ({w0_s3[65], w0_s2[65], w0_s1[65], w0_s0[65]}), .c ({new_AGEMA_signal_20878, new_AGEMA_signal_20877, new_AGEMA_signal_20876, y0_1[65]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U605 ( .a ({new_AGEMA_signal_20749, new_AGEMA_signal_20748, new_AGEMA_signal_20747, mcs_out[194]}), .b ({w0_s3[66], w0_s2[66], w0_s1[66], w0_s0[66]}), .c ({new_AGEMA_signal_20881, new_AGEMA_signal_20880, new_AGEMA_signal_20879, y0_1[66]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U606 ( .a ({new_AGEMA_signal_20746, new_AGEMA_signal_20745, new_AGEMA_signal_20744, mcs_out[195]}), .b ({w0_s3[67], w0_s2[67], w0_s1[67], w0_s0[67]}), .c ({new_AGEMA_signal_20884, new_AGEMA_signal_20883, new_AGEMA_signal_20882, y0_1[67]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U607 ( .a ({new_AGEMA_signal_20692, new_AGEMA_signal_20691, new_AGEMA_signal_20690, mcs_out[196]}), .b ({w0_s3[68], w0_s2[68], w0_s1[68], w0_s0[68]}), .c ({new_AGEMA_signal_20887, new_AGEMA_signal_20886, new_AGEMA_signal_20885, y0_1[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U608 ( .a ({new_AGEMA_signal_19921, new_AGEMA_signal_19920, new_AGEMA_signal_19919, mcs_out[197]}), .b ({w0_s3[69], w0_s2[69], w0_s1[69], w0_s0[69]}), .c ({new_AGEMA_signal_20122, new_AGEMA_signal_20121, new_AGEMA_signal_20120, y0_1[69]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U609 ( .a ({new_AGEMA_signal_21313, new_AGEMA_signal_21312, new_AGEMA_signal_21311, mcs_out[134]}), .b ({w0_s3[6], w0_s2[6], w0_s1[6], w0_s0[6]}), .c ({new_AGEMA_signal_21472, new_AGEMA_signal_21471, new_AGEMA_signal_21470, y0_1[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U610 ( .a ({new_AGEMA_signal_19201, new_AGEMA_signal_19200, new_AGEMA_signal_19199, mcs_out[198]}), .b ({w0_s3[70], w0_s2[70], w0_s1[70], w0_s0[70]}), .c ({new_AGEMA_signal_19414, new_AGEMA_signal_19413, new_AGEMA_signal_19412, y0_1[70]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U611 ( .a ({new_AGEMA_signal_20689, new_AGEMA_signal_20688, new_AGEMA_signal_20687, mcs_out[199]}), .b ({w0_s3[71], w0_s2[71], w0_s1[71], w0_s0[71]}), .c ({new_AGEMA_signal_20890, new_AGEMA_signal_20889, new_AGEMA_signal_20888, y0_1[71]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U612 ( .a ({new_AGEMA_signal_21838, new_AGEMA_signal_21837, new_AGEMA_signal_21836, mcs_out[200]}), .b ({w0_s3[72], w0_s2[72], w0_s1[72], w0_s0[72]}), .c ({new_AGEMA_signal_21952, new_AGEMA_signal_21951, new_AGEMA_signal_21950, y0_1[72]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U613 ( .a ({new_AGEMA_signal_18466, new_AGEMA_signal_18465, new_AGEMA_signal_18464, mcs_out[201]}), .b ({w0_s3[73], w0_s2[73], w0_s1[73], w0_s0[73]}), .c ({new_AGEMA_signal_18706, new_AGEMA_signal_18705, new_AGEMA_signal_18704, y0_1[73]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U614 ( .a ({new_AGEMA_signal_19846, new_AGEMA_signal_19845, new_AGEMA_signal_19844, mcs_out[202]}), .b ({w0_s3[74], w0_s2[74], w0_s1[74], w0_s0[74]}), .c ({new_AGEMA_signal_20125, new_AGEMA_signal_20124, new_AGEMA_signal_20123, y0_1[74]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U615 ( .a ({new_AGEMA_signal_21286, new_AGEMA_signal_21285, new_AGEMA_signal_21284, mcs_out[203]}), .b ({w0_s3[75], w0_s2[75], w0_s1[75], w0_s0[75]}), .c ({new_AGEMA_signal_21475, new_AGEMA_signal_21474, new_AGEMA_signal_21473, y0_1[75]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U616 ( .a ({new_AGEMA_signal_21262, new_AGEMA_signal_21261, new_AGEMA_signal_21260, mcs_out[204]}), .b ({w0_s3[76], w0_s2[76], w0_s1[76], w0_s0[76]}), .c ({new_AGEMA_signal_21478, new_AGEMA_signal_21477, new_AGEMA_signal_21476, y0_1[76]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U617 ( .a ({new_AGEMA_signal_21259, new_AGEMA_signal_21258, new_AGEMA_signal_21257, mcs_out[205]}), .b ({w0_s3[77], w0_s2[77], w0_s1[77], w0_s0[77]}), .c ({new_AGEMA_signal_21481, new_AGEMA_signal_21480, new_AGEMA_signal_21479, y0_1[77]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U618 ( .a ({new_AGEMA_signal_21256, new_AGEMA_signal_21255, new_AGEMA_signal_21254, mcs_out[206]}), .b ({w0_s3[78], w0_s2[78], w0_s1[78], w0_s0[78]}), .c ({new_AGEMA_signal_21484, new_AGEMA_signal_21483, new_AGEMA_signal_21482, y0_1[78]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U619 ( .a ({new_AGEMA_signal_21253, new_AGEMA_signal_21252, new_AGEMA_signal_21251, mcs_out[207]}), .b ({w0_s3[79], w0_s2[79], w0_s1[79], w0_s0[79]}), .c ({new_AGEMA_signal_21487, new_AGEMA_signal_21486, new_AGEMA_signal_21485, y0_1[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U620 ( .a ({new_AGEMA_signal_20695, new_AGEMA_signal_20694, new_AGEMA_signal_20693, mcs_out[135]}), .b ({w0_s3[7], w0_s2[7], w0_s1[7], w0_s0[7]}), .c ({new_AGEMA_signal_20893, new_AGEMA_signal_20892, new_AGEMA_signal_20891, y0_1[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U621 ( .a ({new_AGEMA_signal_21229, new_AGEMA_signal_21228, new_AGEMA_signal_21227, mcs_out[208]}), .b ({w0_s3[80], w0_s2[80], w0_s1[80], w0_s0[80]}), .c ({new_AGEMA_signal_21490, new_AGEMA_signal_21489, new_AGEMA_signal_21488, y0_1[80]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U622 ( .a ({new_AGEMA_signal_20545, new_AGEMA_signal_20544, new_AGEMA_signal_20543, mcs_out[209]}), .b ({w0_s3[81], w0_s2[81], w0_s1[81], w0_s0[81]}), .c ({new_AGEMA_signal_20896, new_AGEMA_signal_20895, new_AGEMA_signal_20894, y0_1[81]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U623 ( .a ({new_AGEMA_signal_20542, new_AGEMA_signal_20541, new_AGEMA_signal_20540, mcs_out[210]}), .b ({w0_s3[82], w0_s2[82], w0_s1[82], w0_s0[82]}), .c ({new_AGEMA_signal_20899, new_AGEMA_signal_20898, new_AGEMA_signal_20897, y0_1[82]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U624 ( .a ({new_AGEMA_signal_20539, new_AGEMA_signal_20538, new_AGEMA_signal_20537, mcs_out[211]}), .b ({w0_s3[83], w0_s2[83], w0_s1[83], w0_s0[83]}), .c ({new_AGEMA_signal_20902, new_AGEMA_signal_20901, new_AGEMA_signal_20900, y0_1[83]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U625 ( .a ({new_AGEMA_signal_20485, new_AGEMA_signal_20484, new_AGEMA_signal_20483, mcs_out[212]}), .b ({w0_s3[84], w0_s2[84], w0_s1[84], w0_s0[84]}), .c ({new_AGEMA_signal_20905, new_AGEMA_signal_20904, new_AGEMA_signal_20903, y0_1[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U626 ( .a ({new_AGEMA_signal_19636, new_AGEMA_signal_19635, new_AGEMA_signal_19634, mcs_out[213]}), .b ({w0_s3[85], w0_s2[85], w0_s1[85], w0_s0[85]}), .c ({new_AGEMA_signal_20128, new_AGEMA_signal_20127, new_AGEMA_signal_20126, y0_1[85]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U627 ( .a ({new_AGEMA_signal_18904, new_AGEMA_signal_18903, new_AGEMA_signal_18902, mcs_out[214]}), .b ({w0_s3[86], w0_s2[86], w0_s1[86], w0_s0[86]}), .c ({new_AGEMA_signal_19417, new_AGEMA_signal_19416, new_AGEMA_signal_19415, y0_1[86]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U628 ( .a ({new_AGEMA_signal_20482, new_AGEMA_signal_20481, new_AGEMA_signal_20480, mcs_out[215]}), .b ({w0_s3[87], w0_s2[87], w0_s1[87], w0_s0[87]}), .c ({new_AGEMA_signal_20908, new_AGEMA_signal_20907, new_AGEMA_signal_20906, y0_1[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U629 ( .a ({new_AGEMA_signal_21832, new_AGEMA_signal_21831, new_AGEMA_signal_21830, mcs_out[216]}), .b ({w0_s3[88], w0_s2[88], w0_s1[88], w0_s0[88]}), .c ({new_AGEMA_signal_21955, new_AGEMA_signal_21954, new_AGEMA_signal_21953, y0_1[88]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U630 ( .a ({new_AGEMA_signal_18187, new_AGEMA_signal_18186, new_AGEMA_signal_18185, mcs_out[217]}), .b ({w0_s3[89], w0_s2[89], w0_s1[89], w0_s0[89]}), .c ({new_AGEMA_signal_18709, new_AGEMA_signal_18708, new_AGEMA_signal_18707, y0_1[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U631 ( .a ({new_AGEMA_signal_21700, new_AGEMA_signal_21699, new_AGEMA_signal_21698, mcs_out[136]}), .b ({w0_s3[8], w0_s2[8], w0_s1[8], w0_s0[8]}), .c ({new_AGEMA_signal_21793, new_AGEMA_signal_21792, new_AGEMA_signal_21791, y0_1[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U632 ( .a ({new_AGEMA_signal_19561, new_AGEMA_signal_19560, new_AGEMA_signal_19559, mcs_out[218]}), .b ({w0_s3[90], w0_s2[90], w0_s1[90], w0_s0[90]}), .c ({new_AGEMA_signal_20131, new_AGEMA_signal_20130, new_AGEMA_signal_20129, y0_1[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U633 ( .a ({new_AGEMA_signal_21175, new_AGEMA_signal_21174, new_AGEMA_signal_21173, mcs_out[219]}), .b ({w0_s3[91], w0_s2[91], w0_s1[91], w0_s0[91]}), .c ({new_AGEMA_signal_21493, new_AGEMA_signal_21492, new_AGEMA_signal_21491, y0_1[91]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U634 ( .a ({new_AGEMA_signal_21151, new_AGEMA_signal_21150, new_AGEMA_signal_21149, mcs_out[220]}), .b ({w0_s3[92], w0_s2[92], w0_s1[92], w0_s0[92]}), .c ({new_AGEMA_signal_21496, new_AGEMA_signal_21495, new_AGEMA_signal_21494, y0_1[92]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U635 ( .a ({new_AGEMA_signal_21148, new_AGEMA_signal_21147, new_AGEMA_signal_21146, mcs_out[221]}), .b ({w0_s3[93], w0_s2[93], w0_s1[93], w0_s0[93]}), .c ({new_AGEMA_signal_21499, new_AGEMA_signal_21498, new_AGEMA_signal_21497, y0_1[93]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U636 ( .a ({new_AGEMA_signal_21145, new_AGEMA_signal_21144, new_AGEMA_signal_21143, mcs_out[222]}), .b ({w0_s3[94], w0_s2[94], w0_s1[94], w0_s0[94]}), .c ({new_AGEMA_signal_21502, new_AGEMA_signal_21501, new_AGEMA_signal_21500, y0_1[94]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U637 ( .a ({new_AGEMA_signal_21142, new_AGEMA_signal_21141, new_AGEMA_signal_21140, mcs_out[223]}), .b ({w0_s3[95], w0_s2[95], w0_s1[95], w0_s0[95]}), .c ({new_AGEMA_signal_21505, new_AGEMA_signal_21504, new_AGEMA_signal_21503, y0_1[95]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U638 ( .a ({new_AGEMA_signal_20743, new_AGEMA_signal_20742, new_AGEMA_signal_20741, mcs_out[224]}), .b ({w0_s3[96], w0_s2[96], w0_s1[96], w0_s0[96]}), .c ({new_AGEMA_signal_20911, new_AGEMA_signal_20910, new_AGEMA_signal_20909, y0_1[96]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U639 ( .a ({new_AGEMA_signal_21337, new_AGEMA_signal_21336, new_AGEMA_signal_21335, mcs_out[225]}), .b ({w0_s3[97], w0_s2[97], w0_s1[97], w0_s0[97]}), .c ({new_AGEMA_signal_21508, new_AGEMA_signal_21507, new_AGEMA_signal_21506, y0_1[97]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U640 ( .a ({new_AGEMA_signal_19270, new_AGEMA_signal_19269, new_AGEMA_signal_19268, mcs_out[226]}), .b ({w0_s3[98], w0_s2[98], w0_s1[98], w0_s0[98]}), .c ({new_AGEMA_signal_19420, new_AGEMA_signal_19419, new_AGEMA_signal_19418, y0_1[98]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U641 ( .a ({new_AGEMA_signal_21334, new_AGEMA_signal_21333, new_AGEMA_signal_21332, mcs_out[227]}), .b ({w0_s3[99], w0_s2[99], w0_s1[99], w0_s0[99]}), .c ({new_AGEMA_signal_21511, new_AGEMA_signal_21510, new_AGEMA_signal_21509, y0_1[99]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U642 ( .a ({new_AGEMA_signal_19141, new_AGEMA_signal_19140, new_AGEMA_signal_19139, mcs_out[137]}), .b ({w0_s3[9], w0_s2[9], w0_s1[9], w0_s0[9]}), .c ({new_AGEMA_signal_19423, new_AGEMA_signal_19422, new_AGEMA_signal_19421, y0_1[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U643 ( .a ({temp_s3[0], temp_s2[0], temp_s1[0], temp_s0[0]}), .b ({temp_next_s3[0], temp_next_s2[0], temp_next_s1[0], temp_next_s0[0]}), .c ({y1_s3[0], y1_s2[0], y1_s1[0], y1_s0[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U644 ( .a ({temp_s3[100], temp_s2[100], temp_s1[100], temp_s0[100]}), .b ({temp_next_s3[100], temp_next_s2[100], temp_next_s1[100], temp_next_s0[100]}), .c ({y1_s3[100], y1_s2[100], y1_s1[100], y1_s0[100]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U645 ( .a ({temp_s3[101], temp_s2[101], temp_s1[101], temp_s0[101]}), .b ({temp_next_s3[101], temp_next_s2[101], temp_next_s1[101], temp_next_s0[101]}), .c ({y1_s3[101], y1_s2[101], y1_s1[101], y1_s0[101]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U646 ( .a ({temp_s3[102], temp_s2[102], temp_s1[102], temp_s0[102]}), .b ({temp_next_s3[102], temp_next_s2[102], temp_next_s1[102], temp_next_s0[102]}), .c ({y1_s3[102], y1_s2[102], y1_s1[102], y1_s0[102]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U647 ( .a ({temp_s3[103], temp_s2[103], temp_s1[103], temp_s0[103]}), .b ({temp_next_s3[103], temp_next_s2[103], temp_next_s1[103], temp_next_s0[103]}), .c ({y1_s3[103], y1_s2[103], y1_s1[103], y1_s0[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U648 ( .a ({temp_s3[104], temp_s2[104], temp_s1[104], temp_s0[104]}), .b ({temp_next_s3[104], temp_next_s2[104], temp_next_s1[104], temp_next_s0[104]}), .c ({y1_s3[104], y1_s2[104], y1_s1[104], y1_s0[104]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U649 ( .a ({temp_s3[105], temp_s2[105], temp_s1[105], temp_s0[105]}), .b ({temp_next_s3[105], temp_next_s2[105], temp_next_s1[105], temp_next_s0[105]}), .c ({y1_s3[105], y1_s2[105], y1_s1[105], y1_s0[105]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U650 ( .a ({temp_s3[106], temp_s2[106], temp_s1[106], temp_s0[106]}), .b ({temp_next_s3[106], temp_next_s2[106], temp_next_s1[106], temp_next_s0[106]}), .c ({y1_s3[106], y1_s2[106], y1_s1[106], y1_s0[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U651 ( .a ({temp_s3[107], temp_s2[107], temp_s1[107], temp_s0[107]}), .b ({temp_next_s3[107], temp_next_s2[107], temp_next_s1[107], temp_next_s0[107]}), .c ({y1_s3[107], y1_s2[107], y1_s1[107], y1_s0[107]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U652 ( .a ({temp_s3[108], temp_s2[108], temp_s1[108], temp_s0[108]}), .b ({temp_next_s3[108], temp_next_s2[108], temp_next_s1[108], temp_next_s0[108]}), .c ({y1_s3[108], y1_s2[108], y1_s1[108], y1_s0[108]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U653 ( .a ({temp_s3[109], temp_s2[109], temp_s1[109], temp_s0[109]}), .b ({temp_next_s3[109], temp_next_s2[109], temp_next_s1[109], temp_next_s0[109]}), .c ({y1_s3[109], y1_s2[109], y1_s1[109], y1_s0[109]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U654 ( .a ({temp_s3[10], temp_s2[10], temp_s1[10], temp_s0[10]}), .b ({temp_next_s3[10], temp_next_s2[10], temp_next_s1[10], temp_next_s0[10]}), .c ({y1_s3[10], y1_s2[10], y1_s1[10], y1_s0[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U655 ( .a ({temp_s3[110], temp_s2[110], temp_s1[110], temp_s0[110]}), .b ({temp_next_s3[110], temp_next_s2[110], temp_next_s1[110], temp_next_s0[110]}), .c ({y1_s3[110], y1_s2[110], y1_s1[110], y1_s0[110]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U656 ( .a ({temp_s3[111], temp_s2[111], temp_s1[111], temp_s0[111]}), .b ({temp_next_s3[111], temp_next_s2[111], temp_next_s1[111], temp_next_s0[111]}), .c ({y1_s3[111], y1_s2[111], y1_s1[111], y1_s0[111]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U657 ( .a ({temp_s3[112], temp_s2[112], temp_s1[112], temp_s0[112]}), .b ({temp_next_s3[112], temp_next_s2[112], temp_next_s1[112], temp_next_s0[112]}), .c ({y1_s3[112], y1_s2[112], y1_s1[112], y1_s0[112]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U658 ( .a ({temp_s3[113], temp_s2[113], temp_s1[113], temp_s0[113]}), .b ({temp_next_s3[113], temp_next_s2[113], temp_next_s1[113], temp_next_s0[113]}), .c ({y1_s3[113], y1_s2[113], y1_s1[113], y1_s0[113]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U659 ( .a ({temp_s3[114], temp_s2[114], temp_s1[114], temp_s0[114]}), .b ({temp_next_s3[114], temp_next_s2[114], temp_next_s1[114], temp_next_s0[114]}), .c ({y1_s3[114], y1_s2[114], y1_s1[114], y1_s0[114]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U660 ( .a ({temp_s3[115], temp_s2[115], temp_s1[115], temp_s0[115]}), .b ({temp_next_s3[115], temp_next_s2[115], temp_next_s1[115], temp_next_s0[115]}), .c ({y1_s3[115], y1_s2[115], y1_s1[115], y1_s0[115]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U661 ( .a ({temp_s3[116], temp_s2[116], temp_s1[116], temp_s0[116]}), .b ({temp_next_s3[116], temp_next_s2[116], temp_next_s1[116], temp_next_s0[116]}), .c ({y1_s3[116], y1_s2[116], y1_s1[116], y1_s0[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U662 ( .a ({temp_s3[117], temp_s2[117], temp_s1[117], temp_s0[117]}), .b ({temp_next_s3[117], temp_next_s2[117], temp_next_s1[117], temp_next_s0[117]}), .c ({y1_s3[117], y1_s2[117], y1_s1[117], y1_s0[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U663 ( .a ({temp_s3[118], temp_s2[118], temp_s1[118], temp_s0[118]}), .b ({temp_next_s3[118], temp_next_s2[118], temp_next_s1[118], temp_next_s0[118]}), .c ({y1_s3[118], y1_s2[118], y1_s1[118], y1_s0[118]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U664 ( .a ({temp_s3[119], temp_s2[119], temp_s1[119], temp_s0[119]}), .b ({temp_next_s3[119], temp_next_s2[119], temp_next_s1[119], temp_next_s0[119]}), .c ({y1_s3[119], y1_s2[119], y1_s1[119], y1_s0[119]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U665 ( .a ({temp_s3[11], temp_s2[11], temp_s1[11], temp_s0[11]}), .b ({temp_next_s3[11], temp_next_s2[11], temp_next_s1[11], temp_next_s0[11]}), .c ({y1_s3[11], y1_s2[11], y1_s1[11], y1_s0[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U666 ( .a ({temp_s3[120], temp_s2[120], temp_s1[120], temp_s0[120]}), .b ({temp_next_s3[120], temp_next_s2[120], temp_next_s1[120], temp_next_s0[120]}), .c ({y1_s3[120], y1_s2[120], y1_s1[120], y1_s0[120]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U667 ( .a ({temp_s3[121], temp_s2[121], temp_s1[121], temp_s0[121]}), .b ({temp_next_s3[121], temp_next_s2[121], temp_next_s1[121], temp_next_s0[121]}), .c ({y1_s3[121], y1_s2[121], y1_s1[121], y1_s0[121]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U668 ( .a ({temp_s3[122], temp_s2[122], temp_s1[122], temp_s0[122]}), .b ({temp_next_s3[122], temp_next_s2[122], temp_next_s1[122], temp_next_s0[122]}), .c ({y1_s3[122], y1_s2[122], y1_s1[122], y1_s0[122]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U669 ( .a ({temp_s3[123], temp_s2[123], temp_s1[123], temp_s0[123]}), .b ({temp_next_s3[123], temp_next_s2[123], temp_next_s1[123], temp_next_s0[123]}), .c ({y1_s3[123], y1_s2[123], y1_s1[123], y1_s0[123]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U670 ( .a ({temp_s3[124], temp_s2[124], temp_s1[124], temp_s0[124]}), .b ({temp_next_s3[124], temp_next_s2[124], temp_next_s1[124], temp_next_s0[124]}), .c ({y1_s3[124], y1_s2[124], y1_s1[124], y1_s0[124]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U671 ( .a ({temp_s3[125], temp_s2[125], temp_s1[125], temp_s0[125]}), .b ({temp_next_s3[125], temp_next_s2[125], temp_next_s1[125], temp_next_s0[125]}), .c ({y1_s3[125], y1_s2[125], y1_s1[125], y1_s0[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U672 ( .a ({temp_s3[126], temp_s2[126], temp_s1[126], temp_s0[126]}), .b ({temp_next_s3[126], temp_next_s2[126], temp_next_s1[126], temp_next_s0[126]}), .c ({y1_s3[126], y1_s2[126], y1_s1[126], y1_s0[126]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U673 ( .a ({temp_s3[127], temp_s2[127], temp_s1[127], temp_s0[127]}), .b ({temp_next_s3[127], temp_next_s2[127], temp_next_s1[127], temp_next_s0[127]}), .c ({y1_s3[127], y1_s2[127], y1_s1[127], y1_s0[127]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U674 ( .a ({temp_s3[12], temp_s2[12], temp_s1[12], temp_s0[12]}), .b ({temp_next_s3[12], temp_next_s2[12], temp_next_s1[12], temp_next_s0[12]}), .c ({y1_s3[12], y1_s2[12], y1_s1[12], y1_s0[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U675 ( .a ({temp_s3[13], temp_s2[13], temp_s1[13], temp_s0[13]}), .b ({temp_next_s3[13], temp_next_s2[13], temp_next_s1[13], temp_next_s0[13]}), .c ({y1_s3[13], y1_s2[13], y1_s1[13], y1_s0[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U676 ( .a ({temp_s3[14], temp_s2[14], temp_s1[14], temp_s0[14]}), .b ({temp_next_s3[14], temp_next_s2[14], temp_next_s1[14], temp_next_s0[14]}), .c ({y1_s3[14], y1_s2[14], y1_s1[14], y1_s0[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U677 ( .a ({temp_s3[15], temp_s2[15], temp_s1[15], temp_s0[15]}), .b ({temp_next_s3[15], temp_next_s2[15], temp_next_s1[15], temp_next_s0[15]}), .c ({y1_s3[15], y1_s2[15], y1_s1[15], y1_s0[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U678 ( .a ({temp_s3[16], temp_s2[16], temp_s1[16], temp_s0[16]}), .b ({temp_next_s3[16], temp_next_s2[16], temp_next_s1[16], temp_next_s0[16]}), .c ({y1_s3[16], y1_s2[16], y1_s1[16], y1_s0[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U679 ( .a ({temp_s3[17], temp_s2[17], temp_s1[17], temp_s0[17]}), .b ({temp_next_s3[17], temp_next_s2[17], temp_next_s1[17], temp_next_s0[17]}), .c ({y1_s3[17], y1_s2[17], y1_s1[17], y1_s0[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U680 ( .a ({temp_s3[18], temp_s2[18], temp_s1[18], temp_s0[18]}), .b ({temp_next_s3[18], temp_next_s2[18], temp_next_s1[18], temp_next_s0[18]}), .c ({y1_s3[18], y1_s2[18], y1_s1[18], y1_s0[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U681 ( .a ({temp_s3[19], temp_s2[19], temp_s1[19], temp_s0[19]}), .b ({temp_next_s3[19], temp_next_s2[19], temp_next_s1[19], temp_next_s0[19]}), .c ({y1_s3[19], y1_s2[19], y1_s1[19], y1_s0[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U682 ( .a ({temp_s3[1], temp_s2[1], temp_s1[1], temp_s0[1]}), .b ({temp_next_s3[1], temp_next_s2[1], temp_next_s1[1], temp_next_s0[1]}), .c ({y1_s3[1], y1_s2[1], y1_s1[1], y1_s0[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U683 ( .a ({temp_s3[20], temp_s2[20], temp_s1[20], temp_s0[20]}), .b ({temp_next_s3[20], temp_next_s2[20], temp_next_s1[20], temp_next_s0[20]}), .c ({y1_s3[20], y1_s2[20], y1_s1[20], y1_s0[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U684 ( .a ({temp_s3[21], temp_s2[21], temp_s1[21], temp_s0[21]}), .b ({temp_next_s3[21], temp_next_s2[21], temp_next_s1[21], temp_next_s0[21]}), .c ({y1_s3[21], y1_s2[21], y1_s1[21], y1_s0[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U685 ( .a ({temp_s3[22], temp_s2[22], temp_s1[22], temp_s0[22]}), .b ({temp_next_s3[22], temp_next_s2[22], temp_next_s1[22], temp_next_s0[22]}), .c ({y1_s3[22], y1_s2[22], y1_s1[22], y1_s0[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U686 ( .a ({temp_s3[23], temp_s2[23], temp_s1[23], temp_s0[23]}), .b ({temp_next_s3[23], temp_next_s2[23], temp_next_s1[23], temp_next_s0[23]}), .c ({y1_s3[23], y1_s2[23], y1_s1[23], y1_s0[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U687 ( .a ({temp_s3[24], temp_s2[24], temp_s1[24], temp_s0[24]}), .b ({temp_next_s3[24], temp_next_s2[24], temp_next_s1[24], temp_next_s0[24]}), .c ({y1_s3[24], y1_s2[24], y1_s1[24], y1_s0[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U688 ( .a ({temp_s3[25], temp_s2[25], temp_s1[25], temp_s0[25]}), .b ({temp_next_s3[25], temp_next_s2[25], temp_next_s1[25], temp_next_s0[25]}), .c ({y1_s3[25], y1_s2[25], y1_s1[25], y1_s0[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U689 ( .a ({temp_s3[26], temp_s2[26], temp_s1[26], temp_s0[26]}), .b ({temp_next_s3[26], temp_next_s2[26], temp_next_s1[26], temp_next_s0[26]}), .c ({y1_s3[26], y1_s2[26], y1_s1[26], y1_s0[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U690 ( .a ({temp_s3[27], temp_s2[27], temp_s1[27], temp_s0[27]}), .b ({temp_next_s3[27], temp_next_s2[27], temp_next_s1[27], temp_next_s0[27]}), .c ({y1_s3[27], y1_s2[27], y1_s1[27], y1_s0[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U691 ( .a ({temp_s3[28], temp_s2[28], temp_s1[28], temp_s0[28]}), .b ({temp_next_s3[28], temp_next_s2[28], temp_next_s1[28], temp_next_s0[28]}), .c ({y1_s3[28], y1_s2[28], y1_s1[28], y1_s0[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U692 ( .a ({temp_s3[29], temp_s2[29], temp_s1[29], temp_s0[29]}), .b ({temp_next_s3[29], temp_next_s2[29], temp_next_s1[29], temp_next_s0[29]}), .c ({y1_s3[29], y1_s2[29], y1_s1[29], y1_s0[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U693 ( .a ({temp_s3[2], temp_s2[2], temp_s1[2], temp_s0[2]}), .b ({temp_next_s3[2], temp_next_s2[2], temp_next_s1[2], temp_next_s0[2]}), .c ({y1_s3[2], y1_s2[2], y1_s1[2], y1_s0[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U694 ( .a ({temp_s3[30], temp_s2[30], temp_s1[30], temp_s0[30]}), .b ({temp_next_s3[30], temp_next_s2[30], temp_next_s1[30], temp_next_s0[30]}), .c ({y1_s3[30], y1_s2[30], y1_s1[30], y1_s0[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U695 ( .a ({temp_s3[31], temp_s2[31], temp_s1[31], temp_s0[31]}), .b ({temp_next_s3[31], temp_next_s2[31], temp_next_s1[31], temp_next_s0[31]}), .c ({y1_s3[31], y1_s2[31], y1_s1[31], y1_s0[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U696 ( .a ({temp_s3[32], temp_s2[32], temp_s1[32], temp_s0[32]}), .b ({temp_next_s3[32], temp_next_s2[32], temp_next_s1[32], temp_next_s0[32]}), .c ({y1_s3[32], y1_s2[32], y1_s1[32], y1_s0[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U697 ( .a ({temp_s3[33], temp_s2[33], temp_s1[33], temp_s0[33]}), .b ({temp_next_s3[33], temp_next_s2[33], temp_next_s1[33], temp_next_s0[33]}), .c ({y1_s3[33], y1_s2[33], y1_s1[33], y1_s0[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U698 ( .a ({temp_s3[34], temp_s2[34], temp_s1[34], temp_s0[34]}), .b ({temp_next_s3[34], temp_next_s2[34], temp_next_s1[34], temp_next_s0[34]}), .c ({y1_s3[34], y1_s2[34], y1_s1[34], y1_s0[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U699 ( .a ({temp_s3[35], temp_s2[35], temp_s1[35], temp_s0[35]}), .b ({temp_next_s3[35], temp_next_s2[35], temp_next_s1[35], temp_next_s0[35]}), .c ({y1_s3[35], y1_s2[35], y1_s1[35], y1_s0[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U700 ( .a ({temp_s3[36], temp_s2[36], temp_s1[36], temp_s0[36]}), .b ({temp_next_s3[36], temp_next_s2[36], temp_next_s1[36], temp_next_s0[36]}), .c ({y1_s3[36], y1_s2[36], y1_s1[36], y1_s0[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U701 ( .a ({temp_s3[37], temp_s2[37], temp_s1[37], temp_s0[37]}), .b ({temp_next_s3[37], temp_next_s2[37], temp_next_s1[37], temp_next_s0[37]}), .c ({y1_s3[37], y1_s2[37], y1_s1[37], y1_s0[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U702 ( .a ({temp_s3[38], temp_s2[38], temp_s1[38], temp_s0[38]}), .b ({temp_next_s3[38], temp_next_s2[38], temp_next_s1[38], temp_next_s0[38]}), .c ({y1_s3[38], y1_s2[38], y1_s1[38], y1_s0[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U703 ( .a ({temp_s3[39], temp_s2[39], temp_s1[39], temp_s0[39]}), .b ({temp_next_s3[39], temp_next_s2[39], temp_next_s1[39], temp_next_s0[39]}), .c ({y1_s3[39], y1_s2[39], y1_s1[39], y1_s0[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U704 ( .a ({temp_s3[3], temp_s2[3], temp_s1[3], temp_s0[3]}), .b ({temp_next_s3[3], temp_next_s2[3], temp_next_s1[3], temp_next_s0[3]}), .c ({y1_s3[3], y1_s2[3], y1_s1[3], y1_s0[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U705 ( .a ({temp_s3[40], temp_s2[40], temp_s1[40], temp_s0[40]}), .b ({temp_next_s3[40], temp_next_s2[40], temp_next_s1[40], temp_next_s0[40]}), .c ({y1_s3[40], y1_s2[40], y1_s1[40], y1_s0[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U706 ( .a ({temp_s3[41], temp_s2[41], temp_s1[41], temp_s0[41]}), .b ({temp_next_s3[41], temp_next_s2[41], temp_next_s1[41], temp_next_s0[41]}), .c ({y1_s3[41], y1_s2[41], y1_s1[41], y1_s0[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U707 ( .a ({temp_s3[42], temp_s2[42], temp_s1[42], temp_s0[42]}), .b ({temp_next_s3[42], temp_next_s2[42], temp_next_s1[42], temp_next_s0[42]}), .c ({y1_s3[42], y1_s2[42], y1_s1[42], y1_s0[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U708 ( .a ({temp_s3[43], temp_s2[43], temp_s1[43], temp_s0[43]}), .b ({temp_next_s3[43], temp_next_s2[43], temp_next_s1[43], temp_next_s0[43]}), .c ({y1_s3[43], y1_s2[43], y1_s1[43], y1_s0[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U709 ( .a ({temp_s3[44], temp_s2[44], temp_s1[44], temp_s0[44]}), .b ({temp_next_s3[44], temp_next_s2[44], temp_next_s1[44], temp_next_s0[44]}), .c ({y1_s3[44], y1_s2[44], y1_s1[44], y1_s0[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U710 ( .a ({temp_s3[45], temp_s2[45], temp_s1[45], temp_s0[45]}), .b ({temp_next_s3[45], temp_next_s2[45], temp_next_s1[45], temp_next_s0[45]}), .c ({y1_s3[45], y1_s2[45], y1_s1[45], y1_s0[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U711 ( .a ({temp_s3[46], temp_s2[46], temp_s1[46], temp_s0[46]}), .b ({temp_next_s3[46], temp_next_s2[46], temp_next_s1[46], temp_next_s0[46]}), .c ({y1_s3[46], y1_s2[46], y1_s1[46], y1_s0[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U712 ( .a ({temp_s3[47], temp_s2[47], temp_s1[47], temp_s0[47]}), .b ({temp_next_s3[47], temp_next_s2[47], temp_next_s1[47], temp_next_s0[47]}), .c ({y1_s3[47], y1_s2[47], y1_s1[47], y1_s0[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U713 ( .a ({temp_s3[48], temp_s2[48], temp_s1[48], temp_s0[48]}), .b ({temp_next_s3[48], temp_next_s2[48], temp_next_s1[48], temp_next_s0[48]}), .c ({y1_s3[48], y1_s2[48], y1_s1[48], y1_s0[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U714 ( .a ({temp_s3[49], temp_s2[49], temp_s1[49], temp_s0[49]}), .b ({temp_next_s3[49], temp_next_s2[49], temp_next_s1[49], temp_next_s0[49]}), .c ({y1_s3[49], y1_s2[49], y1_s1[49], y1_s0[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U715 ( .a ({temp_s3[4], temp_s2[4], temp_s1[4], temp_s0[4]}), .b ({temp_next_s3[4], temp_next_s2[4], temp_next_s1[4], temp_next_s0[4]}), .c ({y1_s3[4], y1_s2[4], y1_s1[4], y1_s0[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U716 ( .a ({temp_s3[50], temp_s2[50], temp_s1[50], temp_s0[50]}), .b ({temp_next_s3[50], temp_next_s2[50], temp_next_s1[50], temp_next_s0[50]}), .c ({y1_s3[50], y1_s2[50], y1_s1[50], y1_s0[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U717 ( .a ({temp_s3[51], temp_s2[51], temp_s1[51], temp_s0[51]}), .b ({temp_next_s3[51], temp_next_s2[51], temp_next_s1[51], temp_next_s0[51]}), .c ({y1_s3[51], y1_s2[51], y1_s1[51], y1_s0[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U718 ( .a ({temp_s3[52], temp_s2[52], temp_s1[52], temp_s0[52]}), .b ({temp_next_s3[52], temp_next_s2[52], temp_next_s1[52], temp_next_s0[52]}), .c ({y1_s3[52], y1_s2[52], y1_s1[52], y1_s0[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U719 ( .a ({temp_s3[53], temp_s2[53], temp_s1[53], temp_s0[53]}), .b ({temp_next_s3[53], temp_next_s2[53], temp_next_s1[53], temp_next_s0[53]}), .c ({y1_s3[53], y1_s2[53], y1_s1[53], y1_s0[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U720 ( .a ({temp_s3[54], temp_s2[54], temp_s1[54], temp_s0[54]}), .b ({temp_next_s3[54], temp_next_s2[54], temp_next_s1[54], temp_next_s0[54]}), .c ({y1_s3[54], y1_s2[54], y1_s1[54], y1_s0[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U721 ( .a ({temp_s3[55], temp_s2[55], temp_s1[55], temp_s0[55]}), .b ({temp_next_s3[55], temp_next_s2[55], temp_next_s1[55], temp_next_s0[55]}), .c ({y1_s3[55], y1_s2[55], y1_s1[55], y1_s0[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U722 ( .a ({temp_s3[56], temp_s2[56], temp_s1[56], temp_s0[56]}), .b ({temp_next_s3[56], temp_next_s2[56], temp_next_s1[56], temp_next_s0[56]}), .c ({y1_s3[56], y1_s2[56], y1_s1[56], y1_s0[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U723 ( .a ({temp_s3[57], temp_s2[57], temp_s1[57], temp_s0[57]}), .b ({temp_next_s3[57], temp_next_s2[57], temp_next_s1[57], temp_next_s0[57]}), .c ({y1_s3[57], y1_s2[57], y1_s1[57], y1_s0[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U724 ( .a ({temp_s3[58], temp_s2[58], temp_s1[58], temp_s0[58]}), .b ({temp_next_s3[58], temp_next_s2[58], temp_next_s1[58], temp_next_s0[58]}), .c ({y1_s3[58], y1_s2[58], y1_s1[58], y1_s0[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U725 ( .a ({temp_s3[59], temp_s2[59], temp_s1[59], temp_s0[59]}), .b ({temp_next_s3[59], temp_next_s2[59], temp_next_s1[59], temp_next_s0[59]}), .c ({y1_s3[59], y1_s2[59], y1_s1[59], y1_s0[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U726 ( .a ({temp_s3[5], temp_s2[5], temp_s1[5], temp_s0[5]}), .b ({temp_next_s3[5], temp_next_s2[5], temp_next_s1[5], temp_next_s0[5]}), .c ({y1_s3[5], y1_s2[5], y1_s1[5], y1_s0[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U727 ( .a ({temp_s3[60], temp_s2[60], temp_s1[60], temp_s0[60]}), .b ({temp_next_s3[60], temp_next_s2[60], temp_next_s1[60], temp_next_s0[60]}), .c ({y1_s3[60], y1_s2[60], y1_s1[60], y1_s0[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U728 ( .a ({temp_s3[61], temp_s2[61], temp_s1[61], temp_s0[61]}), .b ({temp_next_s3[61], temp_next_s2[61], temp_next_s1[61], temp_next_s0[61]}), .c ({y1_s3[61], y1_s2[61], y1_s1[61], y1_s0[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U729 ( .a ({temp_s3[62], temp_s2[62], temp_s1[62], temp_s0[62]}), .b ({temp_next_s3[62], temp_next_s2[62], temp_next_s1[62], temp_next_s0[62]}), .c ({y1_s3[62], y1_s2[62], y1_s1[62], y1_s0[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U730 ( .a ({temp_s3[63], temp_s2[63], temp_s1[63], temp_s0[63]}), .b ({temp_next_s3[63], temp_next_s2[63], temp_next_s1[63], temp_next_s0[63]}), .c ({y1_s3[63], y1_s2[63], y1_s1[63], y1_s0[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U731 ( .a ({temp_s3[64], temp_s2[64], temp_s1[64], temp_s0[64]}), .b ({temp_next_s3[64], temp_next_s2[64], temp_next_s1[64], temp_next_s0[64]}), .c ({y1_s3[64], y1_s2[64], y1_s1[64], y1_s0[64]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U732 ( .a ({temp_s3[65], temp_s2[65], temp_s1[65], temp_s0[65]}), .b ({temp_next_s3[65], temp_next_s2[65], temp_next_s1[65], temp_next_s0[65]}), .c ({y1_s3[65], y1_s2[65], y1_s1[65], y1_s0[65]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U733 ( .a ({temp_s3[66], temp_s2[66], temp_s1[66], temp_s0[66]}), .b ({temp_next_s3[66], temp_next_s2[66], temp_next_s1[66], temp_next_s0[66]}), .c ({y1_s3[66], y1_s2[66], y1_s1[66], y1_s0[66]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U734 ( .a ({temp_s3[67], temp_s2[67], temp_s1[67], temp_s0[67]}), .b ({temp_next_s3[67], temp_next_s2[67], temp_next_s1[67], temp_next_s0[67]}), .c ({y1_s3[67], y1_s2[67], y1_s1[67], y1_s0[67]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U735 ( .a ({temp_s3[68], temp_s2[68], temp_s1[68], temp_s0[68]}), .b ({temp_next_s3[68], temp_next_s2[68], temp_next_s1[68], temp_next_s0[68]}), .c ({y1_s3[68], y1_s2[68], y1_s1[68], y1_s0[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U736 ( .a ({temp_s3[69], temp_s2[69], temp_s1[69], temp_s0[69]}), .b ({temp_next_s3[69], temp_next_s2[69], temp_next_s1[69], temp_next_s0[69]}), .c ({y1_s3[69], y1_s2[69], y1_s1[69], y1_s0[69]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U737 ( .a ({temp_s3[6], temp_s2[6], temp_s1[6], temp_s0[6]}), .b ({temp_next_s3[6], temp_next_s2[6], temp_next_s1[6], temp_next_s0[6]}), .c ({y1_s3[6], y1_s2[6], y1_s1[6], y1_s0[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U738 ( .a ({temp_s3[70], temp_s2[70], temp_s1[70], temp_s0[70]}), .b ({temp_next_s3[70], temp_next_s2[70], temp_next_s1[70], temp_next_s0[70]}), .c ({y1_s3[70], y1_s2[70], y1_s1[70], y1_s0[70]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U739 ( .a ({temp_s3[71], temp_s2[71], temp_s1[71], temp_s0[71]}), .b ({temp_next_s3[71], temp_next_s2[71], temp_next_s1[71], temp_next_s0[71]}), .c ({y1_s3[71], y1_s2[71], y1_s1[71], y1_s0[71]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U740 ( .a ({temp_s3[72], temp_s2[72], temp_s1[72], temp_s0[72]}), .b ({temp_next_s3[72], temp_next_s2[72], temp_next_s1[72], temp_next_s0[72]}), .c ({y1_s3[72], y1_s2[72], y1_s1[72], y1_s0[72]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U741 ( .a ({temp_s3[73], temp_s2[73], temp_s1[73], temp_s0[73]}), .b ({temp_next_s3[73], temp_next_s2[73], temp_next_s1[73], temp_next_s0[73]}), .c ({y1_s3[73], y1_s2[73], y1_s1[73], y1_s0[73]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U742 ( .a ({temp_s3[74], temp_s2[74], temp_s1[74], temp_s0[74]}), .b ({temp_next_s3[74], temp_next_s2[74], temp_next_s1[74], temp_next_s0[74]}), .c ({y1_s3[74], y1_s2[74], y1_s1[74], y1_s0[74]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U743 ( .a ({temp_s3[75], temp_s2[75], temp_s1[75], temp_s0[75]}), .b ({temp_next_s3[75], temp_next_s2[75], temp_next_s1[75], temp_next_s0[75]}), .c ({y1_s3[75], y1_s2[75], y1_s1[75], y1_s0[75]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U744 ( .a ({temp_s3[76], temp_s2[76], temp_s1[76], temp_s0[76]}), .b ({temp_next_s3[76], temp_next_s2[76], temp_next_s1[76], temp_next_s0[76]}), .c ({y1_s3[76], y1_s2[76], y1_s1[76], y1_s0[76]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U745 ( .a ({temp_s3[77], temp_s2[77], temp_s1[77], temp_s0[77]}), .b ({temp_next_s3[77], temp_next_s2[77], temp_next_s1[77], temp_next_s0[77]}), .c ({y1_s3[77], y1_s2[77], y1_s1[77], y1_s0[77]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U746 ( .a ({temp_s3[78], temp_s2[78], temp_s1[78], temp_s0[78]}), .b ({temp_next_s3[78], temp_next_s2[78], temp_next_s1[78], temp_next_s0[78]}), .c ({y1_s3[78], y1_s2[78], y1_s1[78], y1_s0[78]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U747 ( .a ({temp_s3[79], temp_s2[79], temp_s1[79], temp_s0[79]}), .b ({temp_next_s3[79], temp_next_s2[79], temp_next_s1[79], temp_next_s0[79]}), .c ({y1_s3[79], y1_s2[79], y1_s1[79], y1_s0[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U748 ( .a ({temp_s3[7], temp_s2[7], temp_s1[7], temp_s0[7]}), .b ({temp_next_s3[7], temp_next_s2[7], temp_next_s1[7], temp_next_s0[7]}), .c ({y1_s3[7], y1_s2[7], y1_s1[7], y1_s0[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U749 ( .a ({temp_s3[80], temp_s2[80], temp_s1[80], temp_s0[80]}), .b ({temp_next_s3[80], temp_next_s2[80], temp_next_s1[80], temp_next_s0[80]}), .c ({y1_s3[80], y1_s2[80], y1_s1[80], y1_s0[80]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U750 ( .a ({temp_s3[81], temp_s2[81], temp_s1[81], temp_s0[81]}), .b ({temp_next_s3[81], temp_next_s2[81], temp_next_s1[81], temp_next_s0[81]}), .c ({y1_s3[81], y1_s2[81], y1_s1[81], y1_s0[81]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U751 ( .a ({temp_s3[82], temp_s2[82], temp_s1[82], temp_s0[82]}), .b ({temp_next_s3[82], temp_next_s2[82], temp_next_s1[82], temp_next_s0[82]}), .c ({y1_s3[82], y1_s2[82], y1_s1[82], y1_s0[82]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U752 ( .a ({temp_s3[83], temp_s2[83], temp_s1[83], temp_s0[83]}), .b ({temp_next_s3[83], temp_next_s2[83], temp_next_s1[83], temp_next_s0[83]}), .c ({y1_s3[83], y1_s2[83], y1_s1[83], y1_s0[83]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U753 ( .a ({temp_s3[84], temp_s2[84], temp_s1[84], temp_s0[84]}), .b ({temp_next_s3[84], temp_next_s2[84], temp_next_s1[84], temp_next_s0[84]}), .c ({y1_s3[84], y1_s2[84], y1_s1[84], y1_s0[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U754 ( .a ({temp_s3[85], temp_s2[85], temp_s1[85], temp_s0[85]}), .b ({temp_next_s3[85], temp_next_s2[85], temp_next_s1[85], temp_next_s0[85]}), .c ({y1_s3[85], y1_s2[85], y1_s1[85], y1_s0[85]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U755 ( .a ({temp_s3[86], temp_s2[86], temp_s1[86], temp_s0[86]}), .b ({temp_next_s3[86], temp_next_s2[86], temp_next_s1[86], temp_next_s0[86]}), .c ({y1_s3[86], y1_s2[86], y1_s1[86], y1_s0[86]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U756 ( .a ({temp_s3[87], temp_s2[87], temp_s1[87], temp_s0[87]}), .b ({temp_next_s3[87], temp_next_s2[87], temp_next_s1[87], temp_next_s0[87]}), .c ({y1_s3[87], y1_s2[87], y1_s1[87], y1_s0[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U757 ( .a ({temp_s3[88], temp_s2[88], temp_s1[88], temp_s0[88]}), .b ({temp_next_s3[88], temp_next_s2[88], temp_next_s1[88], temp_next_s0[88]}), .c ({y1_s3[88], y1_s2[88], y1_s1[88], y1_s0[88]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U758 ( .a ({temp_s3[89], temp_s2[89], temp_s1[89], temp_s0[89]}), .b ({temp_next_s3[89], temp_next_s2[89], temp_next_s1[89], temp_next_s0[89]}), .c ({y1_s3[89], y1_s2[89], y1_s1[89], y1_s0[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U759 ( .a ({temp_s3[8], temp_s2[8], temp_s1[8], temp_s0[8]}), .b ({temp_next_s3[8], temp_next_s2[8], temp_next_s1[8], temp_next_s0[8]}), .c ({y1_s3[8], y1_s2[8], y1_s1[8], y1_s0[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U760 ( .a ({temp_s3[90], temp_s2[90], temp_s1[90], temp_s0[90]}), .b ({temp_next_s3[90], temp_next_s2[90], temp_next_s1[90], temp_next_s0[90]}), .c ({y1_s3[90], y1_s2[90], y1_s1[90], y1_s0[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U761 ( .a ({temp_s3[91], temp_s2[91], temp_s1[91], temp_s0[91]}), .b ({temp_next_s3[91], temp_next_s2[91], temp_next_s1[91], temp_next_s0[91]}), .c ({y1_s3[91], y1_s2[91], y1_s1[91], y1_s0[91]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U762 ( .a ({temp_s3[92], temp_s2[92], temp_s1[92], temp_s0[92]}), .b ({temp_next_s3[92], temp_next_s2[92], temp_next_s1[92], temp_next_s0[92]}), .c ({y1_s3[92], y1_s2[92], y1_s1[92], y1_s0[92]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U763 ( .a ({temp_s3[93], temp_s2[93], temp_s1[93], temp_s0[93]}), .b ({temp_next_s3[93], temp_next_s2[93], temp_next_s1[93], temp_next_s0[93]}), .c ({y1_s3[93], y1_s2[93], y1_s1[93], y1_s0[93]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U764 ( .a ({temp_s3[94], temp_s2[94], temp_s1[94], temp_s0[94]}), .b ({temp_next_s3[94], temp_next_s2[94], temp_next_s1[94], temp_next_s0[94]}), .c ({y1_s3[94], y1_s2[94], y1_s1[94], y1_s0[94]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U765 ( .a ({temp_s3[95], temp_s2[95], temp_s1[95], temp_s0[95]}), .b ({temp_next_s3[95], temp_next_s2[95], temp_next_s1[95], temp_next_s0[95]}), .c ({y1_s3[95], y1_s2[95], y1_s1[95], y1_s0[95]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U766 ( .a ({temp_s3[96], temp_s2[96], temp_s1[96], temp_s0[96]}), .b ({temp_next_s3[96], temp_next_s2[96], temp_next_s1[96], temp_next_s0[96]}), .c ({y1_s3[96], y1_s2[96], y1_s1[96], y1_s0[96]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U767 ( .a ({temp_s3[97], temp_s2[97], temp_s1[97], temp_s0[97]}), .b ({temp_next_s3[97], temp_next_s2[97], temp_next_s1[97], temp_next_s0[97]}), .c ({y1_s3[97], y1_s2[97], y1_s1[97], y1_s0[97]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U768 ( .a ({temp_s3[98], temp_s2[98], temp_s1[98], temp_s0[98]}), .b ({temp_next_s3[98], temp_next_s2[98], temp_next_s1[98], temp_next_s0[98]}), .c ({y1_s3[98], y1_s2[98], y1_s1[98], y1_s0[98]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U769 ( .a ({temp_s3[99], temp_s2[99], temp_s1[99], temp_s0[99]}), .b ({temp_next_s3[99], temp_next_s2[99], temp_next_s1[99], temp_next_s0[99]}), .c ({y1_s3[99], y1_s2[99], y1_s1[99], y1_s0[99]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U770 ( .a ({temp_s3[9], temp_s2[9], temp_s1[9], temp_s0[9]}), .b ({temp_next_s3[9], temp_next_s2[9], temp_next_s1[9], temp_next_s0[9]}), .c ({y1_s3[9], y1_s2[9], y1_s1[9], y1_s0[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U96 ( .a ({new_AGEMA_signal_16630, new_AGEMA_signal_16629, new_AGEMA_signal_16628, mcs1_mcs_mat1_0_n128}), .b ({new_AGEMA_signal_18118, new_AGEMA_signal_18117, new_AGEMA_signal_18116, mcs1_mcs_mat1_0_n127}), .c ({temp_next_s3[93], temp_next_s2[93], temp_next_s1[93], temp_next_s0[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U95 ( .a ({new_AGEMA_signal_14407, new_AGEMA_signal_14406, new_AGEMA_signal_14405, mcs1_mcs_mat1_0_mcs_out[41]}), .b ({new_AGEMA_signal_17446, new_AGEMA_signal_17445, new_AGEMA_signal_17444, mcs1_mcs_mat1_0_mcs_out[45]}), .c ({new_AGEMA_signal_18118, new_AGEMA_signal_18117, new_AGEMA_signal_18116, mcs1_mcs_mat1_0_n127}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U94 ( .a ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, new_AGEMA_signal_10280, mcs1_mcs_mat1_0_mcs_out[33]}), .b ({new_AGEMA_signal_15790, new_AGEMA_signal_15789, new_AGEMA_signal_15788, mcs1_mcs_mat1_0_mcs_out[37]}), .c ({new_AGEMA_signal_16630, new_AGEMA_signal_16629, new_AGEMA_signal_16628, mcs1_mcs_mat1_0_n128}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U93 ( .a ({new_AGEMA_signal_17392, new_AGEMA_signal_17391, new_AGEMA_signal_17390, mcs1_mcs_mat1_0_n126}), .b ({new_AGEMA_signal_21130, new_AGEMA_signal_21129, new_AGEMA_signal_21128, mcs1_mcs_mat1_0_n125}), .c ({temp_next_s3[92], temp_next_s2[92], temp_next_s1[92], temp_next_s0[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U92 ( .a ({new_AGEMA_signal_12955, new_AGEMA_signal_12954, new_AGEMA_signal_12953, mcs1_mcs_mat1_0_mcs_out[40]}), .b ({new_AGEMA_signal_20413, new_AGEMA_signal_20412, new_AGEMA_signal_20411, mcs1_mcs_mat1_0_mcs_out[44]}), .c ({new_AGEMA_signal_21130, new_AGEMA_signal_21129, new_AGEMA_signal_21128, mcs1_mcs_mat1_0_n125}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U91 ( .a ({new_AGEMA_signal_16711, new_AGEMA_signal_16710, new_AGEMA_signal_16709, mcs1_mcs_mat1_0_mcs_out[32]}), .b ({new_AGEMA_signal_12961, new_AGEMA_signal_12960, new_AGEMA_signal_12959, mcs1_mcs_mat1_0_mcs_out[36]}), .c ({new_AGEMA_signal_17392, new_AGEMA_signal_17391, new_AGEMA_signal_17390, mcs1_mcs_mat1_0_n126}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U90 ( .a ({new_AGEMA_signal_14278, new_AGEMA_signal_14277, new_AGEMA_signal_14276, mcs1_mcs_mat1_0_n124}), .b ({new_AGEMA_signal_20362, new_AGEMA_signal_20361, new_AGEMA_signal_20360, mcs1_mcs_mat1_0_n123}), .c ({temp_next_s3[63], temp_next_s2[63], temp_next_s1[63], temp_next_s0[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U89 ( .a ({new_AGEMA_signal_12973, new_AGEMA_signal_12972, new_AGEMA_signal_12971, mcs1_mcs_mat1_0_mcs_out[27]}), .b ({new_AGEMA_signal_19528, new_AGEMA_signal_19527, new_AGEMA_signal_19526, mcs1_mcs_mat1_0_mcs_out[31]}), .c ({new_AGEMA_signal_20362, new_AGEMA_signal_20361, new_AGEMA_signal_20360, mcs1_mcs_mat1_0_n123}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U88 ( .a ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, new_AGEMA_signal_12989, mcs1_mcs_mat1_0_mcs_out[19]}), .b ({new_AGEMA_signal_12982, new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_0_mcs_out[23]}), .c ({new_AGEMA_signal_14278, new_AGEMA_signal_14277, new_AGEMA_signal_14276, mcs1_mcs_mat1_0_n124}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U87 ( .a ({new_AGEMA_signal_15718, new_AGEMA_signal_15717, new_AGEMA_signal_15716, mcs1_mcs_mat1_0_n122}), .b ({new_AGEMA_signal_19474, new_AGEMA_signal_19473, new_AGEMA_signal_19472, mcs1_mcs_mat1_0_n121}), .c ({temp_next_s3[62], temp_next_s2[62], temp_next_s1[62], temp_next_s0[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U86 ( .a ({new_AGEMA_signal_14422, new_AGEMA_signal_14421, new_AGEMA_signal_14420, mcs1_mcs_mat1_0_mcs_out[26]}), .b ({new_AGEMA_signal_18799, new_AGEMA_signal_18798, new_AGEMA_signal_18797, mcs1_mcs_mat1_0_mcs_out[30]}), .c ({new_AGEMA_signal_19474, new_AGEMA_signal_19473, new_AGEMA_signal_19472, mcs1_mcs_mat1_0_n121}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U85 ( .a ({new_AGEMA_signal_14434, new_AGEMA_signal_14433, new_AGEMA_signal_14432, mcs1_mcs_mat1_0_mcs_out[18]}), .b ({new_AGEMA_signal_14428, new_AGEMA_signal_14427, new_AGEMA_signal_14426, mcs1_mcs_mat1_0_mcs_out[22]}), .c ({new_AGEMA_signal_15718, new_AGEMA_signal_15717, new_AGEMA_signal_15716, mcs1_mcs_mat1_0_n122}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U84 ( .a ({new_AGEMA_signal_16633, new_AGEMA_signal_16632, new_AGEMA_signal_16631, mcs1_mcs_mat1_0_n120}), .b ({new_AGEMA_signal_18751, new_AGEMA_signal_18750, new_AGEMA_signal_18749, mcs1_mcs_mat1_0_n119}), .c ({temp_next_s3[61], temp_next_s2[61], temp_next_s1[61], temp_next_s0[61]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U83 ( .a ({new_AGEMA_signal_15796, new_AGEMA_signal_15795, new_AGEMA_signal_15794, mcs1_mcs_mat1_0_mcs_out[25]}), .b ({new_AGEMA_signal_18169, new_AGEMA_signal_18168, new_AGEMA_signal_18167, mcs1_mcs_mat1_0_mcs_out[29]}), .c ({new_AGEMA_signal_18751, new_AGEMA_signal_18750, new_AGEMA_signal_18749, mcs1_mcs_mat1_0_n119}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U82 ( .a ({new_AGEMA_signal_15802, new_AGEMA_signal_15801, new_AGEMA_signal_15800, mcs1_mcs_mat1_0_mcs_out[17]}), .b ({new_AGEMA_signal_15799, new_AGEMA_signal_15798, new_AGEMA_signal_15797, mcs1_mcs_mat1_0_mcs_out[21]}), .c ({new_AGEMA_signal_16633, new_AGEMA_signal_16632, new_AGEMA_signal_16631, mcs1_mcs_mat1_0_n120}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U81 ( .a ({new_AGEMA_signal_14281, new_AGEMA_signal_14280, new_AGEMA_signal_14279, mcs1_mcs_mat1_0_n118}), .b ({new_AGEMA_signal_20368, new_AGEMA_signal_20367, new_AGEMA_signal_20366, mcs1_mcs_mat1_0_n117}), .c ({temp_next_s3[60], temp_next_s2[60], temp_next_s1[60], temp_next_s0[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U80 ( .a ({new_AGEMA_signal_12979, new_AGEMA_signal_12978, new_AGEMA_signal_12977, mcs1_mcs_mat1_0_mcs_out[24]}), .b ({new_AGEMA_signal_19531, new_AGEMA_signal_19530, new_AGEMA_signal_19529, mcs1_mcs_mat1_0_mcs_out[28]}), .c ({new_AGEMA_signal_20368, new_AGEMA_signal_20367, new_AGEMA_signal_20366, mcs1_mcs_mat1_0_n117}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U79 ( .a ({new_AGEMA_signal_12997, new_AGEMA_signal_12996, new_AGEMA_signal_12995, mcs1_mcs_mat1_0_mcs_out[16]}), .b ({new_AGEMA_signal_12988, new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_0_mcs_out[20]}), .c ({new_AGEMA_signal_14281, new_AGEMA_signal_14280, new_AGEMA_signal_14279, mcs1_mcs_mat1_0_n118}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U78 ( .a ({new_AGEMA_signal_20371, new_AGEMA_signal_20370, new_AGEMA_signal_20369, mcs1_mcs_mat1_0_n116}), .b ({new_AGEMA_signal_16636, new_AGEMA_signal_16635, new_AGEMA_signal_16634, mcs1_mcs_mat1_0_n115}), .c ({temp_next_s3[31], temp_next_s2[31], temp_next_s1[31], temp_next_s0[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U77 ( .a ({new_AGEMA_signal_13012, new_AGEMA_signal_13011, new_AGEMA_signal_13010, mcs1_mcs_mat1_0_mcs_out[3]}), .b ({new_AGEMA_signal_15811, new_AGEMA_signal_15810, new_AGEMA_signal_15809, mcs1_mcs_mat1_0_mcs_out[7]}), .c ({new_AGEMA_signal_16636, new_AGEMA_signal_16635, new_AGEMA_signal_16634, mcs1_mcs_mat1_0_n115}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U76 ( .a ({new_AGEMA_signal_10570, new_AGEMA_signal_10569, new_AGEMA_signal_10568, mcs1_mcs_mat1_0_mcs_out[11]}), .b ({new_AGEMA_signal_19534, new_AGEMA_signal_19533, new_AGEMA_signal_19532, mcs1_mcs_mat1_0_mcs_out[15]}), .c ({new_AGEMA_signal_20371, new_AGEMA_signal_20370, new_AGEMA_signal_20369, mcs1_mcs_mat1_0_n116}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U75 ( .a ({new_AGEMA_signal_16642, new_AGEMA_signal_16641, new_AGEMA_signal_16640, mcs1_mcs_mat1_0_n114}), .b ({new_AGEMA_signal_16639, new_AGEMA_signal_16638, new_AGEMA_signal_16637, mcs1_mcs_mat1_0_n113}), .c ({new_AGEMA_signal_17395, new_AGEMA_signal_17394, new_AGEMA_signal_17393, mcs_out[255]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U74 ( .a ({new_AGEMA_signal_15742, new_AGEMA_signal_15741, new_AGEMA_signal_15740, mcs1_mcs_mat1_0_mcs_out[123]}), .b ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_16639, new_AGEMA_signal_16638, new_AGEMA_signal_16637, mcs1_mcs_mat1_0_n113}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U73 ( .a ({new_AGEMA_signal_14320, new_AGEMA_signal_14319, new_AGEMA_signal_14318, mcs1_mcs_mat1_0_mcs_out[115]}), .b ({new_AGEMA_signal_15748, new_AGEMA_signal_15747, new_AGEMA_signal_15746, mcs1_mcs_mat1_0_mcs_out[119]}), .c ({new_AGEMA_signal_16642, new_AGEMA_signal_16641, new_AGEMA_signal_16640, mcs1_mcs_mat1_0_n114}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U72 ( .a ({new_AGEMA_signal_16645, new_AGEMA_signal_16644, new_AGEMA_signal_16643, mcs1_mcs_mat1_0_n112}), .b ({new_AGEMA_signal_17398, new_AGEMA_signal_17397, new_AGEMA_signal_17396, mcs1_mcs_mat1_0_n111}), .c ({new_AGEMA_signal_18121, new_AGEMA_signal_18120, new_AGEMA_signal_18119, mcs_out[254]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U71 ( .a ({new_AGEMA_signal_11404, new_AGEMA_signal_11403, new_AGEMA_signal_11402, mcs1_mcs_mat1_0_mcs_out[122]}), .b ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_17398, new_AGEMA_signal_17397, new_AGEMA_signal_17396, mcs1_mcs_mat1_0_n111}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U70 ( .a ({new_AGEMA_signal_12856, new_AGEMA_signal_12855, new_AGEMA_signal_12854, mcs1_mcs_mat1_0_mcs_out[114]}), .b ({new_AGEMA_signal_15751, new_AGEMA_signal_15750, new_AGEMA_signal_15749, mcs1_mcs_mat1_0_mcs_out[118]}), .c ({new_AGEMA_signal_16645, new_AGEMA_signal_16644, new_AGEMA_signal_16643, mcs1_mcs_mat1_0_n112}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U69 ( .a ({new_AGEMA_signal_19480, new_AGEMA_signal_19479, new_AGEMA_signal_19478, mcs1_mcs_mat1_0_n110}), .b ({new_AGEMA_signal_14284, new_AGEMA_signal_14283, new_AGEMA_signal_14282, mcs1_mcs_mat1_0_n109}), .c ({temp_next_s3[30], temp_next_s2[30], temp_next_s1[30], temp_next_s0[30]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U68 ( .a ({new_AGEMA_signal_13015, new_AGEMA_signal_13014, new_AGEMA_signal_13013, mcs1_mcs_mat1_0_mcs_out[2]}), .b ({new_AGEMA_signal_13009, new_AGEMA_signal_13008, new_AGEMA_signal_13007, mcs1_mcs_mat1_0_mcs_out[6]}), .c ({new_AGEMA_signal_14284, new_AGEMA_signal_14283, new_AGEMA_signal_14282, mcs1_mcs_mat1_0_n109}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U67 ( .a ({new_AGEMA_signal_14443, new_AGEMA_signal_14442, new_AGEMA_signal_14441, mcs1_mcs_mat1_0_mcs_out[10]}), .b ({new_AGEMA_signal_18805, new_AGEMA_signal_18804, new_AGEMA_signal_18803, mcs1_mcs_mat1_0_mcs_out[14]}), .c ({new_AGEMA_signal_19480, new_AGEMA_signal_19479, new_AGEMA_signal_19478, mcs1_mcs_mat1_0_n110}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U66 ( .a ({new_AGEMA_signal_15721, new_AGEMA_signal_15720, new_AGEMA_signal_15719, mcs1_mcs_mat1_0_n108}), .b ({new_AGEMA_signal_17401, new_AGEMA_signal_17400, new_AGEMA_signal_17399, mcs1_mcs_mat1_0_n107}), .c ({new_AGEMA_signal_18124, new_AGEMA_signal_18123, new_AGEMA_signal_18122, mcs_out[253]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U65 ( .a ({new_AGEMA_signal_15745, new_AGEMA_signal_15744, new_AGEMA_signal_15743, mcs1_mcs_mat1_0_mcs_out[121]}), .b ({new_AGEMA_signal_16678, new_AGEMA_signal_16677, new_AGEMA_signal_16676, mcs1_mcs_mat1_0_mcs_out[125]}), .c ({new_AGEMA_signal_17401, new_AGEMA_signal_17400, new_AGEMA_signal_17399, mcs1_mcs_mat1_0_n107}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U64 ( .a ({new_AGEMA_signal_11419, new_AGEMA_signal_11418, new_AGEMA_signal_11417, mcs1_mcs_mat1_0_mcs_out[113]}), .b ({new_AGEMA_signal_14317, new_AGEMA_signal_14316, new_AGEMA_signal_14315, mcs1_mcs_mat1_0_mcs_out[117]}), .c ({new_AGEMA_signal_15721, new_AGEMA_signal_15720, new_AGEMA_signal_15719, mcs1_mcs_mat1_0_n108}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U63 ( .a ({new_AGEMA_signal_16651, new_AGEMA_signal_16650, new_AGEMA_signal_16649, mcs1_mcs_mat1_0_n106}), .b ({new_AGEMA_signal_16648, new_AGEMA_signal_16647, new_AGEMA_signal_16646, mcs1_mcs_mat1_0_n105}), .c ({new_AGEMA_signal_17404, new_AGEMA_signal_17403, new_AGEMA_signal_17402, mcs_out[252]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U62 ( .a ({new_AGEMA_signal_14308, new_AGEMA_signal_14307, new_AGEMA_signal_14306, mcs1_mcs_mat1_0_mcs_out[120]}), .b ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_16648, new_AGEMA_signal_16647, new_AGEMA_signal_16646, mcs1_mcs_mat1_0_n105}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U61 ( .a ({new_AGEMA_signal_15754, new_AGEMA_signal_15753, new_AGEMA_signal_15752, mcs1_mcs_mat1_0_mcs_out[112]}), .b ({new_AGEMA_signal_12853, new_AGEMA_signal_12852, new_AGEMA_signal_12851, mcs1_mcs_mat1_0_mcs_out[116]}), .c ({new_AGEMA_signal_16651, new_AGEMA_signal_16650, new_AGEMA_signal_16649, mcs1_mcs_mat1_0_n106}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U60 ( .a ({new_AGEMA_signal_15724, new_AGEMA_signal_15723, new_AGEMA_signal_15722, mcs1_mcs_mat1_0_n104}), .b ({new_AGEMA_signal_20377, new_AGEMA_signal_20376, new_AGEMA_signal_20375, mcs1_mcs_mat1_0_n103}), .c ({new_AGEMA_signal_21142, new_AGEMA_signal_21141, new_AGEMA_signal_21140, mcs_out[223]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U59 ( .a ({new_AGEMA_signal_19504, new_AGEMA_signal_19503, new_AGEMA_signal_19502, mcs1_mcs_mat1_0_mcs_out[111]}), .b ({new_AGEMA_signal_15760, new_AGEMA_signal_15759, new_AGEMA_signal_15758, mcs1_mcs_mat1_0_mcs_out[99]}), .c ({new_AGEMA_signal_20377, new_AGEMA_signal_20376, new_AGEMA_signal_20375, mcs1_mcs_mat1_0_n103}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U58 ( .a ({new_AGEMA_signal_14341, new_AGEMA_signal_14340, new_AGEMA_signal_14339, mcs1_mcs_mat1_0_mcs_out[103]}), .b ({new_AGEMA_signal_14329, new_AGEMA_signal_14328, new_AGEMA_signal_14327, mcs1_mcs_mat1_0_mcs_out[107]}), .c ({new_AGEMA_signal_15724, new_AGEMA_signal_15723, new_AGEMA_signal_15722, mcs1_mcs_mat1_0_n104}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U57 ( .a ({new_AGEMA_signal_15727, new_AGEMA_signal_15726, new_AGEMA_signal_15725, mcs1_mcs_mat1_0_n102}), .b ({new_AGEMA_signal_20380, new_AGEMA_signal_20379, new_AGEMA_signal_20378, mcs1_mcs_mat1_0_n101}), .c ({new_AGEMA_signal_21145, new_AGEMA_signal_21144, new_AGEMA_signal_21143, mcs_out[222]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U56 ( .a ({new_AGEMA_signal_19507, new_AGEMA_signal_19506, new_AGEMA_signal_19505, mcs1_mcs_mat1_0_mcs_out[110]}), .b ({new_AGEMA_signal_12883, new_AGEMA_signal_12882, new_AGEMA_signal_12881, mcs1_mcs_mat1_0_mcs_out[98]}), .c ({new_AGEMA_signal_20380, new_AGEMA_signal_20379, new_AGEMA_signal_20378, mcs1_mcs_mat1_0_n101}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U55 ( .a ({new_AGEMA_signal_11434, new_AGEMA_signal_11433, new_AGEMA_signal_11432, mcs1_mcs_mat1_0_mcs_out[102]}), .b ({new_AGEMA_signal_14332, new_AGEMA_signal_14331, new_AGEMA_signal_14330, mcs1_mcs_mat1_0_mcs_out[106]}), .c ({new_AGEMA_signal_15727, new_AGEMA_signal_15726, new_AGEMA_signal_15725, mcs1_mcs_mat1_0_n102}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U54 ( .a ({new_AGEMA_signal_15730, new_AGEMA_signal_15729, new_AGEMA_signal_15728, mcs1_mcs_mat1_0_n100}), .b ({new_AGEMA_signal_20383, new_AGEMA_signal_20382, new_AGEMA_signal_20381, mcs1_mcs_mat1_0_n99}), .c ({new_AGEMA_signal_21148, new_AGEMA_signal_21147, new_AGEMA_signal_21146, mcs_out[221]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U53 ( .a ({new_AGEMA_signal_19510, new_AGEMA_signal_19509, new_AGEMA_signal_19508, mcs1_mcs_mat1_0_mcs_out[109]}), .b ({new_AGEMA_signal_10507, new_AGEMA_signal_10506, new_AGEMA_signal_10505, mcs1_mcs_mat1_0_mcs_out[97]}), .c ({new_AGEMA_signal_20383, new_AGEMA_signal_20382, new_AGEMA_signal_20381, mcs1_mcs_mat1_0_n99}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U52 ( .a ({new_AGEMA_signal_12877, new_AGEMA_signal_12876, new_AGEMA_signal_12875, mcs1_mcs_mat1_0_mcs_out[101]}), .b ({new_AGEMA_signal_14335, new_AGEMA_signal_14334, new_AGEMA_signal_14333, mcs1_mcs_mat1_0_mcs_out[105]}), .c ({new_AGEMA_signal_15730, new_AGEMA_signal_15729, new_AGEMA_signal_15728, mcs1_mcs_mat1_0_n100}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U51 ( .a ({new_AGEMA_signal_16654, new_AGEMA_signal_16653, new_AGEMA_signal_16652, mcs1_mcs_mat1_0_n98}), .b ({new_AGEMA_signal_20386, new_AGEMA_signal_20385, new_AGEMA_signal_20384, mcs1_mcs_mat1_0_n97}), .c ({new_AGEMA_signal_21151, new_AGEMA_signal_21150, new_AGEMA_signal_21149, mcs_out[220]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U50 ( .a ({new_AGEMA_signal_19513, new_AGEMA_signal_19512, new_AGEMA_signal_19511, mcs1_mcs_mat1_0_mcs_out[108]}), .b ({new_AGEMA_signal_17422, new_AGEMA_signal_17421, new_AGEMA_signal_17420, mcs1_mcs_mat1_0_mcs_out[96]}), .c ({new_AGEMA_signal_20386, new_AGEMA_signal_20385, new_AGEMA_signal_20384, mcs1_mcs_mat1_0_n97}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U49 ( .a ({new_AGEMA_signal_14344, new_AGEMA_signal_14343, new_AGEMA_signal_14342, mcs1_mcs_mat1_0_mcs_out[100]}), .b ({new_AGEMA_signal_15757, new_AGEMA_signal_15756, new_AGEMA_signal_15755, mcs1_mcs_mat1_0_mcs_out[104]}), .c ({new_AGEMA_signal_16654, new_AGEMA_signal_16653, new_AGEMA_signal_16652, mcs1_mcs_mat1_0_n98}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U48 ( .a ({new_AGEMA_signal_14287, new_AGEMA_signal_14286, new_AGEMA_signal_14285, mcs1_mcs_mat1_0_n96}), .b ({new_AGEMA_signal_19483, new_AGEMA_signal_19482, new_AGEMA_signal_19481, mcs1_mcs_mat1_0_n95}), .c ({new_AGEMA_signal_20389, new_AGEMA_signal_20388, new_AGEMA_signal_20387, mcs_out[191]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U47 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_18775, new_AGEMA_signal_18774, new_AGEMA_signal_18773, mcs1_mcs_mat1_0_mcs_out[95]}), .c ({new_AGEMA_signal_19483, new_AGEMA_signal_19482, new_AGEMA_signal_19481, mcs1_mcs_mat1_0_n95}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U46 ( .a ({new_AGEMA_signal_12892, new_AGEMA_signal_12891, new_AGEMA_signal_12890, mcs1_mcs_mat1_0_mcs_out[83]}), .b ({new_AGEMA_signal_11449, new_AGEMA_signal_11448, new_AGEMA_signal_11447, mcs1_mcs_mat1_0_mcs_out[87]}), .c ({new_AGEMA_signal_14287, new_AGEMA_signal_14286, new_AGEMA_signal_14285, mcs1_mcs_mat1_0_n96}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U45 ( .a ({new_AGEMA_signal_14290, new_AGEMA_signal_14289, new_AGEMA_signal_14288, mcs1_mcs_mat1_0_n94}), .b ({new_AGEMA_signal_18127, new_AGEMA_signal_18126, new_AGEMA_signal_18125, mcs1_mcs_mat1_0_n93}), .c ({new_AGEMA_signal_18754, new_AGEMA_signal_18753, new_AGEMA_signal_18752, mcs_out[190]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U43 ( .a ({new_AGEMA_signal_12895, new_AGEMA_signal_12894, new_AGEMA_signal_12893, mcs1_mcs_mat1_0_mcs_out[82]}), .b ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_14290, new_AGEMA_signal_14289, new_AGEMA_signal_14288, mcs1_mcs_mat1_0_n94}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U42 ( .a ({new_AGEMA_signal_14293, new_AGEMA_signal_14292, new_AGEMA_signal_14291, mcs1_mcs_mat1_0_n92}), .b ({new_AGEMA_signal_18130, new_AGEMA_signal_18129, new_AGEMA_signal_18128, mcs1_mcs_mat1_0_n91}), .c ({new_AGEMA_signal_18757, new_AGEMA_signal_18756, new_AGEMA_signal_18755, mcs_out[189]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U41 ( .a ({new_AGEMA_signal_10516, new_AGEMA_signal_10515, new_AGEMA_signal_10514, mcs1_mcs_mat1_0_mcs_out[89]}), .b ({new_AGEMA_signal_17428, new_AGEMA_signal_17427, new_AGEMA_signal_17426, mcs1_mcs_mat1_0_mcs_out[93]}), .c ({new_AGEMA_signal_18130, new_AGEMA_signal_18129, new_AGEMA_signal_18128, mcs1_mcs_mat1_0_n91}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U40 ( .a ({new_AGEMA_signal_12898, new_AGEMA_signal_12897, new_AGEMA_signal_12896, mcs1_mcs_mat1_0_mcs_out[81]}), .b ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_14293, new_AGEMA_signal_14292, new_AGEMA_signal_14291, mcs1_mcs_mat1_0_n92}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U39 ( .a ({new_AGEMA_signal_15733, new_AGEMA_signal_15732, new_AGEMA_signal_15731, mcs1_mcs_mat1_0_n90}), .b ({new_AGEMA_signal_20392, new_AGEMA_signal_20391, new_AGEMA_signal_20390, mcs1_mcs_mat1_0_n89}), .c ({new_AGEMA_signal_21154, new_AGEMA_signal_21153, new_AGEMA_signal_21152, mcs_out[188]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U38 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_19516, new_AGEMA_signal_19515, new_AGEMA_signal_19514, mcs1_mcs_mat1_0_mcs_out[92]}), .c ({new_AGEMA_signal_20392, new_AGEMA_signal_20391, new_AGEMA_signal_20390, mcs1_mcs_mat1_0_n89}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U37 ( .a ({new_AGEMA_signal_14353, new_AGEMA_signal_14352, new_AGEMA_signal_14351, mcs1_mcs_mat1_0_mcs_out[80]}), .b ({new_AGEMA_signal_12889, new_AGEMA_signal_12888, new_AGEMA_signal_12887, mcs1_mcs_mat1_0_mcs_out[84]}), .c ({new_AGEMA_signal_15733, new_AGEMA_signal_15732, new_AGEMA_signal_15731, mcs1_mcs_mat1_0_n90}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U36 ( .a ({new_AGEMA_signal_19486, new_AGEMA_signal_19485, new_AGEMA_signal_19484, mcs1_mcs_mat1_0_n88}), .b ({new_AGEMA_signal_14296, new_AGEMA_signal_14295, new_AGEMA_signal_14294, mcs1_mcs_mat1_0_n87}), .c ({temp_next_s3[29], temp_next_s2[29], temp_next_s1[29], temp_next_s0[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U35 ( .a ({new_AGEMA_signal_10576, new_AGEMA_signal_10575, new_AGEMA_signal_10574, mcs1_mcs_mat1_0_mcs_out[5]}), .b ({new_AGEMA_signal_13003, new_AGEMA_signal_13002, new_AGEMA_signal_13001, mcs1_mcs_mat1_0_mcs_out[9]}), .c ({new_AGEMA_signal_14296, new_AGEMA_signal_14295, new_AGEMA_signal_14294, mcs1_mcs_mat1_0_n87}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U34 ( .a ({new_AGEMA_signal_18808, new_AGEMA_signal_18807, new_AGEMA_signal_18806, mcs1_mcs_mat1_0_mcs_out[13]}), .b ({new_AGEMA_signal_14452, new_AGEMA_signal_14451, new_AGEMA_signal_14450, mcs1_mcs_mat1_0_mcs_out[1]}), .c ({new_AGEMA_signal_19486, new_AGEMA_signal_19485, new_AGEMA_signal_19484, mcs1_mcs_mat1_0_n88}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U33 ( .a ({new_AGEMA_signal_16657, new_AGEMA_signal_16656, new_AGEMA_signal_16655, mcs1_mcs_mat1_0_n86}), .b ({new_AGEMA_signal_19489, new_AGEMA_signal_19488, new_AGEMA_signal_19487, mcs1_mcs_mat1_0_n85}), .c ({new_AGEMA_signal_20398, new_AGEMA_signal_20397, new_AGEMA_signal_20396, mcs_out[159]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U32 ( .a ({new_AGEMA_signal_11464, new_AGEMA_signal_11463, new_AGEMA_signal_11462, mcs1_mcs_mat1_0_mcs_out[75]}), .b ({new_AGEMA_signal_18781, new_AGEMA_signal_18780, new_AGEMA_signal_18779, mcs1_mcs_mat1_0_mcs_out[79]}), .c ({new_AGEMA_signal_19489, new_AGEMA_signal_19488, new_AGEMA_signal_19487, mcs1_mcs_mat1_0_n85}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U31 ( .a ({new_AGEMA_signal_15775, new_AGEMA_signal_15774, new_AGEMA_signal_15773, mcs1_mcs_mat1_0_mcs_out[67]}), .b ({new_AGEMA_signal_14368, new_AGEMA_signal_14367, new_AGEMA_signal_14366, mcs1_mcs_mat1_0_mcs_out[71]}), .c ({new_AGEMA_signal_16657, new_AGEMA_signal_16656, new_AGEMA_signal_16655, mcs1_mcs_mat1_0_n86}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U30 ( .a ({new_AGEMA_signal_16663, new_AGEMA_signal_16662, new_AGEMA_signal_16661, mcs1_mcs_mat1_0_n84}), .b ({new_AGEMA_signal_16660, new_AGEMA_signal_16659, new_AGEMA_signal_16658, mcs1_mcs_mat1_0_n83}), .c ({new_AGEMA_signal_17407, new_AGEMA_signal_17406, new_AGEMA_signal_17405, mcs_out[158]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U29 ( .a ({new_AGEMA_signal_15763, new_AGEMA_signal_15762, new_AGEMA_signal_15761, mcs1_mcs_mat1_0_mcs_out[74]}), .b ({new_AGEMA_signal_14356, new_AGEMA_signal_14355, new_AGEMA_signal_14354, mcs1_mcs_mat1_0_mcs_out[78]}), .c ({new_AGEMA_signal_16660, new_AGEMA_signal_16659, new_AGEMA_signal_16658, mcs1_mcs_mat1_0_n83}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U28 ( .a ({new_AGEMA_signal_14377, new_AGEMA_signal_14376, new_AGEMA_signal_14375, mcs1_mcs_mat1_0_mcs_out[66]}), .b ({new_AGEMA_signal_15769, new_AGEMA_signal_15768, new_AGEMA_signal_15767, mcs1_mcs_mat1_0_mcs_out[70]}), .c ({new_AGEMA_signal_16663, new_AGEMA_signal_16662, new_AGEMA_signal_16661, mcs1_mcs_mat1_0_n84}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U27 ( .a ({new_AGEMA_signal_16666, new_AGEMA_signal_16665, new_AGEMA_signal_16664, mcs1_mcs_mat1_0_n82}), .b ({new_AGEMA_signal_18133, new_AGEMA_signal_18132, new_AGEMA_signal_18131, mcs1_mcs_mat1_0_n81}), .c ({new_AGEMA_signal_18760, new_AGEMA_signal_18759, new_AGEMA_signal_18758, mcs_out[157]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U26 ( .a ({new_AGEMA_signal_12907, new_AGEMA_signal_12906, new_AGEMA_signal_12905, mcs1_mcs_mat1_0_mcs_out[73]}), .b ({new_AGEMA_signal_17434, new_AGEMA_signal_17433, new_AGEMA_signal_17432, mcs1_mcs_mat1_0_mcs_out[77]}), .c ({new_AGEMA_signal_18133, new_AGEMA_signal_18132, new_AGEMA_signal_18131, mcs1_mcs_mat1_0_n81}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U25 ( .a ({new_AGEMA_signal_11482, new_AGEMA_signal_11481, new_AGEMA_signal_11480, mcs1_mcs_mat1_0_mcs_out[65]}), .b ({new_AGEMA_signal_15772, new_AGEMA_signal_15771, new_AGEMA_signal_15770, mcs1_mcs_mat1_0_mcs_out[69]}), .c ({new_AGEMA_signal_16666, new_AGEMA_signal_16665, new_AGEMA_signal_16664, mcs1_mcs_mat1_0_n82}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U24 ( .a ({new_AGEMA_signal_17410, new_AGEMA_signal_17409, new_AGEMA_signal_17408, mcs1_mcs_mat1_0_n80}), .b ({new_AGEMA_signal_20401, new_AGEMA_signal_20400, new_AGEMA_signal_20399, mcs1_mcs_mat1_0_n79}), .c ({new_AGEMA_signal_21157, new_AGEMA_signal_21156, new_AGEMA_signal_21155, mcs_out[156]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U23 ( .a ({new_AGEMA_signal_15766, new_AGEMA_signal_15765, new_AGEMA_signal_15764, mcs1_mcs_mat1_0_mcs_out[72]}), .b ({new_AGEMA_signal_19519, new_AGEMA_signal_19518, new_AGEMA_signal_19517, mcs1_mcs_mat1_0_mcs_out[76]}), .c ({new_AGEMA_signal_20401, new_AGEMA_signal_20400, new_AGEMA_signal_20399, mcs1_mcs_mat1_0_n79}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U22 ( .a ({new_AGEMA_signal_16699, new_AGEMA_signal_16698, new_AGEMA_signal_16697, mcs1_mcs_mat1_0_mcs_out[64]}), .b ({new_AGEMA_signal_14374, new_AGEMA_signal_14373, new_AGEMA_signal_14372, mcs1_mcs_mat1_0_mcs_out[68]}), .c ({new_AGEMA_signal_17410, new_AGEMA_signal_17409, new_AGEMA_signal_17408, mcs1_mcs_mat1_0_n80}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U21 ( .a ({new_AGEMA_signal_15736, new_AGEMA_signal_15735, new_AGEMA_signal_15734, mcs1_mcs_mat1_0_n78}), .b ({new_AGEMA_signal_19492, new_AGEMA_signal_19491, new_AGEMA_signal_19490, mcs1_mcs_mat1_0_n77}), .c ({temp_next_s3[127], temp_next_s2[127], temp_next_s1[127], temp_next_s0[127]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U20 ( .a ({new_AGEMA_signal_12925, new_AGEMA_signal_12924, new_AGEMA_signal_12923, mcs1_mcs_mat1_0_mcs_out[59]}), .b ({new_AGEMA_signal_18787, new_AGEMA_signal_18786, new_AGEMA_signal_18785, mcs1_mcs_mat1_0_mcs_out[63]}), .c ({new_AGEMA_signal_19492, new_AGEMA_signal_19491, new_AGEMA_signal_19490, mcs1_mcs_mat1_0_n77}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U19 ( .a ({new_AGEMA_signal_11512, new_AGEMA_signal_11511, new_AGEMA_signal_11510, mcs1_mcs_mat1_0_mcs_out[51]}), .b ({new_AGEMA_signal_14389, new_AGEMA_signal_14388, new_AGEMA_signal_14387, mcs1_mcs_mat1_0_mcs_out[55]}), .c ({new_AGEMA_signal_15736, new_AGEMA_signal_15735, new_AGEMA_signal_15734, mcs1_mcs_mat1_0_n78}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U18 ( .a ({new_AGEMA_signal_16669, new_AGEMA_signal_16668, new_AGEMA_signal_16667, mcs1_mcs_mat1_0_n76}), .b ({new_AGEMA_signal_18763, new_AGEMA_signal_18762, new_AGEMA_signal_18761, mcs1_mcs_mat1_0_n75}), .c ({temp_next_s3[126], temp_next_s2[126], temp_next_s1[126], temp_next_s0[126]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U17 ( .a ({new_AGEMA_signal_11488, new_AGEMA_signal_11487, new_AGEMA_signal_11486, mcs1_mcs_mat1_0_mcs_out[58]}), .b ({new_AGEMA_signal_18154, new_AGEMA_signal_18153, new_AGEMA_signal_18152, mcs1_mcs_mat1_0_mcs_out[62]}), .c ({new_AGEMA_signal_18763, new_AGEMA_signal_18762, new_AGEMA_signal_18761, mcs1_mcs_mat1_0_n75}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U16 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_15781, new_AGEMA_signal_15780, new_AGEMA_signal_15779, mcs1_mcs_mat1_0_mcs_out[54]}), .c ({new_AGEMA_signal_16669, new_AGEMA_signal_16668, new_AGEMA_signal_16667, mcs1_mcs_mat1_0_n76}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U15 ( .a ({new_AGEMA_signal_16672, new_AGEMA_signal_16671, new_AGEMA_signal_16670, mcs1_mcs_mat1_0_n74}), .b ({new_AGEMA_signal_18766, new_AGEMA_signal_18765, new_AGEMA_signal_18764, mcs1_mcs_mat1_0_n73}), .c ({temp_next_s3[125], temp_next_s2[125], temp_next_s1[125], temp_next_s0[125]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U14 ( .a ({new_AGEMA_signal_12928, new_AGEMA_signal_12927, new_AGEMA_signal_12926, mcs1_mcs_mat1_0_mcs_out[57]}), .b ({new_AGEMA_signal_18157, new_AGEMA_signal_18156, new_AGEMA_signal_18155, mcs1_mcs_mat1_0_mcs_out[61]}), .c ({new_AGEMA_signal_18766, new_AGEMA_signal_18765, new_AGEMA_signal_18764, mcs1_mcs_mat1_0_n73}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U13 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({new_AGEMA_signal_15784, new_AGEMA_signal_15783, new_AGEMA_signal_15782, mcs1_mcs_mat1_0_mcs_out[53]}), .c ({new_AGEMA_signal_16672, new_AGEMA_signal_16671, new_AGEMA_signal_16670, mcs1_mcs_mat1_0_n74}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U12 ( .a ({new_AGEMA_signal_15739, new_AGEMA_signal_15738, new_AGEMA_signal_15737, mcs1_mcs_mat1_0_n72}), .b ({new_AGEMA_signal_20407, new_AGEMA_signal_20406, new_AGEMA_signal_20405, mcs1_mcs_mat1_0_n71}), .c ({temp_next_s3[124], temp_next_s2[124], temp_next_s1[124], temp_next_s0[124]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U11 ( .a ({new_AGEMA_signal_14386, new_AGEMA_signal_14385, new_AGEMA_signal_14384, mcs1_mcs_mat1_0_mcs_out[56]}), .b ({new_AGEMA_signal_19522, new_AGEMA_signal_19521, new_AGEMA_signal_19520, mcs1_mcs_mat1_0_mcs_out[60]}), .c ({new_AGEMA_signal_20407, new_AGEMA_signal_20406, new_AGEMA_signal_20405, mcs1_mcs_mat1_0_n71}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U10 ( .a ({new_AGEMA_signal_12940, new_AGEMA_signal_12939, new_AGEMA_signal_12938, mcs1_mcs_mat1_0_mcs_out[48]}), .b ({new_AGEMA_signal_14395, new_AGEMA_signal_14394, new_AGEMA_signal_14393, mcs1_mcs_mat1_0_mcs_out[52]}), .c ({new_AGEMA_signal_15739, new_AGEMA_signal_15738, new_AGEMA_signal_15737, mcs1_mcs_mat1_0_n72}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U9 ( .a ({new_AGEMA_signal_16675, new_AGEMA_signal_16674, new_AGEMA_signal_16673, mcs1_mcs_mat1_0_n70}), .b ({new_AGEMA_signal_19501, new_AGEMA_signal_19500, new_AGEMA_signal_19499, mcs1_mcs_mat1_0_n69}), .c ({temp_next_s3[95], temp_next_s2[95], temp_next_s1[95], temp_next_s0[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U8 ( .a ({new_AGEMA_signal_14401, new_AGEMA_signal_14400, new_AGEMA_signal_14399, mcs1_mcs_mat1_0_mcs_out[43]}), .b ({new_AGEMA_signal_18793, new_AGEMA_signal_18792, new_AGEMA_signal_18791, mcs1_mcs_mat1_0_mcs_out[47]}), .c ({new_AGEMA_signal_19501, new_AGEMA_signal_19500, new_AGEMA_signal_19499, mcs1_mcs_mat1_0_n69}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U7 ( .a ({new_AGEMA_signal_14413, new_AGEMA_signal_14412, new_AGEMA_signal_14411, mcs1_mcs_mat1_0_mcs_out[35]}), .b ({new_AGEMA_signal_15787, new_AGEMA_signal_15786, new_AGEMA_signal_15785, mcs1_mcs_mat1_0_mcs_out[39]}), .c ({new_AGEMA_signal_16675, new_AGEMA_signal_16674, new_AGEMA_signal_16673, mcs1_mcs_mat1_0_n70}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U6 ( .a ({new_AGEMA_signal_14299, new_AGEMA_signal_14298, new_AGEMA_signal_14297, mcs1_mcs_mat1_0_n68}), .b ({new_AGEMA_signal_17413, new_AGEMA_signal_17412, new_AGEMA_signal_17411, mcs1_mcs_mat1_0_n67}), .c ({temp_next_s3[94], temp_next_s2[94], temp_next_s1[94], temp_next_s0[94]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U5 ( .a ({new_AGEMA_signal_14404, new_AGEMA_signal_14403, new_AGEMA_signal_14402, mcs1_mcs_mat1_0_mcs_out[42]}), .b ({new_AGEMA_signal_16705, new_AGEMA_signal_16704, new_AGEMA_signal_16703, mcs1_mcs_mat1_0_mcs_out[46]}), .c ({new_AGEMA_signal_17413, new_AGEMA_signal_17412, new_AGEMA_signal_17411, mcs1_mcs_mat1_0_n67}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U4 ( .a ({new_AGEMA_signal_12964, new_AGEMA_signal_12963, new_AGEMA_signal_12962, mcs1_mcs_mat1_0_mcs_out[34]}), .b ({new_AGEMA_signal_11524, new_AGEMA_signal_11523, new_AGEMA_signal_11522, mcs1_mcs_mat1_0_mcs_out[38]}), .c ({new_AGEMA_signal_14299, new_AGEMA_signal_14298, new_AGEMA_signal_14297, mcs1_mcs_mat1_0_n68}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U3 ( .a ({new_AGEMA_signal_21163, new_AGEMA_signal_21162, new_AGEMA_signal_21161, mcs1_mcs_mat1_0_n66}), .b ({new_AGEMA_signal_18139, new_AGEMA_signal_18138, new_AGEMA_signal_18137, mcs1_mcs_mat1_0_n65}), .c ({temp_next_s3[28], temp_next_s2[28], temp_next_s1[28], temp_next_s0[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U2 ( .a ({new_AGEMA_signal_17467, new_AGEMA_signal_17466, new_AGEMA_signal_17465, mcs1_mcs_mat1_0_mcs_out[4]}), .b ({new_AGEMA_signal_15808, new_AGEMA_signal_15807, new_AGEMA_signal_15806, mcs1_mcs_mat1_0_mcs_out[8]}), .c ({new_AGEMA_signal_18139, new_AGEMA_signal_18138, new_AGEMA_signal_18137, mcs1_mcs_mat1_0_n65}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_U1 ( .a ({new_AGEMA_signal_14455, new_AGEMA_signal_14454, new_AGEMA_signal_14453, mcs1_mcs_mat1_0_mcs_out[0]}), .b ({new_AGEMA_signal_20416, new_AGEMA_signal_20415, new_AGEMA_signal_20414, mcs1_mcs_mat1_0_mcs_out[12]}), .c ({new_AGEMA_signal_21163, new_AGEMA_signal_21162, new_AGEMA_signal_21161, mcs1_mcs_mat1_0_n66}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_14302, new_AGEMA_signal_14301, new_AGEMA_signal_14300, mcs1_mcs_mat1_0_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_15742, new_AGEMA_signal_15741, new_AGEMA_signal_15740, mcs1_mcs_mat1_0_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_12844, new_AGEMA_signal_12843, new_AGEMA_signal_12842, mcs1_mcs_mat1_0_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_8638, new_AGEMA_signal_8637, new_AGEMA_signal_8636, mcs1_mcs_mat1_0_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_14302, new_AGEMA_signal_14301, new_AGEMA_signal_14300, mcs1_mcs_mat1_0_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_9394, new_AGEMA_signal_9393, new_AGEMA_signal_9392, mcs1_mcs_mat1_0_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_10474, new_AGEMA_signal_10473, new_AGEMA_signal_10472, mcs1_mcs_mat1_0_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_11404, new_AGEMA_signal_11403, new_AGEMA_signal_11402, mcs1_mcs_mat1_0_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_9397, new_AGEMA_signal_9396, new_AGEMA_signal_9395, mcs1_mcs_mat1_0_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .c ({new_AGEMA_signal_10474, new_AGEMA_signal_10473, new_AGEMA_signal_10472, mcs1_mcs_mat1_0_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_14305, new_AGEMA_signal_14304, new_AGEMA_signal_14303, mcs1_mcs_mat1_0_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .c ({new_AGEMA_signal_15745, new_AGEMA_signal_15744, new_AGEMA_signal_15743, mcs1_mcs_mat1_0_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_12844, new_AGEMA_signal_12843, new_AGEMA_signal_12842, mcs1_mcs_mat1_0_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_14305, new_AGEMA_signal_14304, new_AGEMA_signal_14303, mcs1_mcs_mat1_0_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_11407, new_AGEMA_signal_11406, new_AGEMA_signal_11405, mcs1_mcs_mat1_0_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_10477, new_AGEMA_signal_10476, new_AGEMA_signal_10475, mcs1_mcs_mat1_0_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_12844, new_AGEMA_signal_12843, new_AGEMA_signal_12842, mcs1_mcs_mat1_0_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_12847, new_AGEMA_signal_12846, new_AGEMA_signal_12845, mcs1_mcs_mat1_0_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_14308, new_AGEMA_signal_14307, new_AGEMA_signal_14306, mcs1_mcs_mat1_0_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_11407, new_AGEMA_signal_11406, new_AGEMA_signal_11405, mcs1_mcs_mat1_0_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9397, new_AGEMA_signal_9396, new_AGEMA_signal_9395, mcs1_mcs_mat1_0_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_12847, new_AGEMA_signal_12846, new_AGEMA_signal_12845, mcs1_mcs_mat1_0_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688]}), .c ({new_AGEMA_signal_11407, new_AGEMA_signal_11406, new_AGEMA_signal_11405, mcs1_mcs_mat1_0_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694]}), .c ({new_AGEMA_signal_9397, new_AGEMA_signal_9396, new_AGEMA_signal_9395, mcs1_mcs_mat1_0_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({new_AGEMA_signal_10477, new_AGEMA_signal_10476, new_AGEMA_signal_10475, mcs1_mcs_mat1_0_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_14311, new_AGEMA_signal_14310, new_AGEMA_signal_14309, mcs1_mcs_mat1_0_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .c ({new_AGEMA_signal_15748, new_AGEMA_signal_15747, new_AGEMA_signal_15746, mcs1_mcs_mat1_0_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_12850, new_AGEMA_signal_12849, new_AGEMA_signal_12848, mcs1_mcs_mat1_0_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10486, new_AGEMA_signal_10485, new_AGEMA_signal_10484, mcs1_mcs_mat1_0_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_14311, new_AGEMA_signal_14310, new_AGEMA_signal_14309, mcs1_mcs_mat1_0_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_14314, new_AGEMA_signal_14313, new_AGEMA_signal_14312, mcs1_mcs_mat1_0_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_11413, new_AGEMA_signal_11412, new_AGEMA_signal_11411, mcs1_mcs_mat1_0_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_15751, new_AGEMA_signal_15750, new_AGEMA_signal_15749, mcs1_mcs_mat1_0_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_12850, new_AGEMA_signal_12849, new_AGEMA_signal_12848, mcs1_mcs_mat1_0_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .c ({new_AGEMA_signal_14314, new_AGEMA_signal_14313, new_AGEMA_signal_14312, mcs1_mcs_mat1_0_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_12850, new_AGEMA_signal_12849, new_AGEMA_signal_12848, mcs1_mcs_mat1_0_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_11410, new_AGEMA_signal_11409, new_AGEMA_signal_11408, mcs1_mcs_mat1_0_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_14317, new_AGEMA_signal_14316, new_AGEMA_signal_14315, mcs1_mcs_mat1_0_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_11416, new_AGEMA_signal_11415, new_AGEMA_signal_11414, mcs1_mcs_mat1_0_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_9400, new_AGEMA_signal_9399, new_AGEMA_signal_9398, mcs1_mcs_mat1_0_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_12850, new_AGEMA_signal_12849, new_AGEMA_signal_12848, mcs1_mcs_mat1_0_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_10483, new_AGEMA_signal_10482, new_AGEMA_signal_10481, mcs1_mcs_mat1_0_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_11413, new_AGEMA_signal_11412, new_AGEMA_signal_11411, mcs1_mcs_mat1_0_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_12853, new_AGEMA_signal_12852, new_AGEMA_signal_12851, mcs1_mcs_mat1_0_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_8641, new_AGEMA_signal_8640, new_AGEMA_signal_8639, mcs1_mcs_mat1_0_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_10486, new_AGEMA_signal_10485, new_AGEMA_signal_10484, mcs1_mcs_mat1_0_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_11413, new_AGEMA_signal_11412, new_AGEMA_signal_11411, mcs1_mcs_mat1_0_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_9400, new_AGEMA_signal_9399, new_AGEMA_signal_9398, mcs1_mcs_mat1_0_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_10483, new_AGEMA_signal_10482, new_AGEMA_signal_10481, mcs1_mcs_mat1_0_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706]}), .c ({new_AGEMA_signal_11416, new_AGEMA_signal_11415, new_AGEMA_signal_11414, mcs1_mcs_mat1_0_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712]}), .c ({new_AGEMA_signal_9400, new_AGEMA_signal_9399, new_AGEMA_signal_9398, mcs1_mcs_mat1_0_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718]}), .c ({new_AGEMA_signal_10486, new_AGEMA_signal_10485, new_AGEMA_signal_10484, mcs1_mcs_mat1_0_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_12859, new_AGEMA_signal_12858, new_AGEMA_signal_12857, mcs1_mcs_mat1_0_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_9403, new_AGEMA_signal_9402, new_AGEMA_signal_9401, mcs1_mcs_mat1_0_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_14320, new_AGEMA_signal_14319, new_AGEMA_signal_14318, mcs1_mcs_mat1_0_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_10489, new_AGEMA_signal_10488, new_AGEMA_signal_10487, mcs1_mcs_mat1_0_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_10492, new_AGEMA_signal_10491, new_AGEMA_signal_10490, mcs1_mcs_mat1_0_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_11419, new_AGEMA_signal_11418, new_AGEMA_signal_11417, mcs1_mcs_mat1_0_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_12862, new_AGEMA_signal_12861, new_AGEMA_signal_12860, mcs1_mcs_mat1_0_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_14323, new_AGEMA_signal_14322, new_AGEMA_signal_14321, mcs1_mcs_mat1_0_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_15754, new_AGEMA_signal_15753, new_AGEMA_signal_15752, mcs1_mcs_mat1_0_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_12859, new_AGEMA_signal_12858, new_AGEMA_signal_12857, mcs1_mcs_mat1_0_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_14323, new_AGEMA_signal_14322, new_AGEMA_signal_14321, mcs1_mcs_mat1_0_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_8644, new_AGEMA_signal_8643, new_AGEMA_signal_8642, mcs1_mcs_mat1_0_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_11425, new_AGEMA_signal_11424, new_AGEMA_signal_11423, mcs1_mcs_mat1_0_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_12859, new_AGEMA_signal_12858, new_AGEMA_signal_12857, mcs1_mcs_mat1_0_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_9406, new_AGEMA_signal_9405, new_AGEMA_signal_9404, mcs1_mcs_mat1_0_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_11422, new_AGEMA_signal_11421, new_AGEMA_signal_11420, mcs1_mcs_mat1_0_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_12862, new_AGEMA_signal_12861, new_AGEMA_signal_12860, mcs1_mcs_mat1_0_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724]}), .c ({new_AGEMA_signal_11425, new_AGEMA_signal_11424, new_AGEMA_signal_11423, mcs1_mcs_mat1_0_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({new_AGEMA_signal_9406, new_AGEMA_signal_9405, new_AGEMA_signal_9404, mcs1_mcs_mat1_0_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736]}), .c ({new_AGEMA_signal_10492, new_AGEMA_signal_10491, new_AGEMA_signal_10490, mcs1_mcs_mat1_0_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({new_AGEMA_signal_18769, new_AGEMA_signal_18768, new_AGEMA_signal_18767, mcs1_mcs_mat1_0_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_19504, new_AGEMA_signal_19503, new_AGEMA_signal_19502, mcs1_mcs_mat1_0_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({new_AGEMA_signal_18772, new_AGEMA_signal_18771, new_AGEMA_signal_18770, mcs1_mcs_mat1_0_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_19507, new_AGEMA_signal_19506, new_AGEMA_signal_19505, mcs1_mcs_mat1_0_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_16681, new_AGEMA_signal_16680, new_AGEMA_signal_16679, mcs1_mcs_mat1_0_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_18769, new_AGEMA_signal_18768, new_AGEMA_signal_18767, mcs1_mcs_mat1_0_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_19510, new_AGEMA_signal_19509, new_AGEMA_signal_19508, mcs1_mcs_mat1_0_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_14326, new_AGEMA_signal_14325, new_AGEMA_signal_14324, mcs1_mcs_mat1_0_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_18142, new_AGEMA_signal_18141, new_AGEMA_signal_18140, mcs1_mcs_mat1_0_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_18769, new_AGEMA_signal_18768, new_AGEMA_signal_18767, mcs1_mcs_mat1_0_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_17416, new_AGEMA_signal_17415, new_AGEMA_signal_17414, mcs1_mcs_mat1_0_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_18772, new_AGEMA_signal_18771, new_AGEMA_signal_18770, mcs1_mcs_mat1_0_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_19513, new_AGEMA_signal_19512, new_AGEMA_signal_19511, mcs1_mcs_mat1_0_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_18145, new_AGEMA_signal_18144, new_AGEMA_signal_18143, mcs1_mcs_mat1_0_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_18772, new_AGEMA_signal_18771, new_AGEMA_signal_18770, mcs1_mcs_mat1_0_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_16681, new_AGEMA_signal_16680, new_AGEMA_signal_16679, mcs1_mcs_mat1_0_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_17419, new_AGEMA_signal_17418, new_AGEMA_signal_17417, mcs1_mcs_mat1_0_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_18145, new_AGEMA_signal_18144, new_AGEMA_signal_18143, mcs1_mcs_mat1_0_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742]}), .c ({new_AGEMA_signal_17419, new_AGEMA_signal_17418, new_AGEMA_signal_17417, mcs1_mcs_mat1_0_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748]}), .c ({new_AGEMA_signal_14326, new_AGEMA_signal_14325, new_AGEMA_signal_14324, mcs1_mcs_mat1_0_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754]}), .c ({new_AGEMA_signal_16681, new_AGEMA_signal_16680, new_AGEMA_signal_16679, mcs1_mcs_mat1_0_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_12871, new_AGEMA_signal_12870, new_AGEMA_signal_12869, mcs1_mcs_mat1_0_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_12868, new_AGEMA_signal_12867, new_AGEMA_signal_12866, mcs1_mcs_mat1_0_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_14329, new_AGEMA_signal_14328, new_AGEMA_signal_14327, mcs1_mcs_mat1_0_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_12868, new_AGEMA_signal_12867, new_AGEMA_signal_12866, mcs1_mcs_mat1_0_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_10495, new_AGEMA_signal_10494, new_AGEMA_signal_10493, mcs1_mcs_mat1_0_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_14332, new_AGEMA_signal_14331, new_AGEMA_signal_14330, mcs1_mcs_mat1_0_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_9409, new_AGEMA_signal_9408, new_AGEMA_signal_9407, mcs1_mcs_mat1_0_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .c ({new_AGEMA_signal_10495, new_AGEMA_signal_10494, new_AGEMA_signal_10493, mcs1_mcs_mat1_0_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({new_AGEMA_signal_12868, new_AGEMA_signal_12867, new_AGEMA_signal_12866, mcs1_mcs_mat1_0_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_14335, new_AGEMA_signal_14334, new_AGEMA_signal_14333, mcs1_mcs_mat1_0_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_11431, new_AGEMA_signal_11430, new_AGEMA_signal_11429, mcs1_mcs_mat1_0_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_8647, new_AGEMA_signal_8646, new_AGEMA_signal_8645, mcs1_mcs_mat1_0_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_12868, new_AGEMA_signal_12867, new_AGEMA_signal_12866, mcs1_mcs_mat1_0_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_14338, new_AGEMA_signal_14337, new_AGEMA_signal_14336, mcs1_mcs_mat1_0_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_15757, new_AGEMA_signal_15756, new_AGEMA_signal_15755, mcs1_mcs_mat1_0_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_12871, new_AGEMA_signal_12870, new_AGEMA_signal_12869, mcs1_mcs_mat1_0_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_11431, new_AGEMA_signal_11430, new_AGEMA_signal_11429, mcs1_mcs_mat1_0_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_14338, new_AGEMA_signal_14337, new_AGEMA_signal_14336, mcs1_mcs_mat1_0_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_11428, new_AGEMA_signal_11427, new_AGEMA_signal_11426, mcs1_mcs_mat1_0_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .c ({new_AGEMA_signal_12871, new_AGEMA_signal_12870, new_AGEMA_signal_12869, mcs1_mcs_mat1_0_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_9409, new_AGEMA_signal_9408, new_AGEMA_signal_9407, mcs1_mcs_mat1_0_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_10498, new_AGEMA_signal_10497, new_AGEMA_signal_10496, mcs1_mcs_mat1_0_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_11428, new_AGEMA_signal_11427, new_AGEMA_signal_11426, mcs1_mcs_mat1_0_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({new_AGEMA_signal_11431, new_AGEMA_signal_11430, new_AGEMA_signal_11429, mcs1_mcs_mat1_0_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766]}), .c ({new_AGEMA_signal_9409, new_AGEMA_signal_9408, new_AGEMA_signal_9407, mcs1_mcs_mat1_0_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772]}), .c ({new_AGEMA_signal_10498, new_AGEMA_signal_10497, new_AGEMA_signal_10496, mcs1_mcs_mat1_0_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_10501, new_AGEMA_signal_10500, new_AGEMA_signal_10499, mcs1_mcs_mat1_0_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_12874, new_AGEMA_signal_12873, new_AGEMA_signal_12872, mcs1_mcs_mat1_0_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_14341, new_AGEMA_signal_14340, new_AGEMA_signal_14339, mcs1_mcs_mat1_0_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_11443, new_AGEMA_signal_11442, new_AGEMA_signal_11441, mcs1_mcs_mat1_0_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_12874, new_AGEMA_signal_12873, new_AGEMA_signal_12872, mcs1_mcs_mat1_0_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_11437, new_AGEMA_signal_11436, new_AGEMA_signal_11435, mcs1_mcs_mat1_0_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_10504, new_AGEMA_signal_10503, new_AGEMA_signal_10502, mcs1_mcs_mat1_0_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_12877, new_AGEMA_signal_12876, new_AGEMA_signal_12875, mcs1_mcs_mat1_0_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_11440, new_AGEMA_signal_11439, new_AGEMA_signal_11438, mcs1_mcs_mat1_0_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_12880, new_AGEMA_signal_12879, new_AGEMA_signal_12878, mcs1_mcs_mat1_0_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_14344, new_AGEMA_signal_14343, new_AGEMA_signal_14342, mcs1_mcs_mat1_0_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_8650, new_AGEMA_signal_8649, new_AGEMA_signal_8648, mcs1_mcs_mat1_0_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_11443, new_AGEMA_signal_11442, new_AGEMA_signal_11441, mcs1_mcs_mat1_0_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_12880, new_AGEMA_signal_12879, new_AGEMA_signal_12878, mcs1_mcs_mat1_0_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_9412, new_AGEMA_signal_9411, new_AGEMA_signal_9410, mcs1_mcs_mat1_0_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .c ({new_AGEMA_signal_11440, new_AGEMA_signal_11439, new_AGEMA_signal_11438, mcs1_mcs_mat1_0_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778]}), .c ({new_AGEMA_signal_11443, new_AGEMA_signal_11442, new_AGEMA_signal_11441, mcs1_mcs_mat1_0_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784]}), .c ({new_AGEMA_signal_9412, new_AGEMA_signal_9411, new_AGEMA_signal_9410, mcs1_mcs_mat1_0_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({new_AGEMA_signal_10504, new_AGEMA_signal_10503, new_AGEMA_signal_10502, mcs1_mcs_mat1_0_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_16684, new_AGEMA_signal_16683, new_AGEMA_signal_16682, mcs1_mcs_mat1_0_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_10510, new_AGEMA_signal_10509, new_AGEMA_signal_10508, mcs1_mcs_mat1_0_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_17422, new_AGEMA_signal_17421, new_AGEMA_signal_17420, mcs1_mcs_mat1_0_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_15760, new_AGEMA_signal_15759, new_AGEMA_signal_15758, mcs1_mcs_mat1_0_mcs_out[99]}), .b ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .c ({new_AGEMA_signal_16684, new_AGEMA_signal_16683, new_AGEMA_signal_16682, mcs1_mcs_mat1_0_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_14347, new_AGEMA_signal_14346, new_AGEMA_signal_14345, mcs1_mcs_mat1_0_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .c ({new_AGEMA_signal_15760, new_AGEMA_signal_15759, new_AGEMA_signal_15758, mcs1_mcs_mat1_0_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_12883, new_AGEMA_signal_12882, new_AGEMA_signal_12881, mcs1_mcs_mat1_0_mcs_out[98]}), .b ({new_AGEMA_signal_9418, new_AGEMA_signal_9417, new_AGEMA_signal_9416, mcs1_mcs_mat1_0_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_14347, new_AGEMA_signal_14346, new_AGEMA_signal_14345, mcs1_mcs_mat1_0_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_9415, new_AGEMA_signal_9414, new_AGEMA_signal_9413, mcs1_mcs_mat1_0_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_11446, new_AGEMA_signal_11445, new_AGEMA_signal_11444, mcs1_mcs_mat1_0_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_12883, new_AGEMA_signal_12882, new_AGEMA_signal_12881, mcs1_mcs_mat1_0_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796]}), .c ({new_AGEMA_signal_11446, new_AGEMA_signal_11445, new_AGEMA_signal_11444, mcs1_mcs_mat1_0_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802]}), .c ({new_AGEMA_signal_9418, new_AGEMA_signal_9417, new_AGEMA_signal_9416, mcs1_mcs_mat1_0_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808]}), .c ({new_AGEMA_signal_10510, new_AGEMA_signal_10509, new_AGEMA_signal_10508, mcs1_mcs_mat1_0_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_18148, new_AGEMA_signal_18147, new_AGEMA_signal_18146, mcs1_mcs_mat1_0_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_18775, new_AGEMA_signal_18774, new_AGEMA_signal_18773, mcs1_mcs_mat1_0_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_16690, new_AGEMA_signal_16689, new_AGEMA_signal_16688, mcs1_mcs_mat1_0_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_16693, new_AGEMA_signal_16692, new_AGEMA_signal_16691, mcs1_mcs_mat1_0_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_17428, new_AGEMA_signal_17427, new_AGEMA_signal_17426, mcs1_mcs_mat1_0_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_18778, new_AGEMA_signal_18777, new_AGEMA_signal_18776, mcs1_mcs_mat1_0_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_14350, new_AGEMA_signal_14349, new_AGEMA_signal_14348, mcs1_mcs_mat1_0_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_19516, new_AGEMA_signal_19515, new_AGEMA_signal_19514, mcs1_mcs_mat1_0_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_18148, new_AGEMA_signal_18147, new_AGEMA_signal_18146, mcs1_mcs_mat1_0_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .c ({new_AGEMA_signal_18778, new_AGEMA_signal_18777, new_AGEMA_signal_18776, mcs1_mcs_mat1_0_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_12886, new_AGEMA_signal_12885, new_AGEMA_signal_12884, mcs1_mcs_mat1_0_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_17431, new_AGEMA_signal_17430, new_AGEMA_signal_17429, mcs1_mcs_mat1_0_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_18148, new_AGEMA_signal_18147, new_AGEMA_signal_18146, mcs1_mcs_mat1_0_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814]}), .c ({new_AGEMA_signal_17431, new_AGEMA_signal_17430, new_AGEMA_signal_17429, mcs1_mcs_mat1_0_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({new_AGEMA_signal_14350, new_AGEMA_signal_14349, new_AGEMA_signal_14348, mcs1_mcs_mat1_0_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826]}), .c ({new_AGEMA_signal_16693, new_AGEMA_signal_16692, new_AGEMA_signal_16691, mcs1_mcs_mat1_0_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_11458, new_AGEMA_signal_11457, new_AGEMA_signal_11456, mcs1_mcs_mat1_0_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_11461, new_AGEMA_signal_11460, new_AGEMA_signal_11459, mcs1_mcs_mat1_0_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_12892, new_AGEMA_signal_12891, new_AGEMA_signal_12890, mcs1_mcs_mat1_0_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_11452, new_AGEMA_signal_11451, new_AGEMA_signal_11450, mcs1_mcs_mat1_0_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_8656, new_AGEMA_signal_8655, new_AGEMA_signal_8654, mcs1_mcs_mat1_0_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_12895, new_AGEMA_signal_12894, new_AGEMA_signal_12893, mcs1_mcs_mat1_0_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_10519, new_AGEMA_signal_10518, new_AGEMA_signal_10517, mcs1_mcs_mat1_0_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_11452, new_AGEMA_signal_11451, new_AGEMA_signal_11450, mcs1_mcs_mat1_0_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_11455, new_AGEMA_signal_11454, new_AGEMA_signal_11453, mcs1_mcs_mat1_0_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_12898, new_AGEMA_signal_12897, new_AGEMA_signal_12896, mcs1_mcs_mat1_0_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_9421, new_AGEMA_signal_9420, new_AGEMA_signal_9419, mcs1_mcs_mat1_0_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_10519, new_AGEMA_signal_10518, new_AGEMA_signal_10517, mcs1_mcs_mat1_0_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_11455, new_AGEMA_signal_11454, new_AGEMA_signal_11453, mcs1_mcs_mat1_0_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_12901, new_AGEMA_signal_12900, new_AGEMA_signal_12899, mcs1_mcs_mat1_0_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .c ({new_AGEMA_signal_14353, new_AGEMA_signal_14352, new_AGEMA_signal_14351, mcs1_mcs_mat1_0_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_11458, new_AGEMA_signal_11457, new_AGEMA_signal_11456, mcs1_mcs_mat1_0_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_9421, new_AGEMA_signal_9420, new_AGEMA_signal_9419, mcs1_mcs_mat1_0_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_12901, new_AGEMA_signal_12900, new_AGEMA_signal_12899, mcs1_mcs_mat1_0_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832]}), .c ({new_AGEMA_signal_11461, new_AGEMA_signal_11460, new_AGEMA_signal_11459, mcs1_mcs_mat1_0_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838]}), .c ({new_AGEMA_signal_9421, new_AGEMA_signal_9420, new_AGEMA_signal_9419, mcs1_mcs_mat1_0_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844]}), .c ({new_AGEMA_signal_10519, new_AGEMA_signal_10518, new_AGEMA_signal_10517, mcs1_mcs_mat1_0_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_18151, new_AGEMA_signal_18150, new_AGEMA_signal_18149, mcs1_mcs_mat1_0_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_18781, new_AGEMA_signal_18780, new_AGEMA_signal_18779, mcs1_mcs_mat1_0_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_16696, new_AGEMA_signal_16695, new_AGEMA_signal_16694, mcs1_mcs_mat1_0_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_17434, new_AGEMA_signal_17433, new_AGEMA_signal_17432, mcs1_mcs_mat1_0_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_18784, new_AGEMA_signal_18783, new_AGEMA_signal_18782, mcs1_mcs_mat1_0_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_14359, new_AGEMA_signal_14358, new_AGEMA_signal_14357, mcs1_mcs_mat1_0_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_19519, new_AGEMA_signal_19518, new_AGEMA_signal_19517, mcs1_mcs_mat1_0_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_18151, new_AGEMA_signal_18150, new_AGEMA_signal_18149, mcs1_mcs_mat1_0_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .c ({new_AGEMA_signal_18784, new_AGEMA_signal_18783, new_AGEMA_signal_18782, mcs1_mcs_mat1_0_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_12904, new_AGEMA_signal_12903, new_AGEMA_signal_12902, mcs1_mcs_mat1_0_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_17437, new_AGEMA_signal_17436, new_AGEMA_signal_17435, mcs1_mcs_mat1_0_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_18151, new_AGEMA_signal_18150, new_AGEMA_signal_18149, mcs1_mcs_mat1_0_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({new_AGEMA_signal_17437, new_AGEMA_signal_17436, new_AGEMA_signal_17435, mcs1_mcs_mat1_0_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856]}), .c ({new_AGEMA_signal_14359, new_AGEMA_signal_14358, new_AGEMA_signal_14357, mcs1_mcs_mat1_0_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862]}), .c ({new_AGEMA_signal_16696, new_AGEMA_signal_16695, new_AGEMA_signal_16694, mcs1_mcs_mat1_0_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_14362, new_AGEMA_signal_14361, new_AGEMA_signal_14360, mcs1_mcs_mat1_0_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_15763, new_AGEMA_signal_15762, new_AGEMA_signal_15761, mcs1_mcs_mat1_0_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_12910, new_AGEMA_signal_12909, new_AGEMA_signal_12908, mcs1_mcs_mat1_0_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_11467, new_AGEMA_signal_11466, new_AGEMA_signal_11465, mcs1_mcs_mat1_0_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_14362, new_AGEMA_signal_14361, new_AGEMA_signal_14360, mcs1_mcs_mat1_0_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, new_AGEMA_signal_10274, mcs1_mcs_mat1_0_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_11464, new_AGEMA_signal_11463, new_AGEMA_signal_11462, mcs1_mcs_mat1_0_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_11467, new_AGEMA_signal_11466, new_AGEMA_signal_11465, mcs1_mcs_mat1_0_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, new_AGEMA_signal_10274, mcs1_mcs_mat1_0_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_12907, new_AGEMA_signal_12906, new_AGEMA_signal_12905, mcs1_mcs_mat1_0_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_9424, new_AGEMA_signal_9423, new_AGEMA_signal_9422, mcs1_mcs_mat1_0_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_9427, new_AGEMA_signal_9426, new_AGEMA_signal_9425, mcs1_mcs_mat1_0_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_10276, new_AGEMA_signal_10275, new_AGEMA_signal_10274, mcs1_mcs_mat1_0_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_10522, new_AGEMA_signal_10521, new_AGEMA_signal_10520, mcs1_mcs_mat1_0_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .c ({new_AGEMA_signal_11467, new_AGEMA_signal_11466, new_AGEMA_signal_11465, mcs1_mcs_mat1_0_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_14365, new_AGEMA_signal_14364, new_AGEMA_signal_14363, mcs1_mcs_mat1_0_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_9424, new_AGEMA_signal_9423, new_AGEMA_signal_9422, mcs1_mcs_mat1_0_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_15766, new_AGEMA_signal_15765, new_AGEMA_signal_15764, mcs1_mcs_mat1_0_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_12910, new_AGEMA_signal_12909, new_AGEMA_signal_12908, mcs1_mcs_mat1_0_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_10522, new_AGEMA_signal_10521, new_AGEMA_signal_10520, mcs1_mcs_mat1_0_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_14365, new_AGEMA_signal_14364, new_AGEMA_signal_14363, mcs1_mcs_mat1_0_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .b ({new_AGEMA_signal_11470, new_AGEMA_signal_11469, new_AGEMA_signal_11468, mcs1_mcs_mat1_0_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_12910, new_AGEMA_signal_12909, new_AGEMA_signal_12908, mcs1_mcs_mat1_0_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868]}), .c ({new_AGEMA_signal_11470, new_AGEMA_signal_11469, new_AGEMA_signal_11468, mcs1_mcs_mat1_0_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874]}), .c ({new_AGEMA_signal_9427, new_AGEMA_signal_9426, new_AGEMA_signal_9425, mcs1_mcs_mat1_0_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({new_AGEMA_signal_10522, new_AGEMA_signal_10521, new_AGEMA_signal_10520, mcs1_mcs_mat1_0_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_12913, new_AGEMA_signal_12912, new_AGEMA_signal_12911, mcs1_mcs_mat1_0_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_10525, new_AGEMA_signal_10524, new_AGEMA_signal_10523, mcs1_mcs_mat1_0_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_14368, new_AGEMA_signal_14367, new_AGEMA_signal_14366, mcs1_mcs_mat1_0_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_11476, new_AGEMA_signal_11475, new_AGEMA_signal_11474, mcs1_mcs_mat1_0_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_14371, new_AGEMA_signal_14370, new_AGEMA_signal_14369, mcs1_mcs_mat1_0_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_15769, new_AGEMA_signal_15768, new_AGEMA_signal_15767, mcs1_mcs_mat1_0_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_12913, new_AGEMA_signal_12912, new_AGEMA_signal_12911, mcs1_mcs_mat1_0_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_14371, new_AGEMA_signal_14370, new_AGEMA_signal_14369, mcs1_mcs_mat1_0_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_15772, new_AGEMA_signal_15771, new_AGEMA_signal_15770, mcs1_mcs_mat1_0_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_10525, new_AGEMA_signal_10524, new_AGEMA_signal_10523, mcs1_mcs_mat1_0_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_12916, new_AGEMA_signal_12915, new_AGEMA_signal_12914, mcs1_mcs_mat1_0_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_14371, new_AGEMA_signal_14370, new_AGEMA_signal_14369, mcs1_mcs_mat1_0_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({new_AGEMA_signal_9430, new_AGEMA_signal_9429, new_AGEMA_signal_9428, mcs1_mcs_mat1_0_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_10525, new_AGEMA_signal_10524, new_AGEMA_signal_10523, mcs1_mcs_mat1_0_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_11473, new_AGEMA_signal_11472, new_AGEMA_signal_11471, mcs1_mcs_mat1_0_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .c ({new_AGEMA_signal_12913, new_AGEMA_signal_12912, new_AGEMA_signal_12911, mcs1_mcs_mat1_0_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_10528, new_AGEMA_signal_10527, new_AGEMA_signal_10526, mcs1_mcs_mat1_0_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8662, new_AGEMA_signal_8661, new_AGEMA_signal_8660, mcs1_mcs_mat1_0_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_11473, new_AGEMA_signal_11472, new_AGEMA_signal_11471, mcs1_mcs_mat1_0_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_12916, new_AGEMA_signal_12915, new_AGEMA_signal_12914, mcs1_mcs_mat1_0_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_11476, new_AGEMA_signal_11475, new_AGEMA_signal_11474, mcs1_mcs_mat1_0_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_14374, new_AGEMA_signal_14373, new_AGEMA_signal_14372, mcs1_mcs_mat1_0_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_10528, new_AGEMA_signal_10527, new_AGEMA_signal_10526, mcs1_mcs_mat1_0_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_11476, new_AGEMA_signal_11475, new_AGEMA_signal_11474, mcs1_mcs_mat1_0_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({new_AGEMA_signal_11479, new_AGEMA_signal_11478, new_AGEMA_signal_11477, mcs1_mcs_mat1_0_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_12916, new_AGEMA_signal_12915, new_AGEMA_signal_12914, mcs1_mcs_mat1_0_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886]}), .c ({new_AGEMA_signal_11479, new_AGEMA_signal_11478, new_AGEMA_signal_11477, mcs1_mcs_mat1_0_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892]}), .c ({new_AGEMA_signal_9430, new_AGEMA_signal_9429, new_AGEMA_signal_9428, mcs1_mcs_mat1_0_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898]}), .c ({new_AGEMA_signal_10528, new_AGEMA_signal_10527, new_AGEMA_signal_10526, mcs1_mcs_mat1_0_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_14380, new_AGEMA_signal_14379, new_AGEMA_signal_14378, mcs1_mcs_mat1_0_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .c ({new_AGEMA_signal_15775, new_AGEMA_signal_15774, new_AGEMA_signal_15773, mcs1_mcs_mat1_0_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({new_AGEMA_signal_12919, new_AGEMA_signal_12918, new_AGEMA_signal_12917, mcs1_mcs_mat1_0_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_14377, new_AGEMA_signal_14376, new_AGEMA_signal_14375, mcs1_mcs_mat1_0_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_15778, new_AGEMA_signal_15777, new_AGEMA_signal_15776, mcs1_mcs_mat1_0_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_10531, new_AGEMA_signal_10530, new_AGEMA_signal_10529, mcs1_mcs_mat1_0_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_16699, new_AGEMA_signal_16698, new_AGEMA_signal_16697, mcs1_mcs_mat1_0_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_14380, new_AGEMA_signal_14379, new_AGEMA_signal_14378, mcs1_mcs_mat1_0_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .c ({new_AGEMA_signal_15778, new_AGEMA_signal_15777, new_AGEMA_signal_15776, mcs1_mcs_mat1_0_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_9433, new_AGEMA_signal_9432, new_AGEMA_signal_9431, mcs1_mcs_mat1_0_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_12919, new_AGEMA_signal_12918, new_AGEMA_signal_12917, mcs1_mcs_mat1_0_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_14380, new_AGEMA_signal_14379, new_AGEMA_signal_14378, mcs1_mcs_mat1_0_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_8665, new_AGEMA_signal_8664, new_AGEMA_signal_8663, mcs1_mcs_mat1_0_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_11485, new_AGEMA_signal_11484, new_AGEMA_signal_11483, mcs1_mcs_mat1_0_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_12919, new_AGEMA_signal_12918, new_AGEMA_signal_12917, mcs1_mcs_mat1_0_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904]}), .c ({new_AGEMA_signal_11485, new_AGEMA_signal_11484, new_AGEMA_signal_11483, mcs1_mcs_mat1_0_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({new_AGEMA_signal_9433, new_AGEMA_signal_9432, new_AGEMA_signal_9431, mcs1_mcs_mat1_0_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916]}), .c ({new_AGEMA_signal_10531, new_AGEMA_signal_10530, new_AGEMA_signal_10529, mcs1_mcs_mat1_0_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_18160, new_AGEMA_signal_18159, new_AGEMA_signal_18158, mcs1_mcs_mat1_0_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_16702, new_AGEMA_signal_16701, new_AGEMA_signal_16700, mcs1_mcs_mat1_0_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_18787, new_AGEMA_signal_18786, new_AGEMA_signal_18785, mcs1_mcs_mat1_0_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_14383, new_AGEMA_signal_14382, new_AGEMA_signal_14381, mcs1_mcs_mat1_0_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_17440, new_AGEMA_signal_17439, new_AGEMA_signal_17438, mcs1_mcs_mat1_0_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_18154, new_AGEMA_signal_18153, new_AGEMA_signal_18152, mcs1_mcs_mat1_0_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({new_AGEMA_signal_17443, new_AGEMA_signal_17442, new_AGEMA_signal_17441, mcs1_mcs_mat1_0_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_18157, new_AGEMA_signal_18156, new_AGEMA_signal_18155, mcs1_mcs_mat1_0_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922]}), .c ({new_AGEMA_signal_17443, new_AGEMA_signal_17442, new_AGEMA_signal_17441, mcs1_mcs_mat1_0_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928]}), .c ({new_AGEMA_signal_14383, new_AGEMA_signal_14382, new_AGEMA_signal_14381, mcs1_mcs_mat1_0_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934]}), .c ({new_AGEMA_signal_16702, new_AGEMA_signal_16701, new_AGEMA_signal_16700, mcs1_mcs_mat1_0_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_9439, new_AGEMA_signal_9438, new_AGEMA_signal_9437, mcs1_mcs_mat1_0_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_10534, new_AGEMA_signal_10533, new_AGEMA_signal_10532, mcs1_mcs_mat1_0_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_11488, new_AGEMA_signal_11487, new_AGEMA_signal_11486, mcs1_mcs_mat1_0_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_9442, new_AGEMA_signal_9441, new_AGEMA_signal_9440, mcs1_mcs_mat1_0_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_11491, new_AGEMA_signal_11490, new_AGEMA_signal_11489, mcs1_mcs_mat1_0_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_12928, new_AGEMA_signal_12927, new_AGEMA_signal_12926, mcs1_mcs_mat1_0_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_12931, new_AGEMA_signal_12930, new_AGEMA_signal_12929, mcs1_mcs_mat1_0_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_11494, new_AGEMA_signal_11493, new_AGEMA_signal_11492, mcs1_mcs_mat1_0_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_14386, new_AGEMA_signal_14385, new_AGEMA_signal_14384, mcs1_mcs_mat1_0_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_11497, new_AGEMA_signal_11496, new_AGEMA_signal_11495, mcs1_mcs_mat1_0_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_12931, new_AGEMA_signal_12930, new_AGEMA_signal_12929, mcs1_mcs_mat1_0_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({new_AGEMA_signal_11497, new_AGEMA_signal_11496, new_AGEMA_signal_11495, mcs1_mcs_mat1_0_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946]}), .c ({new_AGEMA_signal_9442, new_AGEMA_signal_9441, new_AGEMA_signal_9440, mcs1_mcs_mat1_0_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952]}), .c ({new_AGEMA_signal_10534, new_AGEMA_signal_10533, new_AGEMA_signal_10532, mcs1_mcs_mat1_0_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_11503, new_AGEMA_signal_11502, new_AGEMA_signal_11501, mcs1_mcs_mat1_0_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_12934, new_AGEMA_signal_12933, new_AGEMA_signal_12932, mcs1_mcs_mat1_0_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_14389, new_AGEMA_signal_14388, new_AGEMA_signal_14387, mcs1_mcs_mat1_0_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_14392, new_AGEMA_signal_14391, new_AGEMA_signal_14390, mcs1_mcs_mat1_0_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_11500, new_AGEMA_signal_11499, new_AGEMA_signal_11498, mcs1_mcs_mat1_0_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_15781, new_AGEMA_signal_15780, new_AGEMA_signal_15779, mcs1_mcs_mat1_0_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_10537, new_AGEMA_signal_10536, new_AGEMA_signal_10535, mcs1_mcs_mat1_0_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_11500, new_AGEMA_signal_11499, new_AGEMA_signal_11498, mcs1_mcs_mat1_0_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({new_AGEMA_signal_14392, new_AGEMA_signal_14391, new_AGEMA_signal_14390, mcs1_mcs_mat1_0_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_15784, new_AGEMA_signal_15783, new_AGEMA_signal_15782, mcs1_mcs_mat1_0_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_8671, new_AGEMA_signal_8670, new_AGEMA_signal_8669, mcs1_mcs_mat1_0_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_12934, new_AGEMA_signal_12933, new_AGEMA_signal_12932, mcs1_mcs_mat1_0_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_14392, new_AGEMA_signal_14391, new_AGEMA_signal_14390, mcs1_mcs_mat1_0_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_9445, new_AGEMA_signal_9444, new_AGEMA_signal_9443, mcs1_mcs_mat1_0_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_11509, new_AGEMA_signal_11508, new_AGEMA_signal_11507, mcs1_mcs_mat1_0_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_12934, new_AGEMA_signal_12933, new_AGEMA_signal_12932, mcs1_mcs_mat1_0_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_11506, new_AGEMA_signal_11505, new_AGEMA_signal_11504, mcs1_mcs_mat1_0_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_12937, new_AGEMA_signal_12936, new_AGEMA_signal_12935, mcs1_mcs_mat1_0_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_14395, new_AGEMA_signal_14394, new_AGEMA_signal_14393, mcs1_mcs_mat1_0_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_11503, new_AGEMA_signal_11502, new_AGEMA_signal_11501, mcs1_mcs_mat1_0_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_9445, new_AGEMA_signal_9444, new_AGEMA_signal_9443, mcs1_mcs_mat1_0_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_12937, new_AGEMA_signal_12936, new_AGEMA_signal_12935, mcs1_mcs_mat1_0_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_10537, new_AGEMA_signal_10536, new_AGEMA_signal_10535, mcs1_mcs_mat1_0_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_11503, new_AGEMA_signal_11502, new_AGEMA_signal_11501, mcs1_mcs_mat1_0_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958]}), .c ({new_AGEMA_signal_11509, new_AGEMA_signal_11508, new_AGEMA_signal_11507, mcs1_mcs_mat1_0_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964]}), .c ({new_AGEMA_signal_9445, new_AGEMA_signal_9444, new_AGEMA_signal_9443, mcs1_mcs_mat1_0_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({new_AGEMA_signal_10537, new_AGEMA_signal_10536, new_AGEMA_signal_10535, mcs1_mcs_mat1_0_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_16708, new_AGEMA_signal_16707, new_AGEMA_signal_16706, mcs1_mcs_mat1_0_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_17446, new_AGEMA_signal_17445, new_AGEMA_signal_17444, mcs1_mcs_mat1_0_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_19525, new_AGEMA_signal_19524, new_AGEMA_signal_19523, mcs1_mcs_mat1_0_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_14398, new_AGEMA_signal_14397, new_AGEMA_signal_14396, mcs1_mcs_mat1_0_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_20413, new_AGEMA_signal_20412, new_AGEMA_signal_20411, mcs1_mcs_mat1_0_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_18793, new_AGEMA_signal_18792, new_AGEMA_signal_18791, mcs1_mcs_mat1_0_mcs_out[47]}), .b ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .c ({new_AGEMA_signal_19525, new_AGEMA_signal_19524, new_AGEMA_signal_19523, mcs1_mcs_mat1_0_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_18163, new_AGEMA_signal_18162, new_AGEMA_signal_18161, mcs1_mcs_mat1_0_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .c ({new_AGEMA_signal_18793, new_AGEMA_signal_18792, new_AGEMA_signal_18791, mcs1_mcs_mat1_0_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_12943, new_AGEMA_signal_12942, new_AGEMA_signal_12941, mcs1_mcs_mat1_0_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_17449, new_AGEMA_signal_17448, new_AGEMA_signal_17447, mcs1_mcs_mat1_0_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_18163, new_AGEMA_signal_18162, new_AGEMA_signal_18161, mcs1_mcs_mat1_0_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976]}), .c ({new_AGEMA_signal_17449, new_AGEMA_signal_17448, new_AGEMA_signal_17447, mcs1_mcs_mat1_0_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982]}), .c ({new_AGEMA_signal_14398, new_AGEMA_signal_14397, new_AGEMA_signal_14396, mcs1_mcs_mat1_0_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988]}), .c ({new_AGEMA_signal_16708, new_AGEMA_signal_16707, new_AGEMA_signal_16706, mcs1_mcs_mat1_0_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_12946, new_AGEMA_signal_12945, new_AGEMA_signal_12944, mcs1_mcs_mat1_0_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_10540, new_AGEMA_signal_10539, new_AGEMA_signal_10538, mcs1_mcs_mat1_0_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_14401, new_AGEMA_signal_14400, new_AGEMA_signal_14399, mcs1_mcs_mat1_0_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_11515, new_AGEMA_signal_11514, new_AGEMA_signal_11513, mcs1_mcs_mat1_0_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9448, new_AGEMA_signal_9447, new_AGEMA_signal_9446, mcs1_mcs_mat1_0_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_12946, new_AGEMA_signal_12945, new_AGEMA_signal_12944, mcs1_mcs_mat1_0_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_12949, new_AGEMA_signal_12948, new_AGEMA_signal_12947, mcs1_mcs_mat1_0_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_11521, new_AGEMA_signal_11520, new_AGEMA_signal_11519, mcs1_mcs_mat1_0_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_14404, new_AGEMA_signal_14403, new_AGEMA_signal_14402, mcs1_mcs_mat1_0_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_12952, new_AGEMA_signal_12951, new_AGEMA_signal_12950, mcs1_mcs_mat1_0_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_8674, new_AGEMA_signal_8673, new_AGEMA_signal_8672, mcs1_mcs_mat1_0_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_14407, new_AGEMA_signal_14406, new_AGEMA_signal_14405, mcs1_mcs_mat1_0_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_11515, new_AGEMA_signal_11514, new_AGEMA_signal_11513, mcs1_mcs_mat1_0_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_10543, new_AGEMA_signal_10542, new_AGEMA_signal_10541, mcs1_mcs_mat1_0_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_12952, new_AGEMA_signal_12951, new_AGEMA_signal_12950, mcs1_mcs_mat1_0_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_11518, new_AGEMA_signal_11517, new_AGEMA_signal_11516, mcs1_mcs_mat1_0_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_10543, new_AGEMA_signal_10542, new_AGEMA_signal_10541, mcs1_mcs_mat1_0_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_12955, new_AGEMA_signal_12954, new_AGEMA_signal_12953, mcs1_mcs_mat1_0_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994]}), .c ({new_AGEMA_signal_11521, new_AGEMA_signal_11520, new_AGEMA_signal_11519, mcs1_mcs_mat1_0_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({new_AGEMA_signal_9448, new_AGEMA_signal_9447, new_AGEMA_signal_9446, mcs1_mcs_mat1_0_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006]}), .c ({new_AGEMA_signal_10543, new_AGEMA_signal_10542, new_AGEMA_signal_10541, mcs1_mcs_mat1_0_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_14410, new_AGEMA_signal_14409, new_AGEMA_signal_14408, mcs1_mcs_mat1_0_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_8677, new_AGEMA_signal_8676, new_AGEMA_signal_8675, mcs1_mcs_mat1_0_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_15787, new_AGEMA_signal_15786, new_AGEMA_signal_15785, mcs1_mcs_mat1_0_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_10549, new_AGEMA_signal_10548, new_AGEMA_signal_10547, mcs1_mcs_mat1_0_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_10546, new_AGEMA_signal_10545, new_AGEMA_signal_10544, mcs1_mcs_mat1_0_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_11524, new_AGEMA_signal_11523, new_AGEMA_signal_11522, mcs1_mcs_mat1_0_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({new_AGEMA_signal_14410, new_AGEMA_signal_14409, new_AGEMA_signal_14408, mcs1_mcs_mat1_0_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_15790, new_AGEMA_signal_15789, new_AGEMA_signal_15788, mcs1_mcs_mat1_0_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_11527, new_AGEMA_signal_11526, new_AGEMA_signal_11525, mcs1_mcs_mat1_0_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_12958, new_AGEMA_signal_12957, new_AGEMA_signal_12956, mcs1_mcs_mat1_0_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_14410, new_AGEMA_signal_14409, new_AGEMA_signal_14408, mcs1_mcs_mat1_0_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_11530, new_AGEMA_signal_11529, new_AGEMA_signal_11528, mcs1_mcs_mat1_0_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_10552, new_AGEMA_signal_10551, new_AGEMA_signal_10550, mcs1_mcs_mat1_0_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_12958, new_AGEMA_signal_12957, new_AGEMA_signal_12956, mcs1_mcs_mat1_0_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_11530, new_AGEMA_signal_11529, new_AGEMA_signal_11528, mcs1_mcs_mat1_0_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_10549, new_AGEMA_signal_10548, new_AGEMA_signal_10547, mcs1_mcs_mat1_0_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_12961, new_AGEMA_signal_12960, new_AGEMA_signal_12959, mcs1_mcs_mat1_0_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .b ({new_AGEMA_signal_10279, new_AGEMA_signal_10278, new_AGEMA_signal_10277, mcs1_mcs_mat1_0_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_10549, new_AGEMA_signal_10548, new_AGEMA_signal_10547, mcs1_mcs_mat1_0_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({new_AGEMA_signal_9451, new_AGEMA_signal_9450, new_AGEMA_signal_9449, mcs1_mcs_mat1_0_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_10279, new_AGEMA_signal_10278, new_AGEMA_signal_10277, mcs1_mcs_mat1_0_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012]}), .c ({new_AGEMA_signal_11530, new_AGEMA_signal_11529, new_AGEMA_signal_11528, mcs1_mcs_mat1_0_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018]}), .c ({new_AGEMA_signal_9451, new_AGEMA_signal_9450, new_AGEMA_signal_9449, mcs1_mcs_mat1_0_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024]}), .c ({new_AGEMA_signal_10552, new_AGEMA_signal_10551, new_AGEMA_signal_10550, mcs1_mcs_mat1_0_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_11533, new_AGEMA_signal_11532, new_AGEMA_signal_11531, mcs1_mcs_mat1_0_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_10555, new_AGEMA_signal_10554, new_AGEMA_signal_10553, mcs1_mcs_mat1_0_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_12964, new_AGEMA_signal_12963, new_AGEMA_signal_12962, mcs1_mcs_mat1_0_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_9454, new_AGEMA_signal_9453, new_AGEMA_signal_9452, mcs1_mcs_mat1_0_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_10282, new_AGEMA_signal_10281, new_AGEMA_signal_10280, mcs1_mcs_mat1_0_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_15793, new_AGEMA_signal_15792, new_AGEMA_signal_15791, mcs1_mcs_mat1_0_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_11536, new_AGEMA_signal_11535, new_AGEMA_signal_11534, mcs1_mcs_mat1_0_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_16711, new_AGEMA_signal_16710, new_AGEMA_signal_16709, mcs1_mcs_mat1_0_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({new_AGEMA_signal_11536, new_AGEMA_signal_11535, new_AGEMA_signal_11534, mcs1_mcs_mat1_0_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036]}), .c ({new_AGEMA_signal_9454, new_AGEMA_signal_9453, new_AGEMA_signal_9452, mcs1_mcs_mat1_0_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042]}), .c ({new_AGEMA_signal_10555, new_AGEMA_signal_10554, new_AGEMA_signal_10553, mcs1_mcs_mat1_0_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_18796, new_AGEMA_signal_18795, new_AGEMA_signal_18794, mcs1_mcs_mat1_0_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_18166, new_AGEMA_signal_18165, new_AGEMA_signal_18164, mcs1_mcs_mat1_0_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_19528, new_AGEMA_signal_19527, new_AGEMA_signal_19526, mcs1_mcs_mat1_0_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_14419, new_AGEMA_signal_14418, new_AGEMA_signal_14417, mcs1_mcs_mat1_0_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_18169, new_AGEMA_signal_18168, new_AGEMA_signal_18167, mcs1_mcs_mat1_0_mcs_out[29]}), .c ({new_AGEMA_signal_18796, new_AGEMA_signal_18795, new_AGEMA_signal_18794, mcs1_mcs_mat1_0_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_14416, new_AGEMA_signal_14415, new_AGEMA_signal_14414, mcs1_mcs_mat1_0_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_18166, new_AGEMA_signal_18165, new_AGEMA_signal_18164, mcs1_mcs_mat1_0_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_18799, new_AGEMA_signal_18798, new_AGEMA_signal_18797, mcs1_mcs_mat1_0_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_17458, new_AGEMA_signal_17457, new_AGEMA_signal_17456, mcs1_mcs_mat1_0_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .c ({new_AGEMA_signal_18166, new_AGEMA_signal_18165, new_AGEMA_signal_18164, mcs1_mcs_mat1_0_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_18802, new_AGEMA_signal_18801, new_AGEMA_signal_18800, mcs1_mcs_mat1_0_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_17452, new_AGEMA_signal_17451, new_AGEMA_signal_17450, mcs1_mcs_mat1_0_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_19531, new_AGEMA_signal_19530, new_AGEMA_signal_19529, mcs1_mcs_mat1_0_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_18172, new_AGEMA_signal_18171, new_AGEMA_signal_18170, mcs1_mcs_mat1_0_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_17455, new_AGEMA_signal_17454, new_AGEMA_signal_17453, mcs1_mcs_mat1_0_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_18802, new_AGEMA_signal_18801, new_AGEMA_signal_18800, mcs1_mcs_mat1_0_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_16714, new_AGEMA_signal_16713, new_AGEMA_signal_16712, mcs1_mcs_mat1_0_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_17455, new_AGEMA_signal_17454, new_AGEMA_signal_17453, mcs1_mcs_mat1_0_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_17458, new_AGEMA_signal_17457, new_AGEMA_signal_17456, mcs1_mcs_mat1_0_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_14419, new_AGEMA_signal_14418, new_AGEMA_signal_14417, mcs1_mcs_mat1_0_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_18172, new_AGEMA_signal_18171, new_AGEMA_signal_18170, mcs1_mcs_mat1_0_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048]}), .c ({new_AGEMA_signal_17458, new_AGEMA_signal_17457, new_AGEMA_signal_17456, mcs1_mcs_mat1_0_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054]}), .c ({new_AGEMA_signal_14419, new_AGEMA_signal_14418, new_AGEMA_signal_14417, mcs1_mcs_mat1_0_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({new_AGEMA_signal_16714, new_AGEMA_signal_16713, new_AGEMA_signal_16712, mcs1_mcs_mat1_0_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_11539, new_AGEMA_signal_11538, new_AGEMA_signal_11537, mcs1_mcs_mat1_0_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_12973, new_AGEMA_signal_12972, new_AGEMA_signal_12971, mcs1_mcs_mat1_0_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_10558, new_AGEMA_signal_10557, new_AGEMA_signal_10556, mcs1_mcs_mat1_0_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_9457, new_AGEMA_signal_9456, new_AGEMA_signal_9455, mcs1_mcs_mat1_0_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_11539, new_AGEMA_signal_11538, new_AGEMA_signal_11537, mcs1_mcs_mat1_0_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_12976, new_AGEMA_signal_12975, new_AGEMA_signal_12974, mcs1_mcs_mat1_0_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_14422, new_AGEMA_signal_14421, new_AGEMA_signal_14420, mcs1_mcs_mat1_0_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_11545, new_AGEMA_signal_11544, new_AGEMA_signal_11543, mcs1_mcs_mat1_0_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_9457, new_AGEMA_signal_9456, new_AGEMA_signal_9455, mcs1_mcs_mat1_0_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_12976, new_AGEMA_signal_12975, new_AGEMA_signal_12974, mcs1_mcs_mat1_0_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_14425, new_AGEMA_signal_14424, new_AGEMA_signal_14423, mcs1_mcs_mat1_0_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .c ({new_AGEMA_signal_15796, new_AGEMA_signal_15795, new_AGEMA_signal_15794, mcs1_mcs_mat1_0_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_11545, new_AGEMA_signal_11544, new_AGEMA_signal_11543, mcs1_mcs_mat1_0_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_12979, new_AGEMA_signal_12978, new_AGEMA_signal_12977, mcs1_mcs_mat1_0_mcs_out[24]}), .c ({new_AGEMA_signal_14425, new_AGEMA_signal_14424, new_AGEMA_signal_14423, mcs1_mcs_mat1_0_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_11542, new_AGEMA_signal_11541, new_AGEMA_signal_11540, mcs1_mcs_mat1_0_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .c ({new_AGEMA_signal_12979, new_AGEMA_signal_12978, new_AGEMA_signal_12977, mcs1_mcs_mat1_0_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_10558, new_AGEMA_signal_10557, new_AGEMA_signal_10556, mcs1_mcs_mat1_0_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8683, new_AGEMA_signal_8682, new_AGEMA_signal_8681, mcs1_mcs_mat1_0_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_11542, new_AGEMA_signal_11541, new_AGEMA_signal_11540, mcs1_mcs_mat1_0_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066]}), .c ({new_AGEMA_signal_11545, new_AGEMA_signal_11544, new_AGEMA_signal_11543, mcs1_mcs_mat1_0_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072]}), .c ({new_AGEMA_signal_9457, new_AGEMA_signal_9456, new_AGEMA_signal_9455, mcs1_mcs_mat1_0_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078]}), .c ({new_AGEMA_signal_10558, new_AGEMA_signal_10557, new_AGEMA_signal_10556, mcs1_mcs_mat1_0_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_11548, new_AGEMA_signal_11547, new_AGEMA_signal_11546, mcs1_mcs_mat1_0_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .c ({new_AGEMA_signal_12982, new_AGEMA_signal_12981, new_AGEMA_signal_12980, mcs1_mcs_mat1_0_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_10561, new_AGEMA_signal_10560, new_AGEMA_signal_10559, mcs1_mcs_mat1_0_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_9460, new_AGEMA_signal_9459, new_AGEMA_signal_9458, mcs1_mcs_mat1_0_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_11548, new_AGEMA_signal_11547, new_AGEMA_signal_11546, mcs1_mcs_mat1_0_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, new_AGEMA_signal_12983, mcs1_mcs_mat1_0_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .c ({new_AGEMA_signal_14428, new_AGEMA_signal_14427, new_AGEMA_signal_14426, mcs1_mcs_mat1_0_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_11554, new_AGEMA_signal_11553, new_AGEMA_signal_11552, mcs1_mcs_mat1_0_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_9460, new_AGEMA_signal_9459, new_AGEMA_signal_9458, mcs1_mcs_mat1_0_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_12985, new_AGEMA_signal_12984, new_AGEMA_signal_12983, mcs1_mcs_mat1_0_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_14431, new_AGEMA_signal_14430, new_AGEMA_signal_14429, mcs1_mcs_mat1_0_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_8413, new_AGEMA_signal_8412, new_AGEMA_signal_8411, mcs1_mcs_mat1_0_mcs_out[86]}), .c ({new_AGEMA_signal_15799, new_AGEMA_signal_15798, new_AGEMA_signal_15797, mcs1_mcs_mat1_0_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_11554, new_AGEMA_signal_11553, new_AGEMA_signal_11552, mcs1_mcs_mat1_0_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_12988, new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_0_mcs_out[20]}), .c ({new_AGEMA_signal_14431, new_AGEMA_signal_14430, new_AGEMA_signal_14429, mcs1_mcs_mat1_0_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_11551, new_AGEMA_signal_11550, new_AGEMA_signal_11549, mcs1_mcs_mat1_0_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .c ({new_AGEMA_signal_12988, new_AGEMA_signal_12987, new_AGEMA_signal_12986, mcs1_mcs_mat1_0_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_10561, new_AGEMA_signal_10560, new_AGEMA_signal_10559, mcs1_mcs_mat1_0_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8686, new_AGEMA_signal_8685, new_AGEMA_signal_8684, mcs1_mcs_mat1_0_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_11551, new_AGEMA_signal_11550, new_AGEMA_signal_11549, mcs1_mcs_mat1_0_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084]}), .c ({new_AGEMA_signal_11554, new_AGEMA_signal_11553, new_AGEMA_signal_11552, mcs1_mcs_mat1_0_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({new_AGEMA_signal_9460, new_AGEMA_signal_9459, new_AGEMA_signal_9458, mcs1_mcs_mat1_0_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096]}), .c ({new_AGEMA_signal_10561, new_AGEMA_signal_10560, new_AGEMA_signal_10559, mcs1_mcs_mat1_0_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_11557, new_AGEMA_signal_11556, new_AGEMA_signal_11555, mcs1_mcs_mat1_0_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_11566, new_AGEMA_signal_11565, new_AGEMA_signal_11564, mcs1_mcs_mat1_0_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_12991, new_AGEMA_signal_12990, new_AGEMA_signal_12989, mcs1_mcs_mat1_0_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_12994, new_AGEMA_signal_12993, new_AGEMA_signal_12992, mcs1_mcs_mat1_0_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_8689, new_AGEMA_signal_8688, new_AGEMA_signal_8687, mcs1_mcs_mat1_0_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_14434, new_AGEMA_signal_14433, new_AGEMA_signal_14432, mcs1_mcs_mat1_0_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_14437, new_AGEMA_signal_14436, new_AGEMA_signal_14435, mcs1_mcs_mat1_0_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_9463, new_AGEMA_signal_9462, new_AGEMA_signal_9461, mcs1_mcs_mat1_0_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_15802, new_AGEMA_signal_15801, new_AGEMA_signal_15800, mcs1_mcs_mat1_0_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_8431, new_AGEMA_signal_8430, new_AGEMA_signal_8429, mcs1_mcs_mat1_0_mcs_out[50]}), .b ({new_AGEMA_signal_12994, new_AGEMA_signal_12993, new_AGEMA_signal_12992, mcs1_mcs_mat1_0_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_14437, new_AGEMA_signal_14436, new_AGEMA_signal_14435, mcs1_mcs_mat1_0_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_11560, new_AGEMA_signal_11559, new_AGEMA_signal_11558, mcs1_mcs_mat1_0_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .c ({new_AGEMA_signal_12994, new_AGEMA_signal_12993, new_AGEMA_signal_12992, mcs1_mcs_mat1_0_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_10564, new_AGEMA_signal_10563, new_AGEMA_signal_10562, mcs1_mcs_mat1_0_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_10567, new_AGEMA_signal_10566, new_AGEMA_signal_10565, mcs1_mcs_mat1_0_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_11560, new_AGEMA_signal_11559, new_AGEMA_signal_11558, mcs1_mcs_mat1_0_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_11563, new_AGEMA_signal_11562, new_AGEMA_signal_11561, mcs1_mcs_mat1_0_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_9463, new_AGEMA_signal_9462, new_AGEMA_signal_9461, mcs1_mcs_mat1_0_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_12997, new_AGEMA_signal_12996, new_AGEMA_signal_12995, mcs1_mcs_mat1_0_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102]}), .c ({new_AGEMA_signal_11566, new_AGEMA_signal_11565, new_AGEMA_signal_11564, mcs1_mcs_mat1_0_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108]}), .c ({new_AGEMA_signal_9463, new_AGEMA_signal_9462, new_AGEMA_signal_9461, mcs1_mcs_mat1_0_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114]}), .c ({new_AGEMA_signal_10567, new_AGEMA_signal_10566, new_AGEMA_signal_10565, mcs1_mcs_mat1_0_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_18811, new_AGEMA_signal_18810, new_AGEMA_signal_18809, mcs1_mcs_mat1_0_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_15805, new_AGEMA_signal_15804, new_AGEMA_signal_15803, mcs1_mcs_mat1_0_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_19534, new_AGEMA_signal_19533, new_AGEMA_signal_19532, mcs1_mcs_mat1_0_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_18181, new_AGEMA_signal_18180, new_AGEMA_signal_18179, mcs1_mcs_mat1_0_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_18175, new_AGEMA_signal_18174, new_AGEMA_signal_18173, mcs1_mcs_mat1_0_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_18805, new_AGEMA_signal_18804, new_AGEMA_signal_18803, mcs1_mcs_mat1_0_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_17464, new_AGEMA_signal_17463, new_AGEMA_signal_17462, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_14440, new_AGEMA_signal_14439, new_AGEMA_signal_14438, mcs1_mcs_mat1_0_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_18175, new_AGEMA_signal_18174, new_AGEMA_signal_18173, mcs1_mcs_mat1_0_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_15805, new_AGEMA_signal_15804, new_AGEMA_signal_15803, mcs1_mcs_mat1_0_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_18178, new_AGEMA_signal_18177, new_AGEMA_signal_18176, mcs1_mcs_mat1_0_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_18808, new_AGEMA_signal_18807, new_AGEMA_signal_18806, mcs1_mcs_mat1_0_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_17461, new_AGEMA_signal_17460, new_AGEMA_signal_17459, mcs1_mcs_mat1_0_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_17464, new_AGEMA_signal_17463, new_AGEMA_signal_17462, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_18178, new_AGEMA_signal_18177, new_AGEMA_signal_18176, mcs1_mcs_mat1_0_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_13000, new_AGEMA_signal_12999, new_AGEMA_signal_12998, mcs1_mcs_mat1_0_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_14440, new_AGEMA_signal_14439, new_AGEMA_signal_14438, mcs1_mcs_mat1_0_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_15805, new_AGEMA_signal_15804, new_AGEMA_signal_15803, mcs1_mcs_mat1_0_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_19537, new_AGEMA_signal_19536, new_AGEMA_signal_19535, mcs1_mcs_mat1_0_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .c ({new_AGEMA_signal_20416, new_AGEMA_signal_20415, new_AGEMA_signal_20414, mcs1_mcs_mat1_0_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_18811, new_AGEMA_signal_18810, new_AGEMA_signal_18809, mcs1_mcs_mat1_0_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_17464, new_AGEMA_signal_17463, new_AGEMA_signal_17462, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_19537, new_AGEMA_signal_19536, new_AGEMA_signal_19535, mcs1_mcs_mat1_0_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({new_AGEMA_signal_18181, new_AGEMA_signal_18180, new_AGEMA_signal_18179, mcs1_mcs_mat1_0_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_18811, new_AGEMA_signal_18810, new_AGEMA_signal_18809, mcs1_mcs_mat1_0_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({new_AGEMA_signal_17461, new_AGEMA_signal_17460, new_AGEMA_signal_17459, mcs1_mcs_mat1_0_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_18181, new_AGEMA_signal_18180, new_AGEMA_signal_18179, mcs1_mcs_mat1_0_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_11383, new_AGEMA_signal_11382, new_AGEMA_signal_11381, shiftr_out[124]}), .b ({new_AGEMA_signal_16717, new_AGEMA_signal_16716, new_AGEMA_signal_16715, mcs1_mcs_mat1_0_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_17461, new_AGEMA_signal_17460, new_AGEMA_signal_17459, mcs1_mcs_mat1_0_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16609, new_AGEMA_signal_16608, new_AGEMA_signal_16607, mcs1_mcs_mat1_0_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({new_AGEMA_signal_17464, new_AGEMA_signal_17463, new_AGEMA_signal_17462, mcs1_mcs_mat1_0_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12823, new_AGEMA_signal_12822, new_AGEMA_signal_12821, mcs1_mcs_mat1_0_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126]}), .c ({new_AGEMA_signal_14440, new_AGEMA_signal_14439, new_AGEMA_signal_14438, mcs1_mcs_mat1_0_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15697, new_AGEMA_signal_15696, new_AGEMA_signal_15695, mcs1_mcs_mat1_0_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132]}), .c ({new_AGEMA_signal_16717, new_AGEMA_signal_16716, new_AGEMA_signal_16715, mcs1_mcs_mat1_0_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_10285, new_AGEMA_signal_10284, new_AGEMA_signal_10283, mcs1_mcs_mat1_0_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .c ({new_AGEMA_signal_10570, new_AGEMA_signal_10569, new_AGEMA_signal_10568, mcs1_mcs_mat1_0_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_13006, new_AGEMA_signal_13005, new_AGEMA_signal_13004, mcs1_mcs_mat1_0_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .c ({new_AGEMA_signal_14443, new_AGEMA_signal_14442, new_AGEMA_signal_14441, mcs1_mcs_mat1_0_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_11569, new_AGEMA_signal_11568, new_AGEMA_signal_11567, mcs1_mcs_mat1_0_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .c ({new_AGEMA_signal_13003, new_AGEMA_signal_13002, new_AGEMA_signal_13001, mcs1_mcs_mat1_0_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_10573, new_AGEMA_signal_10572, new_AGEMA_signal_10571, mcs1_mcs_mat1_0_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_10285, new_AGEMA_signal_10284, new_AGEMA_signal_10283, mcs1_mcs_mat1_0_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_11569, new_AGEMA_signal_11568, new_AGEMA_signal_11567, mcs1_mcs_mat1_0_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_8692, new_AGEMA_signal_8691, new_AGEMA_signal_8690, mcs1_mcs_mat1_0_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_9466, new_AGEMA_signal_9465, new_AGEMA_signal_9464, mcs1_mcs_mat1_0_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_10285, new_AGEMA_signal_10284, new_AGEMA_signal_10283, mcs1_mcs_mat1_0_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_14446, new_AGEMA_signal_14445, new_AGEMA_signal_14444, mcs1_mcs_mat1_0_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_8395, new_AGEMA_signal_8394, new_AGEMA_signal_8393, shiftr_out[92]}), .c ({new_AGEMA_signal_15808, new_AGEMA_signal_15807, new_AGEMA_signal_15806, mcs1_mcs_mat1_0_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_8692, new_AGEMA_signal_8691, new_AGEMA_signal_8690, mcs1_mcs_mat1_0_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_13006, new_AGEMA_signal_13005, new_AGEMA_signal_13004, mcs1_mcs_mat1_0_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_14446, new_AGEMA_signal_14445, new_AGEMA_signal_14444, mcs1_mcs_mat1_0_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_11572, new_AGEMA_signal_11571, new_AGEMA_signal_11570, mcs1_mcs_mat1_0_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_10573, new_AGEMA_signal_10572, new_AGEMA_signal_10571, mcs1_mcs_mat1_0_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_13006, new_AGEMA_signal_13005, new_AGEMA_signal_13004, mcs1_mcs_mat1_0_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10435, new_AGEMA_signal_10434, new_AGEMA_signal_10433, mcs1_mcs_mat1_0_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138]}), .c ({new_AGEMA_signal_11572, new_AGEMA_signal_11571, new_AGEMA_signal_11570, mcs1_mcs_mat1_0_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8599, new_AGEMA_signal_8598, new_AGEMA_signal_8597, mcs1_mcs_mat1_0_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144]}), .c ({new_AGEMA_signal_9466, new_AGEMA_signal_9465, new_AGEMA_signal_9464, mcs1_mcs_mat1_0_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10236, new_AGEMA_signal_10235, shiftr_out[95]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({new_AGEMA_signal_10573, new_AGEMA_signal_10572, new_AGEMA_signal_10571, mcs1_mcs_mat1_0_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_16720, new_AGEMA_signal_16719, new_AGEMA_signal_16718, mcs1_mcs_mat1_0_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_10579, new_AGEMA_signal_10578, new_AGEMA_signal_10577, mcs1_mcs_mat1_0_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_17467, new_AGEMA_signal_17466, new_AGEMA_signal_17465, mcs1_mcs_mat1_0_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_15811, new_AGEMA_signal_15810, new_AGEMA_signal_15809, mcs1_mcs_mat1_0_mcs_out[7]}), .b ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .c ({new_AGEMA_signal_16720, new_AGEMA_signal_16719, new_AGEMA_signal_16718, mcs1_mcs_mat1_0_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_14449, new_AGEMA_signal_14448, new_AGEMA_signal_14447, mcs1_mcs_mat1_0_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .c ({new_AGEMA_signal_15811, new_AGEMA_signal_15810, new_AGEMA_signal_15809, mcs1_mcs_mat1_0_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_13009, new_AGEMA_signal_13008, new_AGEMA_signal_13007, mcs1_mcs_mat1_0_mcs_out[6]}), .b ({new_AGEMA_signal_9472, new_AGEMA_signal_9471, new_AGEMA_signal_9470, mcs1_mcs_mat1_0_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_14449, new_AGEMA_signal_14448, new_AGEMA_signal_14447, mcs1_mcs_mat1_0_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_9469, new_AGEMA_signal_9468, new_AGEMA_signal_9467, mcs1_mcs_mat1_0_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_11575, new_AGEMA_signal_11574, new_AGEMA_signal_11573, mcs1_mcs_mat1_0_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_13009, new_AGEMA_signal_13008, new_AGEMA_signal_13007, mcs1_mcs_mat1_0_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10452, new_AGEMA_signal_10451, shiftr_out[61]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156]}), .c ({new_AGEMA_signal_11575, new_AGEMA_signal_11574, new_AGEMA_signal_11573, mcs1_mcs_mat1_0_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8616, new_AGEMA_signal_8615, shiftr_out[62]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162]}), .c ({new_AGEMA_signal_9472, new_AGEMA_signal_9471, new_AGEMA_signal_9470, mcs1_mcs_mat1_0_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10255, new_AGEMA_signal_10254, new_AGEMA_signal_10253, mcs1_mcs_mat1_0_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168]}), .c ({new_AGEMA_signal_10579, new_AGEMA_signal_10578, new_AGEMA_signal_10577, mcs1_mcs_mat1_0_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_10582, new_AGEMA_signal_10581, new_AGEMA_signal_10580, mcs1_mcs_mat1_0_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_11578, new_AGEMA_signal_11577, new_AGEMA_signal_11576, mcs1_mcs_mat1_0_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_13015, new_AGEMA_signal_13014, new_AGEMA_signal_13013, mcs1_mcs_mat1_0_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .b ({new_AGEMA_signal_10585, new_AGEMA_signal_10584, new_AGEMA_signal_10583, mcs1_mcs_mat1_0_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_11578, new_AGEMA_signal_11577, new_AGEMA_signal_11576, mcs1_mcs_mat1_0_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_13018, new_AGEMA_signal_13017, new_AGEMA_signal_13016, mcs1_mcs_mat1_0_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_9475, new_AGEMA_signal_9474, new_AGEMA_signal_9473, mcs1_mcs_mat1_0_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_14452, new_AGEMA_signal_14451, new_AGEMA_signal_14450, mcs1_mcs_mat1_0_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_13021, new_AGEMA_signal_13020, new_AGEMA_signal_13019, mcs1_mcs_mat1_0_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_11584, new_AGEMA_signal_11583, new_AGEMA_signal_11582, mcs1_mcs_mat1_0_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_14455, new_AGEMA_signal_14454, new_AGEMA_signal_14453, mcs1_mcs_mat1_0_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_11587, new_AGEMA_signal_11586, new_AGEMA_signal_11585, mcs1_mcs_mat1_0_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_8698, new_AGEMA_signal_8697, new_AGEMA_signal_8696, mcs1_mcs_mat1_0_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_13021, new_AGEMA_signal_13020, new_AGEMA_signal_13019, mcs1_mcs_mat1_0_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10471, new_AGEMA_signal_10470, new_AGEMA_signal_10469, shiftr_out[29]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174]}), .c ({new_AGEMA_signal_11587, new_AGEMA_signal_11586, new_AGEMA_signal_11585, mcs1_mcs_mat1_0_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8635, new_AGEMA_signal_8634, new_AGEMA_signal_8633, shiftr_out[30]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({new_AGEMA_signal_9475, new_AGEMA_signal_9474, new_AGEMA_signal_9473, mcs1_mcs_mat1_0_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_0_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10272, new_AGEMA_signal_10271, mcs1_mcs_mat1_0_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186]}), .c ({new_AGEMA_signal_10585, new_AGEMA_signal_10584, new_AGEMA_signal_10583, mcs1_mcs_mat1_0_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U96 ( .a ({new_AGEMA_signal_16723, new_AGEMA_signal_16722, new_AGEMA_signal_16721, mcs1_mcs_mat1_1_n128}), .b ({new_AGEMA_signal_15814, new_AGEMA_signal_15813, new_AGEMA_signal_15812, mcs1_mcs_mat1_1_n127}), .c ({temp_next_s3[89], temp_next_s2[89], temp_next_s1[89], temp_next_s0[89]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U95 ( .a ({new_AGEMA_signal_14584, new_AGEMA_signal_14583, new_AGEMA_signal_14582, mcs1_mcs_mat1_1_mcs_out[41]}), .b ({new_AGEMA_signal_11695, new_AGEMA_signal_11694, new_AGEMA_signal_11693, mcs1_mcs_mat1_1_mcs_out[45]}), .c ({new_AGEMA_signal_15814, new_AGEMA_signal_15813, new_AGEMA_signal_15812, mcs1_mcs_mat1_1_n127}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U94 ( .a ({new_AGEMA_signal_15913, new_AGEMA_signal_15912, new_AGEMA_signal_15911, mcs1_mcs_mat1_1_mcs_out[33]}), .b ({new_AGEMA_signal_15910, new_AGEMA_signal_15909, new_AGEMA_signal_15908, mcs1_mcs_mat1_1_mcs_out[37]}), .c ({new_AGEMA_signal_16723, new_AGEMA_signal_16722, new_AGEMA_signal_16721, mcs1_mcs_mat1_1_n128}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U93 ( .a ({new_AGEMA_signal_21166, new_AGEMA_signal_21165, new_AGEMA_signal_21164, mcs1_mcs_mat1_1_n126}), .b ({new_AGEMA_signal_17473, new_AGEMA_signal_17472, new_AGEMA_signal_17471, mcs1_mcs_mat1_1_n125}), .c ({temp_next_s3[88], temp_next_s2[88], temp_next_s1[88], temp_next_s0[88]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U92 ( .a ({new_AGEMA_signal_13135, new_AGEMA_signal_13134, new_AGEMA_signal_13133, mcs1_mcs_mat1_1_mcs_out[40]}), .b ({new_AGEMA_signal_16783, new_AGEMA_signal_16782, new_AGEMA_signal_16781, mcs1_mcs_mat1_1_mcs_out[44]}), .c ({new_AGEMA_signal_17473, new_AGEMA_signal_17472, new_AGEMA_signal_17471, mcs1_mcs_mat1_1_n125}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U91 ( .a ({new_AGEMA_signal_20458, new_AGEMA_signal_20457, new_AGEMA_signal_20456, mcs1_mcs_mat1_1_mcs_out[32]}), .b ({new_AGEMA_signal_13141, new_AGEMA_signal_13140, new_AGEMA_signal_13139, mcs1_mcs_mat1_1_mcs_out[36]}), .c ({new_AGEMA_signal_21166, new_AGEMA_signal_21165, new_AGEMA_signal_21164, mcs1_mcs_mat1_1_n126}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U90 ( .a ({new_AGEMA_signal_18814, new_AGEMA_signal_18813, new_AGEMA_signal_18812, mcs1_mcs_mat1_1_n124}), .b ({new_AGEMA_signal_16726, new_AGEMA_signal_16725, new_AGEMA_signal_16724, mcs1_mcs_mat1_1_n123}), .c ({temp_next_s3[59], temp_next_s2[59], temp_next_s1[59], temp_next_s0[59]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U89 ( .a ({new_AGEMA_signal_13156, new_AGEMA_signal_13155, new_AGEMA_signal_13154, mcs1_mcs_mat1_1_mcs_out[27]}), .b ({new_AGEMA_signal_15916, new_AGEMA_signal_15915, new_AGEMA_signal_15914, mcs1_mcs_mat1_1_mcs_out[31]}), .c ({new_AGEMA_signal_16726, new_AGEMA_signal_16725, new_AGEMA_signal_16724, mcs1_mcs_mat1_1_n123}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U88 ( .a ({new_AGEMA_signal_18235, new_AGEMA_signal_18234, new_AGEMA_signal_18233, mcs1_mcs_mat1_1_mcs_out[19]}), .b ({new_AGEMA_signal_13165, new_AGEMA_signal_13164, new_AGEMA_signal_13163, mcs1_mcs_mat1_1_mcs_out[23]}), .c ({new_AGEMA_signal_18814, new_AGEMA_signal_18813, new_AGEMA_signal_18812, mcs1_mcs_mat1_1_n124}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U87 ( .a ({new_AGEMA_signal_19543, new_AGEMA_signal_19542, new_AGEMA_signal_19541, mcs1_mcs_mat1_1_n122}), .b ({new_AGEMA_signal_15817, new_AGEMA_signal_15816, new_AGEMA_signal_15815, mcs1_mcs_mat1_1_n121}), .c ({temp_next_s3[58], temp_next_s2[58], temp_next_s1[58], temp_next_s0[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U86 ( .a ({new_AGEMA_signal_14602, new_AGEMA_signal_14601, new_AGEMA_signal_14600, mcs1_mcs_mat1_1_mcs_out[26]}), .b ({new_AGEMA_signal_14596, new_AGEMA_signal_14595, new_AGEMA_signal_14594, mcs1_mcs_mat1_1_mcs_out[30]}), .c ({new_AGEMA_signal_15817, new_AGEMA_signal_15816, new_AGEMA_signal_15815, mcs1_mcs_mat1_1_n121}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U85 ( .a ({new_AGEMA_signal_18877, new_AGEMA_signal_18876, new_AGEMA_signal_18875, mcs1_mcs_mat1_1_mcs_out[18]}), .b ({new_AGEMA_signal_14608, new_AGEMA_signal_14607, new_AGEMA_signal_14606, mcs1_mcs_mat1_1_mcs_out[22]}), .c ({new_AGEMA_signal_19543, new_AGEMA_signal_19542, new_AGEMA_signal_19541, mcs1_mcs_mat1_1_n122}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U84 ( .a ({new_AGEMA_signal_20422, new_AGEMA_signal_20421, new_AGEMA_signal_20420, mcs1_mcs_mat1_1_n120}), .b ({new_AGEMA_signal_16729, new_AGEMA_signal_16728, new_AGEMA_signal_16727, mcs1_mcs_mat1_1_n119}), .c ({temp_next_s3[57], temp_next_s2[57], temp_next_s1[57], temp_next_s0[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U83 ( .a ({new_AGEMA_signal_15922, new_AGEMA_signal_15921, new_AGEMA_signal_15920, mcs1_mcs_mat1_1_mcs_out[25]}), .b ({new_AGEMA_signal_13150, new_AGEMA_signal_13149, new_AGEMA_signal_13148, mcs1_mcs_mat1_1_mcs_out[29]}), .c ({new_AGEMA_signal_16729, new_AGEMA_signal_16728, new_AGEMA_signal_16727, mcs1_mcs_mat1_1_n119}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U82 ( .a ({new_AGEMA_signal_19609, new_AGEMA_signal_19608, new_AGEMA_signal_19607, mcs1_mcs_mat1_1_mcs_out[17]}), .b ({new_AGEMA_signal_15925, new_AGEMA_signal_15924, new_AGEMA_signal_15923, mcs1_mcs_mat1_1_mcs_out[21]}), .c ({new_AGEMA_signal_20422, new_AGEMA_signal_20421, new_AGEMA_signal_20420, mcs1_mcs_mat1_1_n120}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U81 ( .a ({new_AGEMA_signal_18817, new_AGEMA_signal_18816, new_AGEMA_signal_18815, mcs1_mcs_mat1_1_n118}), .b ({new_AGEMA_signal_16732, new_AGEMA_signal_16731, new_AGEMA_signal_16730, mcs1_mcs_mat1_1_n117}), .c ({temp_next_s3[56], temp_next_s2[56], temp_next_s1[56], temp_next_s0[56]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U80 ( .a ({new_AGEMA_signal_13162, new_AGEMA_signal_13161, new_AGEMA_signal_13160, mcs1_mcs_mat1_1_mcs_out[24]}), .b ({new_AGEMA_signal_15919, new_AGEMA_signal_15918, new_AGEMA_signal_15917, mcs1_mcs_mat1_1_mcs_out[28]}), .c ({new_AGEMA_signal_16732, new_AGEMA_signal_16731, new_AGEMA_signal_16730, mcs1_mcs_mat1_1_n117}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U79 ( .a ({new_AGEMA_signal_18241, new_AGEMA_signal_18240, new_AGEMA_signal_18239, mcs1_mcs_mat1_1_mcs_out[16]}), .b ({new_AGEMA_signal_13171, new_AGEMA_signal_13170, new_AGEMA_signal_13169, mcs1_mcs_mat1_1_mcs_out[20]}), .c ({new_AGEMA_signal_18817, new_AGEMA_signal_18816, new_AGEMA_signal_18815, mcs1_mcs_mat1_1_n118}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U78 ( .a ({new_AGEMA_signal_16735, new_AGEMA_signal_16734, new_AGEMA_signal_16733, mcs1_mcs_mat1_1_n116}), .b ({new_AGEMA_signal_18820, new_AGEMA_signal_18819, new_AGEMA_signal_18818, mcs1_mcs_mat1_1_n115}), .c ({temp_next_s3[27], temp_next_s2[27], temp_next_s1[27], temp_next_s0[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U77 ( .a ({new_AGEMA_signal_18244, new_AGEMA_signal_18243, new_AGEMA_signal_18242, mcs1_mcs_mat1_1_mcs_out[3]}), .b ({new_AGEMA_signal_15937, new_AGEMA_signal_15936, new_AGEMA_signal_15935, mcs1_mcs_mat1_1_mcs_out[7]}), .c ({new_AGEMA_signal_18820, new_AGEMA_signal_18819, new_AGEMA_signal_18818, mcs1_mcs_mat1_1_n115}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U76 ( .a ({new_AGEMA_signal_10690, new_AGEMA_signal_10689, new_AGEMA_signal_10688, mcs1_mcs_mat1_1_mcs_out[11]}), .b ({new_AGEMA_signal_15928, new_AGEMA_signal_15927, new_AGEMA_signal_15926, mcs1_mcs_mat1_1_mcs_out[15]}), .c ({new_AGEMA_signal_16735, new_AGEMA_signal_16734, new_AGEMA_signal_16733, mcs1_mcs_mat1_1_n116}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U75 ( .a ({new_AGEMA_signal_19552, new_AGEMA_signal_19551, new_AGEMA_signal_19550, mcs1_mcs_mat1_1_n114}), .b ({new_AGEMA_signal_16738, new_AGEMA_signal_16737, new_AGEMA_signal_16736, mcs1_mcs_mat1_1_n113}), .c ({new_AGEMA_signal_20425, new_AGEMA_signal_20424, new_AGEMA_signal_20423, mcs_out[251]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U74 ( .a ({new_AGEMA_signal_15850, new_AGEMA_signal_15849, new_AGEMA_signal_15848, mcs1_mcs_mat1_1_mcs_out[123]}), .b ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_16738, new_AGEMA_signal_16737, new_AGEMA_signal_16736, mcs1_mcs_mat1_1_n113}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U73 ( .a ({new_AGEMA_signal_18856, new_AGEMA_signal_18855, new_AGEMA_signal_18854, mcs1_mcs_mat1_1_mcs_out[115]}), .b ({new_AGEMA_signal_15856, new_AGEMA_signal_15855, new_AGEMA_signal_15854, mcs1_mcs_mat1_1_mcs_out[119]}), .c ({new_AGEMA_signal_19552, new_AGEMA_signal_19551, new_AGEMA_signal_19550, mcs1_mcs_mat1_1_n114}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U72 ( .a ({new_AGEMA_signal_18823, new_AGEMA_signal_18822, new_AGEMA_signal_18821, mcs1_mcs_mat1_1_n112}), .b ({new_AGEMA_signal_13024, new_AGEMA_signal_13023, new_AGEMA_signal_13022, mcs1_mcs_mat1_1_n111}), .c ({new_AGEMA_signal_19555, new_AGEMA_signal_19554, new_AGEMA_signal_19553, mcs_out[250]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U71 ( .a ({new_AGEMA_signal_11590, new_AGEMA_signal_11589, new_AGEMA_signal_11588, mcs1_mcs_mat1_1_mcs_out[122]}), .b ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_13024, new_AGEMA_signal_13023, new_AGEMA_signal_13022, mcs1_mcs_mat1_1_n111}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U70 ( .a ({new_AGEMA_signal_18199, new_AGEMA_signal_18198, new_AGEMA_signal_18197, mcs1_mcs_mat1_1_mcs_out[114]}), .b ({new_AGEMA_signal_15859, new_AGEMA_signal_15858, new_AGEMA_signal_15857, mcs1_mcs_mat1_1_mcs_out[118]}), .c ({new_AGEMA_signal_18823, new_AGEMA_signal_18822, new_AGEMA_signal_18821, mcs1_mcs_mat1_1_n112}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U69 ( .a ({new_AGEMA_signal_15820, new_AGEMA_signal_15819, new_AGEMA_signal_15818, mcs1_mcs_mat1_1_n110}), .b ({new_AGEMA_signal_18826, new_AGEMA_signal_18825, new_AGEMA_signal_18824, mcs1_mcs_mat1_1_n109}), .c ({temp_next_s3[26], temp_next_s2[26], temp_next_s1[26], temp_next_s0[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U68 ( .a ({new_AGEMA_signal_18247, new_AGEMA_signal_18246, new_AGEMA_signal_18245, mcs1_mcs_mat1_1_mcs_out[2]}), .b ({new_AGEMA_signal_13192, new_AGEMA_signal_13191, new_AGEMA_signal_13190, mcs1_mcs_mat1_1_mcs_out[6]}), .c ({new_AGEMA_signal_18826, new_AGEMA_signal_18825, new_AGEMA_signal_18824, mcs1_mcs_mat1_1_n109}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U67 ( .a ({new_AGEMA_signal_14626, new_AGEMA_signal_14625, new_AGEMA_signal_14624, mcs1_mcs_mat1_1_mcs_out[10]}), .b ({new_AGEMA_signal_14617, new_AGEMA_signal_14616, new_AGEMA_signal_14615, mcs1_mcs_mat1_1_mcs_out[14]}), .c ({new_AGEMA_signal_15820, new_AGEMA_signal_15819, new_AGEMA_signal_15818, mcs1_mcs_mat1_1_n110}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U66 ( .a ({new_AGEMA_signal_18184, new_AGEMA_signal_18183, new_AGEMA_signal_18182, mcs1_mcs_mat1_1_n108}), .b ({new_AGEMA_signal_16741, new_AGEMA_signal_16740, new_AGEMA_signal_16739, mcs1_mcs_mat1_1_n107}), .c ({new_AGEMA_signal_18829, new_AGEMA_signal_18828, new_AGEMA_signal_18827, mcs_out[249]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U65 ( .a ({new_AGEMA_signal_15853, new_AGEMA_signal_15852, new_AGEMA_signal_15851, mcs1_mcs_mat1_1_mcs_out[121]}), .b ({new_AGEMA_signal_10588, new_AGEMA_signal_10587, new_AGEMA_signal_10586, mcs1_mcs_mat1_1_mcs_out[125]}), .c ({new_AGEMA_signal_16741, new_AGEMA_signal_16740, new_AGEMA_signal_16739, mcs1_mcs_mat1_1_n107}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U64 ( .a ({new_AGEMA_signal_17485, new_AGEMA_signal_17484, new_AGEMA_signal_17483, mcs1_mcs_mat1_1_mcs_out[113]}), .b ({new_AGEMA_signal_14485, new_AGEMA_signal_14484, new_AGEMA_signal_14483, mcs1_mcs_mat1_1_mcs_out[117]}), .c ({new_AGEMA_signal_18184, new_AGEMA_signal_18183, new_AGEMA_signal_18182, mcs1_mcs_mat1_1_n108}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U63 ( .a ({new_AGEMA_signal_20428, new_AGEMA_signal_20427, new_AGEMA_signal_20426, mcs1_mcs_mat1_1_n106}), .b ({new_AGEMA_signal_15823, new_AGEMA_signal_15822, new_AGEMA_signal_15821, mcs1_mcs_mat1_1_n105}), .c ({new_AGEMA_signal_21172, new_AGEMA_signal_21171, new_AGEMA_signal_21170, mcs_out[248]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U62 ( .a ({new_AGEMA_signal_14476, new_AGEMA_signal_14475, new_AGEMA_signal_14474, mcs1_mcs_mat1_1_mcs_out[120]}), .b ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_15823, new_AGEMA_signal_15822, new_AGEMA_signal_15821, mcs1_mcs_mat1_1_n105}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U61 ( .a ({new_AGEMA_signal_19594, new_AGEMA_signal_19593, new_AGEMA_signal_19592, mcs1_mcs_mat1_1_mcs_out[112]}), .b ({new_AGEMA_signal_13042, new_AGEMA_signal_13041, new_AGEMA_signal_13040, mcs1_mcs_mat1_1_mcs_out[116]}), .c ({new_AGEMA_signal_20428, new_AGEMA_signal_20427, new_AGEMA_signal_20426, mcs1_mcs_mat1_1_n106}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U60 ( .a ({new_AGEMA_signal_15826, new_AGEMA_signal_15825, new_AGEMA_signal_15824, mcs1_mcs_mat1_1_n104}), .b ({new_AGEMA_signal_20431, new_AGEMA_signal_20430, new_AGEMA_signal_20429, mcs1_mcs_mat1_1_n103}), .c ({new_AGEMA_signal_21175, new_AGEMA_signal_21174, new_AGEMA_signal_21173, mcs_out[219]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U59 ( .a ({new_AGEMA_signal_15862, new_AGEMA_signal_15861, new_AGEMA_signal_15860, mcs1_mcs_mat1_1_mcs_out[111]}), .b ({new_AGEMA_signal_19597, new_AGEMA_signal_19596, new_AGEMA_signal_19595, mcs1_mcs_mat1_1_mcs_out[99]}), .c ({new_AGEMA_signal_20431, new_AGEMA_signal_20430, new_AGEMA_signal_20429, mcs1_mcs_mat1_1_n103}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U58 ( .a ({new_AGEMA_signal_14512, new_AGEMA_signal_14511, new_AGEMA_signal_14510, mcs1_mcs_mat1_1_mcs_out[103]}), .b ({new_AGEMA_signal_14500, new_AGEMA_signal_14499, new_AGEMA_signal_14498, mcs1_mcs_mat1_1_mcs_out[107]}), .c ({new_AGEMA_signal_15826, new_AGEMA_signal_15825, new_AGEMA_signal_15824, mcs1_mcs_mat1_1_n104}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U57 ( .a ({new_AGEMA_signal_15829, new_AGEMA_signal_15828, new_AGEMA_signal_15827, mcs1_mcs_mat1_1_n102}), .b ({new_AGEMA_signal_18832, new_AGEMA_signal_18831, new_AGEMA_signal_18830, mcs1_mcs_mat1_1_n101}), .c ({new_AGEMA_signal_19561, new_AGEMA_signal_19560, new_AGEMA_signal_19559, mcs_out[218]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U56 ( .a ({new_AGEMA_signal_15865, new_AGEMA_signal_15864, new_AGEMA_signal_15863, mcs1_mcs_mat1_1_mcs_out[110]}), .b ({new_AGEMA_signal_18208, new_AGEMA_signal_18207, new_AGEMA_signal_18206, mcs1_mcs_mat1_1_mcs_out[98]}), .c ({new_AGEMA_signal_18832, new_AGEMA_signal_18831, new_AGEMA_signal_18830, mcs1_mcs_mat1_1_n101}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U55 ( .a ({new_AGEMA_signal_11617, new_AGEMA_signal_11616, new_AGEMA_signal_11615, mcs1_mcs_mat1_1_mcs_out[102]}), .b ({new_AGEMA_signal_14503, new_AGEMA_signal_14502, new_AGEMA_signal_14501, mcs1_mcs_mat1_1_mcs_out[106]}), .c ({new_AGEMA_signal_15829, new_AGEMA_signal_15828, new_AGEMA_signal_15827, mcs1_mcs_mat1_1_n102}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U54 ( .a ({new_AGEMA_signal_15832, new_AGEMA_signal_15831, new_AGEMA_signal_15830, mcs1_mcs_mat1_1_n100}), .b ({new_AGEMA_signal_17476, new_AGEMA_signal_17475, new_AGEMA_signal_17474, mcs1_mcs_mat1_1_n99}), .c ({new_AGEMA_signal_18187, new_AGEMA_signal_18186, new_AGEMA_signal_18185, mcs_out[217]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U53 ( .a ({new_AGEMA_signal_15868, new_AGEMA_signal_15867, new_AGEMA_signal_15866, mcs1_mcs_mat1_1_mcs_out[109]}), .b ({new_AGEMA_signal_16771, new_AGEMA_signal_16770, new_AGEMA_signal_16769, mcs1_mcs_mat1_1_mcs_out[97]}), .c ({new_AGEMA_signal_17476, new_AGEMA_signal_17475, new_AGEMA_signal_17474, mcs1_mcs_mat1_1_n99}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U52 ( .a ({new_AGEMA_signal_13063, new_AGEMA_signal_13062, new_AGEMA_signal_13061, mcs1_mcs_mat1_1_mcs_out[101]}), .b ({new_AGEMA_signal_14506, new_AGEMA_signal_14505, new_AGEMA_signal_14504, mcs1_mcs_mat1_1_mcs_out[105]}), .c ({new_AGEMA_signal_15832, new_AGEMA_signal_15831, new_AGEMA_signal_15830, mcs1_mcs_mat1_1_n100}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U51 ( .a ({new_AGEMA_signal_16744, new_AGEMA_signal_16743, new_AGEMA_signal_16742, mcs1_mcs_mat1_1_n98}), .b ({new_AGEMA_signal_21679, new_AGEMA_signal_21678, new_AGEMA_signal_21677, mcs1_mcs_mat1_1_n97}), .c ({new_AGEMA_signal_21832, new_AGEMA_signal_21831, new_AGEMA_signal_21830, mcs_out[216]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U50 ( .a ({new_AGEMA_signal_15871, new_AGEMA_signal_15870, new_AGEMA_signal_15869, mcs1_mcs_mat1_1_mcs_out[108]}), .b ({new_AGEMA_signal_21184, new_AGEMA_signal_21183, new_AGEMA_signal_21182, mcs1_mcs_mat1_1_mcs_out[96]}), .c ({new_AGEMA_signal_21679, new_AGEMA_signal_21678, new_AGEMA_signal_21677, mcs1_mcs_mat1_1_n97}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U49 ( .a ({new_AGEMA_signal_14515, new_AGEMA_signal_14514, new_AGEMA_signal_14513, mcs1_mcs_mat1_1_mcs_out[100]}), .b ({new_AGEMA_signal_15874, new_AGEMA_signal_15873, new_AGEMA_signal_15872, mcs1_mcs_mat1_1_mcs_out[104]}), .c ({new_AGEMA_signal_16744, new_AGEMA_signal_16743, new_AGEMA_signal_16742, mcs1_mcs_mat1_1_n98}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U48 ( .a ({new_AGEMA_signal_18835, new_AGEMA_signal_18834, new_AGEMA_signal_18833, mcs1_mcs_mat1_1_n96}), .b ({new_AGEMA_signal_15835, new_AGEMA_signal_15834, new_AGEMA_signal_15833, mcs1_mcs_mat1_1_n95}), .c ({new_AGEMA_signal_19564, new_AGEMA_signal_19563, new_AGEMA_signal_19562, mcs_out[187]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U47 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_14524, new_AGEMA_signal_14523, new_AGEMA_signal_14522, mcs1_mcs_mat1_1_mcs_out[95]}), .c ({new_AGEMA_signal_15835, new_AGEMA_signal_15834, new_AGEMA_signal_15833, mcs1_mcs_mat1_1_n95}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U46 ( .a ({new_AGEMA_signal_18211, new_AGEMA_signal_18210, new_AGEMA_signal_18209, mcs1_mcs_mat1_1_mcs_out[83]}), .b ({new_AGEMA_signal_11638, new_AGEMA_signal_11637, new_AGEMA_signal_11636, mcs1_mcs_mat1_1_mcs_out[87]}), .c ({new_AGEMA_signal_18835, new_AGEMA_signal_18834, new_AGEMA_signal_18833, mcs1_mcs_mat1_1_n96}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U45 ( .a ({new_AGEMA_signal_18838, new_AGEMA_signal_18837, new_AGEMA_signal_18836, mcs1_mcs_mat1_1_n94}), .b ({new_AGEMA_signal_13027, new_AGEMA_signal_13026, new_AGEMA_signal_13025, mcs1_mcs_mat1_1_n93}), .c ({new_AGEMA_signal_19567, new_AGEMA_signal_19566, new_AGEMA_signal_19565, mcs_out[186]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U43 ( .a ({new_AGEMA_signal_18214, new_AGEMA_signal_18213, new_AGEMA_signal_18212, mcs1_mcs_mat1_1_mcs_out[82]}), .b ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_18838, new_AGEMA_signal_18837, new_AGEMA_signal_18836, mcs1_mcs_mat1_1_n94}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U42 ( .a ({new_AGEMA_signal_18841, new_AGEMA_signal_18840, new_AGEMA_signal_18839, mcs1_mcs_mat1_1_n92}), .b ({new_AGEMA_signal_13030, new_AGEMA_signal_13029, new_AGEMA_signal_13028, mcs1_mcs_mat1_1_n91}), .c ({new_AGEMA_signal_19570, new_AGEMA_signal_19569, new_AGEMA_signal_19568, mcs_out[185]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U41 ( .a ({new_AGEMA_signal_10633, new_AGEMA_signal_10632, new_AGEMA_signal_10631, mcs1_mcs_mat1_1_mcs_out[89]}), .b ({new_AGEMA_signal_11632, new_AGEMA_signal_11631, new_AGEMA_signal_11630, mcs1_mcs_mat1_1_mcs_out[93]}), .c ({new_AGEMA_signal_13030, new_AGEMA_signal_13029, new_AGEMA_signal_13028, mcs1_mcs_mat1_1_n91}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U40 ( .a ({new_AGEMA_signal_18217, new_AGEMA_signal_18216, new_AGEMA_signal_18215, mcs1_mcs_mat1_1_mcs_out[81]}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_18841, new_AGEMA_signal_18840, new_AGEMA_signal_18839, mcs1_mcs_mat1_1_n92}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U39 ( .a ({new_AGEMA_signal_19573, new_AGEMA_signal_19572, new_AGEMA_signal_19571, mcs1_mcs_mat1_1_n90}), .b ({new_AGEMA_signal_16747, new_AGEMA_signal_16746, new_AGEMA_signal_16745, mcs1_mcs_mat1_1_n89}), .c ({new_AGEMA_signal_20434, new_AGEMA_signal_20433, new_AGEMA_signal_20432, mcs_out[184]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U38 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_15877, new_AGEMA_signal_15876, new_AGEMA_signal_15875, mcs1_mcs_mat1_1_mcs_out[92]}), .c ({new_AGEMA_signal_16747, new_AGEMA_signal_16746, new_AGEMA_signal_16745, mcs1_mcs_mat1_1_n89}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U37 ( .a ({new_AGEMA_signal_18865, new_AGEMA_signal_18864, new_AGEMA_signal_18863, mcs1_mcs_mat1_1_mcs_out[80]}), .b ({new_AGEMA_signal_13075, new_AGEMA_signal_13074, new_AGEMA_signal_13073, mcs1_mcs_mat1_1_mcs_out[84]}), .c ({new_AGEMA_signal_19573, new_AGEMA_signal_19572, new_AGEMA_signal_19571, mcs1_mcs_mat1_1_n90}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U36 ( .a ({new_AGEMA_signal_19576, new_AGEMA_signal_19575, new_AGEMA_signal_19574, mcs1_mcs_mat1_1_n88}), .b ({new_AGEMA_signal_14458, new_AGEMA_signal_14457, new_AGEMA_signal_14456, mcs1_mcs_mat1_1_n87}), .c ({temp_next_s3[25], temp_next_s2[25], temp_next_s1[25], temp_next_s0[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U35 ( .a ({new_AGEMA_signal_10696, new_AGEMA_signal_10695, new_AGEMA_signal_10694, mcs1_mcs_mat1_1_mcs_out[5]}), .b ({new_AGEMA_signal_13186, new_AGEMA_signal_13185, new_AGEMA_signal_13184, mcs1_mcs_mat1_1_mcs_out[9]}), .c ({new_AGEMA_signal_14458, new_AGEMA_signal_14457, new_AGEMA_signal_14456, mcs1_mcs_mat1_1_n87}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U34 ( .a ({new_AGEMA_signal_14620, new_AGEMA_signal_14619, new_AGEMA_signal_14618, mcs1_mcs_mat1_1_mcs_out[13]}), .b ({new_AGEMA_signal_18883, new_AGEMA_signal_18882, new_AGEMA_signal_18881, mcs1_mcs_mat1_1_mcs_out[1]}), .c ({new_AGEMA_signal_19576, new_AGEMA_signal_19575, new_AGEMA_signal_19574, mcs1_mcs_mat1_1_n88}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U33 ( .a ({new_AGEMA_signal_20440, new_AGEMA_signal_20439, new_AGEMA_signal_20438, mcs1_mcs_mat1_1_n86}), .b ({new_AGEMA_signal_15838, new_AGEMA_signal_15837, new_AGEMA_signal_15836, mcs1_mcs_mat1_1_n85}), .c ({new_AGEMA_signal_21178, new_AGEMA_signal_21177, new_AGEMA_signal_21176, mcs_out[155]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U32 ( .a ({new_AGEMA_signal_11647, new_AGEMA_signal_11646, new_AGEMA_signal_11645, mcs1_mcs_mat1_1_mcs_out[75]}), .b ({new_AGEMA_signal_14533, new_AGEMA_signal_14532, new_AGEMA_signal_14531, mcs1_mcs_mat1_1_mcs_out[79]}), .c ({new_AGEMA_signal_15838, new_AGEMA_signal_15837, new_AGEMA_signal_15836, mcs1_mcs_mat1_1_n85}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U31 ( .a ({new_AGEMA_signal_19600, new_AGEMA_signal_19599, new_AGEMA_signal_19598, mcs1_mcs_mat1_1_mcs_out[67]}), .b ({new_AGEMA_signal_14545, new_AGEMA_signal_14544, new_AGEMA_signal_14543, mcs1_mcs_mat1_1_mcs_out[71]}), .c ({new_AGEMA_signal_20440, new_AGEMA_signal_20439, new_AGEMA_signal_20438, mcs1_mcs_mat1_1_n86}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U30 ( .a ({new_AGEMA_signal_19579, new_AGEMA_signal_19578, new_AGEMA_signal_19577, mcs1_mcs_mat1_1_n84}), .b ({new_AGEMA_signal_16750, new_AGEMA_signal_16749, new_AGEMA_signal_16748, mcs1_mcs_mat1_1_n83}), .c ({new_AGEMA_signal_20443, new_AGEMA_signal_20442, new_AGEMA_signal_20441, mcs_out[154]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U29 ( .a ({new_AGEMA_signal_15883, new_AGEMA_signal_15882, new_AGEMA_signal_15881, mcs1_mcs_mat1_1_mcs_out[74]}), .b ({new_AGEMA_signal_9499, new_AGEMA_signal_9498, new_AGEMA_signal_9497, mcs1_mcs_mat1_1_mcs_out[78]}), .c ({new_AGEMA_signal_16750, new_AGEMA_signal_16749, new_AGEMA_signal_16748, mcs1_mcs_mat1_1_n83}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U28 ( .a ({new_AGEMA_signal_18868, new_AGEMA_signal_18867, new_AGEMA_signal_18866, mcs1_mcs_mat1_1_mcs_out[66]}), .b ({new_AGEMA_signal_15889, new_AGEMA_signal_15888, new_AGEMA_signal_15887, mcs1_mcs_mat1_1_mcs_out[70]}), .c ({new_AGEMA_signal_19579, new_AGEMA_signal_19578, new_AGEMA_signal_19577, mcs1_mcs_mat1_1_n84}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U27 ( .a ({new_AGEMA_signal_18190, new_AGEMA_signal_18189, new_AGEMA_signal_18188, mcs1_mcs_mat1_1_n82}), .b ({new_AGEMA_signal_14461, new_AGEMA_signal_14460, new_AGEMA_signal_14459, mcs1_mcs_mat1_1_n81}), .c ({new_AGEMA_signal_18844, new_AGEMA_signal_18843, new_AGEMA_signal_18842, mcs_out[153]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U26 ( .a ({new_AGEMA_signal_13084, new_AGEMA_signal_13083, new_AGEMA_signal_13082, mcs1_mcs_mat1_1_mcs_out[73]}), .b ({new_AGEMA_signal_11641, new_AGEMA_signal_11640, new_AGEMA_signal_11639, mcs1_mcs_mat1_1_mcs_out[77]}), .c ({new_AGEMA_signal_14461, new_AGEMA_signal_14460, new_AGEMA_signal_14459, mcs1_mcs_mat1_1_n81}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U25 ( .a ({new_AGEMA_signal_17509, new_AGEMA_signal_17508, new_AGEMA_signal_17507, mcs1_mcs_mat1_1_mcs_out[65]}), .b ({new_AGEMA_signal_15892, new_AGEMA_signal_15891, new_AGEMA_signal_15890, mcs1_mcs_mat1_1_mcs_out[69]}), .c ({new_AGEMA_signal_18190, new_AGEMA_signal_18189, new_AGEMA_signal_18188, mcs1_mcs_mat1_1_n82}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U24 ( .a ({new_AGEMA_signal_21181, new_AGEMA_signal_21180, new_AGEMA_signal_21179, mcs1_mcs_mat1_1_n80}), .b ({new_AGEMA_signal_16753, new_AGEMA_signal_16752, new_AGEMA_signal_16751, mcs1_mcs_mat1_1_n79}), .c ({new_AGEMA_signal_21682, new_AGEMA_signal_21681, new_AGEMA_signal_21680, mcs_out[152]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U23 ( .a ({new_AGEMA_signal_15886, new_AGEMA_signal_15885, new_AGEMA_signal_15884, mcs1_mcs_mat1_1_mcs_out[72]}), .b ({new_AGEMA_signal_15880, new_AGEMA_signal_15879, new_AGEMA_signal_15878, mcs1_mcs_mat1_1_mcs_out[76]}), .c ({new_AGEMA_signal_16753, new_AGEMA_signal_16752, new_AGEMA_signal_16751, mcs1_mcs_mat1_1_n79}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U22 ( .a ({new_AGEMA_signal_20455, new_AGEMA_signal_20454, new_AGEMA_signal_20453, mcs1_mcs_mat1_1_mcs_out[64]}), .b ({new_AGEMA_signal_14551, new_AGEMA_signal_14550, new_AGEMA_signal_14549, mcs1_mcs_mat1_1_mcs_out[68]}), .c ({new_AGEMA_signal_21181, new_AGEMA_signal_21180, new_AGEMA_signal_21179, mcs1_mcs_mat1_1_n80}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U21 ( .a ({new_AGEMA_signal_18193, new_AGEMA_signal_18192, new_AGEMA_signal_18191, mcs1_mcs_mat1_1_n78}), .b ({new_AGEMA_signal_15841, new_AGEMA_signal_15840, new_AGEMA_signal_15839, mcs1_mcs_mat1_1_n77}), .c ({temp_next_s3[123], temp_next_s2[123], temp_next_s1[123], temp_next_s0[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U20 ( .a ({new_AGEMA_signal_13108, new_AGEMA_signal_13107, new_AGEMA_signal_13106, mcs1_mcs_mat1_1_mcs_out[59]}), .b ({new_AGEMA_signal_14557, new_AGEMA_signal_14556, new_AGEMA_signal_14555, mcs1_mcs_mat1_1_mcs_out[63]}), .c ({new_AGEMA_signal_15841, new_AGEMA_signal_15840, new_AGEMA_signal_15839, mcs1_mcs_mat1_1_n77}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U19 ( .a ({new_AGEMA_signal_17515, new_AGEMA_signal_17514, new_AGEMA_signal_17513, mcs1_mcs_mat1_1_mcs_out[51]}), .b ({new_AGEMA_signal_14566, new_AGEMA_signal_14565, new_AGEMA_signal_14564, mcs1_mcs_mat1_1_mcs_out[55]}), .c ({new_AGEMA_signal_18193, new_AGEMA_signal_18192, new_AGEMA_signal_18191, mcs1_mcs_mat1_1_n78}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U18 ( .a ({new_AGEMA_signal_16756, new_AGEMA_signal_16755, new_AGEMA_signal_16754, mcs1_mcs_mat1_1_n76}), .b ({new_AGEMA_signal_14464, new_AGEMA_signal_14463, new_AGEMA_signal_14462, mcs1_mcs_mat1_1_n75}), .c ({temp_next_s3[122], temp_next_s2[122], temp_next_s1[122], temp_next_s0[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U17 ( .a ({new_AGEMA_signal_11671, new_AGEMA_signal_11670, new_AGEMA_signal_11669, mcs1_mcs_mat1_1_mcs_out[58]}), .b ({new_AGEMA_signal_13099, new_AGEMA_signal_13098, new_AGEMA_signal_13097, mcs1_mcs_mat1_1_mcs_out[62]}), .c ({new_AGEMA_signal_14464, new_AGEMA_signal_14463, new_AGEMA_signal_14462, mcs1_mcs_mat1_1_n75}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U16 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_15898, new_AGEMA_signal_15897, new_AGEMA_signal_15896, mcs1_mcs_mat1_1_mcs_out[54]}), .c ({new_AGEMA_signal_16756, new_AGEMA_signal_16755, new_AGEMA_signal_16754, mcs1_mcs_mat1_1_n76}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U15 ( .a ({new_AGEMA_signal_16759, new_AGEMA_signal_16758, new_AGEMA_signal_16757, mcs1_mcs_mat1_1_n74}), .b ({new_AGEMA_signal_14467, new_AGEMA_signal_14466, new_AGEMA_signal_14465, mcs1_mcs_mat1_1_n73}), .c ({temp_next_s3[121], temp_next_s2[121], temp_next_s1[121], temp_next_s0[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U14 ( .a ({new_AGEMA_signal_13111, new_AGEMA_signal_13110, new_AGEMA_signal_13109, mcs1_mcs_mat1_1_mcs_out[57]}), .b ({new_AGEMA_signal_13102, new_AGEMA_signal_13101, new_AGEMA_signal_13100, mcs1_mcs_mat1_1_mcs_out[61]}), .c ({new_AGEMA_signal_14467, new_AGEMA_signal_14466, new_AGEMA_signal_14465, mcs1_mcs_mat1_1_n73}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U13 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({new_AGEMA_signal_15901, new_AGEMA_signal_15900, new_AGEMA_signal_15899, mcs1_mcs_mat1_1_mcs_out[53]}), .c ({new_AGEMA_signal_16759, new_AGEMA_signal_16758, new_AGEMA_signal_16757, mcs1_mcs_mat1_1_n74}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U12 ( .a ({new_AGEMA_signal_18850, new_AGEMA_signal_18849, new_AGEMA_signal_18848, mcs1_mcs_mat1_1_n72}), .b ({new_AGEMA_signal_16762, new_AGEMA_signal_16761, new_AGEMA_signal_16760, mcs1_mcs_mat1_1_n71}), .c ({temp_next_s3[120], temp_next_s2[120], temp_next_s1[120], temp_next_s0[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U11 ( .a ({new_AGEMA_signal_14563, new_AGEMA_signal_14562, new_AGEMA_signal_14561, mcs1_mcs_mat1_1_mcs_out[56]}), .b ({new_AGEMA_signal_15895, new_AGEMA_signal_15894, new_AGEMA_signal_15893, mcs1_mcs_mat1_1_mcs_out[60]}), .c ({new_AGEMA_signal_16762, new_AGEMA_signal_16761, new_AGEMA_signal_16760, mcs1_mcs_mat1_1_n71}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U10 ( .a ({new_AGEMA_signal_18226, new_AGEMA_signal_18225, new_AGEMA_signal_18224, mcs1_mcs_mat1_1_mcs_out[48]}), .b ({new_AGEMA_signal_14572, new_AGEMA_signal_14571, new_AGEMA_signal_14570, mcs1_mcs_mat1_1_mcs_out[52]}), .c ({new_AGEMA_signal_18850, new_AGEMA_signal_18849, new_AGEMA_signal_18848, mcs1_mcs_mat1_1_n72}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U9 ( .a ({new_AGEMA_signal_19585, new_AGEMA_signal_19584, new_AGEMA_signal_19583, mcs1_mcs_mat1_1_n70}), .b ({new_AGEMA_signal_15844, new_AGEMA_signal_15843, new_AGEMA_signal_15842, mcs1_mcs_mat1_1_n69}), .c ({temp_next_s3[91], temp_next_s2[91], temp_next_s1[91], temp_next_s0[91]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U8 ( .a ({new_AGEMA_signal_14578, new_AGEMA_signal_14577, new_AGEMA_signal_14576, mcs1_mcs_mat1_1_mcs_out[43]}), .b ({new_AGEMA_signal_14575, new_AGEMA_signal_14574, new_AGEMA_signal_14573, mcs1_mcs_mat1_1_mcs_out[47]}), .c ({new_AGEMA_signal_15844, new_AGEMA_signal_15843, new_AGEMA_signal_15842, mcs1_mcs_mat1_1_n69}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U7 ( .a ({new_AGEMA_signal_18874, new_AGEMA_signal_18873, new_AGEMA_signal_18872, mcs1_mcs_mat1_1_mcs_out[35]}), .b ({new_AGEMA_signal_15907, new_AGEMA_signal_15906, new_AGEMA_signal_15905, mcs1_mcs_mat1_1_mcs_out[39]}), .c ({new_AGEMA_signal_19585, new_AGEMA_signal_19584, new_AGEMA_signal_19583, mcs1_mcs_mat1_1_n70}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U6 ( .a ({new_AGEMA_signal_18853, new_AGEMA_signal_18852, new_AGEMA_signal_18851, mcs1_mcs_mat1_1_n68}), .b ({new_AGEMA_signal_15847, new_AGEMA_signal_15846, new_AGEMA_signal_15845, mcs1_mcs_mat1_1_n67}), .c ({temp_next_s3[90], temp_next_s2[90], temp_next_s1[90], temp_next_s0[90]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U5 ( .a ({new_AGEMA_signal_14581, new_AGEMA_signal_14580, new_AGEMA_signal_14579, mcs1_mcs_mat1_1_mcs_out[42]}), .b ({new_AGEMA_signal_10657, new_AGEMA_signal_10656, new_AGEMA_signal_10655, mcs1_mcs_mat1_1_mcs_out[46]}), .c ({new_AGEMA_signal_15847, new_AGEMA_signal_15846, new_AGEMA_signal_15845, mcs1_mcs_mat1_1_n67}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U4 ( .a ({new_AGEMA_signal_18229, new_AGEMA_signal_18228, new_AGEMA_signal_18227, mcs1_mcs_mat1_1_mcs_out[34]}), .b ({new_AGEMA_signal_11710, new_AGEMA_signal_11709, new_AGEMA_signal_11708, mcs1_mcs_mat1_1_mcs_out[38]}), .c ({new_AGEMA_signal_18853, new_AGEMA_signal_18852, new_AGEMA_signal_18851, mcs1_mcs_mat1_1_n68}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U3 ( .a ({new_AGEMA_signal_19591, new_AGEMA_signal_19590, new_AGEMA_signal_19589, mcs1_mcs_mat1_1_n66}), .b ({new_AGEMA_signal_18196, new_AGEMA_signal_18195, new_AGEMA_signal_18194, mcs1_mcs_mat1_1_n65}), .c ({temp_next_s3[24], temp_next_s2[24], temp_next_s1[24], temp_next_s0[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U2 ( .a ({new_AGEMA_signal_17536, new_AGEMA_signal_17535, new_AGEMA_signal_17534, mcs1_mcs_mat1_1_mcs_out[4]}), .b ({new_AGEMA_signal_15934, new_AGEMA_signal_15933, new_AGEMA_signal_15932, mcs1_mcs_mat1_1_mcs_out[8]}), .c ({new_AGEMA_signal_18196, new_AGEMA_signal_18195, new_AGEMA_signal_18194, mcs1_mcs_mat1_1_n65}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_U1 ( .a ({new_AGEMA_signal_18886, new_AGEMA_signal_18885, new_AGEMA_signal_18884, mcs1_mcs_mat1_1_mcs_out[0]}), .b ({new_AGEMA_signal_16795, new_AGEMA_signal_16794, new_AGEMA_signal_16793, mcs1_mcs_mat1_1_mcs_out[12]}), .c ({new_AGEMA_signal_19591, new_AGEMA_signal_19590, new_AGEMA_signal_19589, mcs1_mcs_mat1_1_n66}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_14470, new_AGEMA_signal_14469, new_AGEMA_signal_14468, mcs1_mcs_mat1_1_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_15850, new_AGEMA_signal_15849, new_AGEMA_signal_15848, mcs1_mcs_mat1_1_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_13033, new_AGEMA_signal_13032, new_AGEMA_signal_13031, mcs1_mcs_mat1_1_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_8701, new_AGEMA_signal_8700, new_AGEMA_signal_8699, mcs1_mcs_mat1_1_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_14470, new_AGEMA_signal_14469, new_AGEMA_signal_14468, mcs1_mcs_mat1_1_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_9478, new_AGEMA_signal_9477, new_AGEMA_signal_9476, mcs1_mcs_mat1_1_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_10591, new_AGEMA_signal_10590, new_AGEMA_signal_10589, mcs1_mcs_mat1_1_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_11590, new_AGEMA_signal_11589, new_AGEMA_signal_11588, mcs1_mcs_mat1_1_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_9481, new_AGEMA_signal_9480, new_AGEMA_signal_9479, mcs1_mcs_mat1_1_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .c ({new_AGEMA_signal_10591, new_AGEMA_signal_10590, new_AGEMA_signal_10589, mcs1_mcs_mat1_1_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_14473, new_AGEMA_signal_14472, new_AGEMA_signal_14471, mcs1_mcs_mat1_1_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .c ({new_AGEMA_signal_15853, new_AGEMA_signal_15852, new_AGEMA_signal_15851, mcs1_mcs_mat1_1_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_13033, new_AGEMA_signal_13032, new_AGEMA_signal_13031, mcs1_mcs_mat1_1_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_14473, new_AGEMA_signal_14472, new_AGEMA_signal_14471, mcs1_mcs_mat1_1_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_11593, new_AGEMA_signal_11592, new_AGEMA_signal_11591, mcs1_mcs_mat1_1_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_10594, new_AGEMA_signal_10593, new_AGEMA_signal_10592, mcs1_mcs_mat1_1_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_13033, new_AGEMA_signal_13032, new_AGEMA_signal_13031, mcs1_mcs_mat1_1_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_13036, new_AGEMA_signal_13035, new_AGEMA_signal_13034, mcs1_mcs_mat1_1_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_14476, new_AGEMA_signal_14475, new_AGEMA_signal_14474, mcs1_mcs_mat1_1_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_11593, new_AGEMA_signal_11592, new_AGEMA_signal_11591, mcs1_mcs_mat1_1_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9481, new_AGEMA_signal_9480, new_AGEMA_signal_9479, mcs1_mcs_mat1_1_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_13036, new_AGEMA_signal_13035, new_AGEMA_signal_13034, mcs1_mcs_mat1_1_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192]}), .c ({new_AGEMA_signal_11593, new_AGEMA_signal_11592, new_AGEMA_signal_11591, mcs1_mcs_mat1_1_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198]}), .c ({new_AGEMA_signal_9481, new_AGEMA_signal_9480, new_AGEMA_signal_9479, mcs1_mcs_mat1_1_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204]}), .c ({new_AGEMA_signal_10594, new_AGEMA_signal_10593, new_AGEMA_signal_10592, mcs1_mcs_mat1_1_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_14479, new_AGEMA_signal_14478, new_AGEMA_signal_14477, mcs1_mcs_mat1_1_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .c ({new_AGEMA_signal_15856, new_AGEMA_signal_15855, new_AGEMA_signal_15854, mcs1_mcs_mat1_1_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_13039, new_AGEMA_signal_13038, new_AGEMA_signal_13037, mcs1_mcs_mat1_1_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10603, new_AGEMA_signal_10602, new_AGEMA_signal_10601, mcs1_mcs_mat1_1_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_14479, new_AGEMA_signal_14478, new_AGEMA_signal_14477, mcs1_mcs_mat1_1_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_14482, new_AGEMA_signal_14481, new_AGEMA_signal_14480, mcs1_mcs_mat1_1_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_11599, new_AGEMA_signal_11598, new_AGEMA_signal_11597, mcs1_mcs_mat1_1_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_15859, new_AGEMA_signal_15858, new_AGEMA_signal_15857, mcs1_mcs_mat1_1_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_13039, new_AGEMA_signal_13038, new_AGEMA_signal_13037, mcs1_mcs_mat1_1_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .c ({new_AGEMA_signal_14482, new_AGEMA_signal_14481, new_AGEMA_signal_14480, mcs1_mcs_mat1_1_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_13039, new_AGEMA_signal_13038, new_AGEMA_signal_13037, mcs1_mcs_mat1_1_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_11596, new_AGEMA_signal_11595, new_AGEMA_signal_11594, mcs1_mcs_mat1_1_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_14485, new_AGEMA_signal_14484, new_AGEMA_signal_14483, mcs1_mcs_mat1_1_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_11602, new_AGEMA_signal_11601, new_AGEMA_signal_11600, mcs1_mcs_mat1_1_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, new_AGEMA_signal_9482, mcs1_mcs_mat1_1_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_13039, new_AGEMA_signal_13038, new_AGEMA_signal_13037, mcs1_mcs_mat1_1_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_10600, new_AGEMA_signal_10599, new_AGEMA_signal_10598, mcs1_mcs_mat1_1_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_11599, new_AGEMA_signal_11598, new_AGEMA_signal_11597, mcs1_mcs_mat1_1_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_13042, new_AGEMA_signal_13041, new_AGEMA_signal_13040, mcs1_mcs_mat1_1_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_8704, new_AGEMA_signal_8703, new_AGEMA_signal_8702, mcs1_mcs_mat1_1_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_10603, new_AGEMA_signal_10602, new_AGEMA_signal_10601, mcs1_mcs_mat1_1_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_11599, new_AGEMA_signal_11598, new_AGEMA_signal_11597, mcs1_mcs_mat1_1_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, new_AGEMA_signal_9482, mcs1_mcs_mat1_1_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_10600, new_AGEMA_signal_10599, new_AGEMA_signal_10598, mcs1_mcs_mat1_1_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({new_AGEMA_signal_11602, new_AGEMA_signal_11601, new_AGEMA_signal_11600, mcs1_mcs_mat1_1_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216]}), .c ({new_AGEMA_signal_9484, new_AGEMA_signal_9483, new_AGEMA_signal_9482, mcs1_mcs_mat1_1_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222]}), .c ({new_AGEMA_signal_10603, new_AGEMA_signal_10602, new_AGEMA_signal_10601, mcs1_mcs_mat1_1_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_18202, new_AGEMA_signal_18201, new_AGEMA_signal_18200, mcs1_mcs_mat1_1_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_14488, new_AGEMA_signal_14487, new_AGEMA_signal_14486, mcs1_mcs_mat1_1_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_18856, new_AGEMA_signal_18855, new_AGEMA_signal_18854, mcs1_mcs_mat1_1_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_16765, new_AGEMA_signal_16764, new_AGEMA_signal_16763, mcs1_mcs_mat1_1_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_16768, new_AGEMA_signal_16767, new_AGEMA_signal_16766, mcs1_mcs_mat1_1_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_17485, new_AGEMA_signal_17484, new_AGEMA_signal_17483, mcs1_mcs_mat1_1_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_18205, new_AGEMA_signal_18204, new_AGEMA_signal_18203, mcs1_mcs_mat1_1_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_18859, new_AGEMA_signal_18858, new_AGEMA_signal_18857, mcs1_mcs_mat1_1_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_19594, new_AGEMA_signal_19593, new_AGEMA_signal_19592, mcs1_mcs_mat1_1_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_18202, new_AGEMA_signal_18201, new_AGEMA_signal_18200, mcs1_mcs_mat1_1_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_18859, new_AGEMA_signal_18858, new_AGEMA_signal_18857, mcs1_mcs_mat1_1_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_13045, new_AGEMA_signal_13044, new_AGEMA_signal_13043, mcs1_mcs_mat1_1_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_17491, new_AGEMA_signal_17490, new_AGEMA_signal_17489, mcs1_mcs_mat1_1_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_18202, new_AGEMA_signal_18201, new_AGEMA_signal_18200, mcs1_mcs_mat1_1_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_14491, new_AGEMA_signal_14490, new_AGEMA_signal_14489, mcs1_mcs_mat1_1_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_17488, new_AGEMA_signal_17487, new_AGEMA_signal_17486, mcs1_mcs_mat1_1_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_18205, new_AGEMA_signal_18204, new_AGEMA_signal_18203, mcs1_mcs_mat1_1_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228]}), .c ({new_AGEMA_signal_17491, new_AGEMA_signal_17490, new_AGEMA_signal_17489, mcs1_mcs_mat1_1_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234]}), .c ({new_AGEMA_signal_14491, new_AGEMA_signal_14490, new_AGEMA_signal_14489, mcs1_mcs_mat1_1_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({new_AGEMA_signal_16768, new_AGEMA_signal_16767, new_AGEMA_signal_16766, mcs1_mcs_mat1_1_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({new_AGEMA_signal_14494, new_AGEMA_signal_14493, new_AGEMA_signal_14492, mcs1_mcs_mat1_1_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_15862, new_AGEMA_signal_15861, new_AGEMA_signal_15860, mcs1_mcs_mat1_1_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({new_AGEMA_signal_14497, new_AGEMA_signal_14496, new_AGEMA_signal_14495, mcs1_mcs_mat1_1_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_15865, new_AGEMA_signal_15864, new_AGEMA_signal_15863, mcs1_mcs_mat1_1_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_10606, new_AGEMA_signal_10605, new_AGEMA_signal_10604, mcs1_mcs_mat1_1_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_14494, new_AGEMA_signal_14493, new_AGEMA_signal_14492, mcs1_mcs_mat1_1_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_15868, new_AGEMA_signal_15867, new_AGEMA_signal_15866, mcs1_mcs_mat1_1_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_9487, new_AGEMA_signal_9486, new_AGEMA_signal_9485, mcs1_mcs_mat1_1_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_13048, new_AGEMA_signal_13047, new_AGEMA_signal_13046, mcs1_mcs_mat1_1_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_14494, new_AGEMA_signal_14493, new_AGEMA_signal_14492, mcs1_mcs_mat1_1_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_11605, new_AGEMA_signal_11604, new_AGEMA_signal_11603, mcs1_mcs_mat1_1_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_14497, new_AGEMA_signal_14496, new_AGEMA_signal_14495, mcs1_mcs_mat1_1_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_15871, new_AGEMA_signal_15870, new_AGEMA_signal_15869, mcs1_mcs_mat1_1_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_13051, new_AGEMA_signal_13050, new_AGEMA_signal_13049, mcs1_mcs_mat1_1_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_14497, new_AGEMA_signal_14496, new_AGEMA_signal_14495, mcs1_mcs_mat1_1_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_10606, new_AGEMA_signal_10605, new_AGEMA_signal_10604, mcs1_mcs_mat1_1_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_11608, new_AGEMA_signal_11607, new_AGEMA_signal_11606, mcs1_mcs_mat1_1_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_13051, new_AGEMA_signal_13050, new_AGEMA_signal_13049, mcs1_mcs_mat1_1_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246]}), .c ({new_AGEMA_signal_11608, new_AGEMA_signal_11607, new_AGEMA_signal_11606, mcs1_mcs_mat1_1_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252]}), .c ({new_AGEMA_signal_9487, new_AGEMA_signal_9486, new_AGEMA_signal_9485, mcs1_mcs_mat1_1_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258]}), .c ({new_AGEMA_signal_10606, new_AGEMA_signal_10605, new_AGEMA_signal_10604, mcs1_mcs_mat1_1_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_13057, new_AGEMA_signal_13056, new_AGEMA_signal_13055, mcs1_mcs_mat1_1_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_13054, new_AGEMA_signal_13053, new_AGEMA_signal_13052, mcs1_mcs_mat1_1_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_14500, new_AGEMA_signal_14499, new_AGEMA_signal_14498, mcs1_mcs_mat1_1_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_13054, new_AGEMA_signal_13053, new_AGEMA_signal_13052, mcs1_mcs_mat1_1_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_10609, new_AGEMA_signal_10608, new_AGEMA_signal_10607, mcs1_mcs_mat1_1_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_14503, new_AGEMA_signal_14502, new_AGEMA_signal_14501, mcs1_mcs_mat1_1_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_9490, new_AGEMA_signal_9489, new_AGEMA_signal_9488, mcs1_mcs_mat1_1_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .c ({new_AGEMA_signal_10609, new_AGEMA_signal_10608, new_AGEMA_signal_10607, mcs1_mcs_mat1_1_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({new_AGEMA_signal_13054, new_AGEMA_signal_13053, new_AGEMA_signal_13052, mcs1_mcs_mat1_1_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_14506, new_AGEMA_signal_14505, new_AGEMA_signal_14504, mcs1_mcs_mat1_1_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_11614, new_AGEMA_signal_11613, new_AGEMA_signal_11612, mcs1_mcs_mat1_1_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_8710, new_AGEMA_signal_8709, new_AGEMA_signal_8708, mcs1_mcs_mat1_1_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_13054, new_AGEMA_signal_13053, new_AGEMA_signal_13052, mcs1_mcs_mat1_1_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_14509, new_AGEMA_signal_14508, new_AGEMA_signal_14507, mcs1_mcs_mat1_1_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_15874, new_AGEMA_signal_15873, new_AGEMA_signal_15872, mcs1_mcs_mat1_1_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_13057, new_AGEMA_signal_13056, new_AGEMA_signal_13055, mcs1_mcs_mat1_1_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_11614, new_AGEMA_signal_11613, new_AGEMA_signal_11612, mcs1_mcs_mat1_1_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_14509, new_AGEMA_signal_14508, new_AGEMA_signal_14507, mcs1_mcs_mat1_1_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_11611, new_AGEMA_signal_11610, new_AGEMA_signal_11609, mcs1_mcs_mat1_1_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .c ({new_AGEMA_signal_13057, new_AGEMA_signal_13056, new_AGEMA_signal_13055, mcs1_mcs_mat1_1_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_9490, new_AGEMA_signal_9489, new_AGEMA_signal_9488, mcs1_mcs_mat1_1_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_10612, new_AGEMA_signal_10611, new_AGEMA_signal_10610, mcs1_mcs_mat1_1_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_11611, new_AGEMA_signal_11610, new_AGEMA_signal_11609, mcs1_mcs_mat1_1_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264]}), .c ({new_AGEMA_signal_11614, new_AGEMA_signal_11613, new_AGEMA_signal_11612, mcs1_mcs_mat1_1_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({new_AGEMA_signal_9490, new_AGEMA_signal_9489, new_AGEMA_signal_9488, mcs1_mcs_mat1_1_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276]}), .c ({new_AGEMA_signal_10612, new_AGEMA_signal_10611, new_AGEMA_signal_10610, mcs1_mcs_mat1_1_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_10615, new_AGEMA_signal_10614, new_AGEMA_signal_10613, mcs1_mcs_mat1_1_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_13060, new_AGEMA_signal_13059, new_AGEMA_signal_13058, mcs1_mcs_mat1_1_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_14512, new_AGEMA_signal_14511, new_AGEMA_signal_14510, mcs1_mcs_mat1_1_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_11626, new_AGEMA_signal_11625, new_AGEMA_signal_11624, mcs1_mcs_mat1_1_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_13060, new_AGEMA_signal_13059, new_AGEMA_signal_13058, mcs1_mcs_mat1_1_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_11620, new_AGEMA_signal_11619, new_AGEMA_signal_11618, mcs1_mcs_mat1_1_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_10618, new_AGEMA_signal_10617, new_AGEMA_signal_10616, mcs1_mcs_mat1_1_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_13063, new_AGEMA_signal_13062, new_AGEMA_signal_13061, mcs1_mcs_mat1_1_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_11623, new_AGEMA_signal_11622, new_AGEMA_signal_11621, mcs1_mcs_mat1_1_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_13066, new_AGEMA_signal_13065, new_AGEMA_signal_13064, mcs1_mcs_mat1_1_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_14515, new_AGEMA_signal_14514, new_AGEMA_signal_14513, mcs1_mcs_mat1_1_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8712, new_AGEMA_signal_8711, mcs1_mcs_mat1_1_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_11626, new_AGEMA_signal_11625, new_AGEMA_signal_11624, mcs1_mcs_mat1_1_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_13066, new_AGEMA_signal_13065, new_AGEMA_signal_13064, mcs1_mcs_mat1_1_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_9493, new_AGEMA_signal_9492, new_AGEMA_signal_9491, mcs1_mcs_mat1_1_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .c ({new_AGEMA_signal_11623, new_AGEMA_signal_11622, new_AGEMA_signal_11621, mcs1_mcs_mat1_1_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282]}), .c ({new_AGEMA_signal_11626, new_AGEMA_signal_11625, new_AGEMA_signal_11624, mcs1_mcs_mat1_1_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288]}), .c ({new_AGEMA_signal_9493, new_AGEMA_signal_9492, new_AGEMA_signal_9491, mcs1_mcs_mat1_1_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294]}), .c ({new_AGEMA_signal_10618, new_AGEMA_signal_10617, new_AGEMA_signal_10616, mcs1_mcs_mat1_1_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_20452, new_AGEMA_signal_20451, new_AGEMA_signal_20450, mcs1_mcs_mat1_1_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_16774, new_AGEMA_signal_16773, new_AGEMA_signal_16772, mcs1_mcs_mat1_1_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_21184, new_AGEMA_signal_21183, new_AGEMA_signal_21182, mcs1_mcs_mat1_1_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_19597, new_AGEMA_signal_19596, new_AGEMA_signal_19595, mcs1_mcs_mat1_1_mcs_out[99]}), .b ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .c ({new_AGEMA_signal_20452, new_AGEMA_signal_20451, new_AGEMA_signal_20450, mcs1_mcs_mat1_1_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_18862, new_AGEMA_signal_18861, new_AGEMA_signal_18860, mcs1_mcs_mat1_1_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .c ({new_AGEMA_signal_19597, new_AGEMA_signal_19596, new_AGEMA_signal_19595, mcs1_mcs_mat1_1_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_18208, new_AGEMA_signal_18207, new_AGEMA_signal_18206, mcs1_mcs_mat1_1_mcs_out[98]}), .b ({new_AGEMA_signal_14521, new_AGEMA_signal_14520, new_AGEMA_signal_14519, mcs1_mcs_mat1_1_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_18862, new_AGEMA_signal_18861, new_AGEMA_signal_18860, mcs1_mcs_mat1_1_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_14518, new_AGEMA_signal_14517, new_AGEMA_signal_14516, mcs1_mcs_mat1_1_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_17494, new_AGEMA_signal_17493, new_AGEMA_signal_17492, mcs1_mcs_mat1_1_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_18208, new_AGEMA_signal_18207, new_AGEMA_signal_18206, mcs1_mcs_mat1_1_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({new_AGEMA_signal_17494, new_AGEMA_signal_17493, new_AGEMA_signal_17492, mcs1_mcs_mat1_1_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306]}), .c ({new_AGEMA_signal_14521, new_AGEMA_signal_14520, new_AGEMA_signal_14519, mcs1_mcs_mat1_1_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312]}), .c ({new_AGEMA_signal_16774, new_AGEMA_signal_16773, new_AGEMA_signal_16772, mcs1_mcs_mat1_1_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_13072, new_AGEMA_signal_13071, new_AGEMA_signal_13070, mcs1_mcs_mat1_1_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_14524, new_AGEMA_signal_14523, new_AGEMA_signal_14522, mcs1_mcs_mat1_1_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_10624, new_AGEMA_signal_10623, new_AGEMA_signal_10622, mcs1_mcs_mat1_1_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_10627, new_AGEMA_signal_10626, new_AGEMA_signal_10625, mcs1_mcs_mat1_1_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_11632, new_AGEMA_signal_11631, new_AGEMA_signal_11630, mcs1_mcs_mat1_1_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_14527, new_AGEMA_signal_14526, new_AGEMA_signal_14525, mcs1_mcs_mat1_1_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_9496, new_AGEMA_signal_9495, new_AGEMA_signal_9494, mcs1_mcs_mat1_1_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_15877, new_AGEMA_signal_15876, new_AGEMA_signal_15875, mcs1_mcs_mat1_1_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_13072, new_AGEMA_signal_13071, new_AGEMA_signal_13070, mcs1_mcs_mat1_1_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .c ({new_AGEMA_signal_14527, new_AGEMA_signal_14526, new_AGEMA_signal_14525, mcs1_mcs_mat1_1_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_8716, new_AGEMA_signal_8715, new_AGEMA_signal_8714, mcs1_mcs_mat1_1_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_11635, new_AGEMA_signal_11634, new_AGEMA_signal_11633, mcs1_mcs_mat1_1_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_13072, new_AGEMA_signal_13071, new_AGEMA_signal_13070, mcs1_mcs_mat1_1_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318]}), .c ({new_AGEMA_signal_11635, new_AGEMA_signal_11634, new_AGEMA_signal_11633, mcs1_mcs_mat1_1_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324]}), .c ({new_AGEMA_signal_9496, new_AGEMA_signal_9495, new_AGEMA_signal_9494, mcs1_mcs_mat1_1_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({new_AGEMA_signal_10627, new_AGEMA_signal_10626, new_AGEMA_signal_10625, mcs1_mcs_mat1_1_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_17503, new_AGEMA_signal_17502, new_AGEMA_signal_17501, mcs1_mcs_mat1_1_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_17506, new_AGEMA_signal_17505, new_AGEMA_signal_17504, mcs1_mcs_mat1_1_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_18211, new_AGEMA_signal_18210, new_AGEMA_signal_18209, mcs1_mcs_mat1_1_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_17497, new_AGEMA_signal_17496, new_AGEMA_signal_17495, mcs1_mcs_mat1_1_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_13078, new_AGEMA_signal_13077, new_AGEMA_signal_13076, mcs1_mcs_mat1_1_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_18214, new_AGEMA_signal_18213, new_AGEMA_signal_18212, mcs1_mcs_mat1_1_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_16777, new_AGEMA_signal_16776, new_AGEMA_signal_16775, mcs1_mcs_mat1_1_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_17497, new_AGEMA_signal_17496, new_AGEMA_signal_17495, mcs1_mcs_mat1_1_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_17500, new_AGEMA_signal_17499, new_AGEMA_signal_17498, mcs1_mcs_mat1_1_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_18217, new_AGEMA_signal_18216, new_AGEMA_signal_18215, mcs1_mcs_mat1_1_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_14530, new_AGEMA_signal_14529, new_AGEMA_signal_14528, mcs1_mcs_mat1_1_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_16777, new_AGEMA_signal_16776, new_AGEMA_signal_16775, mcs1_mcs_mat1_1_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_17500, new_AGEMA_signal_17499, new_AGEMA_signal_17498, mcs1_mcs_mat1_1_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_18220, new_AGEMA_signal_18219, new_AGEMA_signal_18218, mcs1_mcs_mat1_1_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .c ({new_AGEMA_signal_18865, new_AGEMA_signal_18864, new_AGEMA_signal_18863, mcs1_mcs_mat1_1_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_17503, new_AGEMA_signal_17502, new_AGEMA_signal_17501, mcs1_mcs_mat1_1_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_14530, new_AGEMA_signal_14529, new_AGEMA_signal_14528, mcs1_mcs_mat1_1_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_18220, new_AGEMA_signal_18219, new_AGEMA_signal_18218, mcs1_mcs_mat1_1_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336]}), .c ({new_AGEMA_signal_17506, new_AGEMA_signal_17505, new_AGEMA_signal_17504, mcs1_mcs_mat1_1_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342]}), .c ({new_AGEMA_signal_14530, new_AGEMA_signal_14529, new_AGEMA_signal_14528, mcs1_mcs_mat1_1_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348]}), .c ({new_AGEMA_signal_16777, new_AGEMA_signal_16776, new_AGEMA_signal_16775, mcs1_mcs_mat1_1_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_13081, new_AGEMA_signal_13080, new_AGEMA_signal_13079, mcs1_mcs_mat1_1_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_14533, new_AGEMA_signal_14532, new_AGEMA_signal_14531, mcs1_mcs_mat1_1_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_10636, new_AGEMA_signal_10635, new_AGEMA_signal_10634, mcs1_mcs_mat1_1_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_11641, new_AGEMA_signal_11640, new_AGEMA_signal_11639, mcs1_mcs_mat1_1_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_14536, new_AGEMA_signal_14535, new_AGEMA_signal_14534, mcs1_mcs_mat1_1_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_9502, new_AGEMA_signal_9501, new_AGEMA_signal_9500, mcs1_mcs_mat1_1_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_15880, new_AGEMA_signal_15879, new_AGEMA_signal_15878, mcs1_mcs_mat1_1_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_13081, new_AGEMA_signal_13080, new_AGEMA_signal_13079, mcs1_mcs_mat1_1_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .c ({new_AGEMA_signal_14536, new_AGEMA_signal_14535, new_AGEMA_signal_14534, mcs1_mcs_mat1_1_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_8719, new_AGEMA_signal_8718, new_AGEMA_signal_8717, mcs1_mcs_mat1_1_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_11644, new_AGEMA_signal_11643, new_AGEMA_signal_11642, mcs1_mcs_mat1_1_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_13081, new_AGEMA_signal_13080, new_AGEMA_signal_13079, mcs1_mcs_mat1_1_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354]}), .c ({new_AGEMA_signal_11644, new_AGEMA_signal_11643, new_AGEMA_signal_11642, mcs1_mcs_mat1_1_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({new_AGEMA_signal_9502, new_AGEMA_signal_9501, new_AGEMA_signal_9500, mcs1_mcs_mat1_1_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366]}), .c ({new_AGEMA_signal_10636, new_AGEMA_signal_10635, new_AGEMA_signal_10634, mcs1_mcs_mat1_1_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_14539, new_AGEMA_signal_14538, new_AGEMA_signal_14537, mcs1_mcs_mat1_1_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_15883, new_AGEMA_signal_15882, new_AGEMA_signal_15881, mcs1_mcs_mat1_1_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_13087, new_AGEMA_signal_13086, new_AGEMA_signal_13085, mcs1_mcs_mat1_1_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_11650, new_AGEMA_signal_11649, new_AGEMA_signal_11648, mcs1_mcs_mat1_1_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_14539, new_AGEMA_signal_14538, new_AGEMA_signal_14537, mcs1_mcs_mat1_1_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, new_AGEMA_signal_10286, mcs1_mcs_mat1_1_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_11647, new_AGEMA_signal_11646, new_AGEMA_signal_11645, mcs1_mcs_mat1_1_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_11650, new_AGEMA_signal_11649, new_AGEMA_signal_11648, mcs1_mcs_mat1_1_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, new_AGEMA_signal_10286, mcs1_mcs_mat1_1_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_13084, new_AGEMA_signal_13083, new_AGEMA_signal_13082, mcs1_mcs_mat1_1_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, new_AGEMA_signal_9503, mcs1_mcs_mat1_1_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_9508, new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_1_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_10288, new_AGEMA_signal_10287, new_AGEMA_signal_10286, mcs1_mcs_mat1_1_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_10639, new_AGEMA_signal_10638, new_AGEMA_signal_10637, mcs1_mcs_mat1_1_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .c ({new_AGEMA_signal_11650, new_AGEMA_signal_11649, new_AGEMA_signal_11648, mcs1_mcs_mat1_1_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_14542, new_AGEMA_signal_14541, new_AGEMA_signal_14540, mcs1_mcs_mat1_1_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_9505, new_AGEMA_signal_9504, new_AGEMA_signal_9503, mcs1_mcs_mat1_1_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_15886, new_AGEMA_signal_15885, new_AGEMA_signal_15884, mcs1_mcs_mat1_1_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_13087, new_AGEMA_signal_13086, new_AGEMA_signal_13085, mcs1_mcs_mat1_1_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_10639, new_AGEMA_signal_10638, new_AGEMA_signal_10637, mcs1_mcs_mat1_1_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_14542, new_AGEMA_signal_14541, new_AGEMA_signal_14540, mcs1_mcs_mat1_1_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .b ({new_AGEMA_signal_11653, new_AGEMA_signal_11652, new_AGEMA_signal_11651, mcs1_mcs_mat1_1_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_13087, new_AGEMA_signal_13086, new_AGEMA_signal_13085, mcs1_mcs_mat1_1_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372]}), .c ({new_AGEMA_signal_11653, new_AGEMA_signal_11652, new_AGEMA_signal_11651, mcs1_mcs_mat1_1_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378]}), .c ({new_AGEMA_signal_9508, new_AGEMA_signal_9507, new_AGEMA_signal_9506, mcs1_mcs_mat1_1_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384]}), .c ({new_AGEMA_signal_10639, new_AGEMA_signal_10638, new_AGEMA_signal_10637, mcs1_mcs_mat1_1_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_13090, new_AGEMA_signal_13089, new_AGEMA_signal_13088, mcs1_mcs_mat1_1_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_10642, new_AGEMA_signal_10641, new_AGEMA_signal_10640, mcs1_mcs_mat1_1_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_14545, new_AGEMA_signal_14544, new_AGEMA_signal_14543, mcs1_mcs_mat1_1_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_11659, new_AGEMA_signal_11658, new_AGEMA_signal_11657, mcs1_mcs_mat1_1_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_14548, new_AGEMA_signal_14547, new_AGEMA_signal_14546, mcs1_mcs_mat1_1_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_15889, new_AGEMA_signal_15888, new_AGEMA_signal_15887, mcs1_mcs_mat1_1_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_13090, new_AGEMA_signal_13089, new_AGEMA_signal_13088, mcs1_mcs_mat1_1_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_14548, new_AGEMA_signal_14547, new_AGEMA_signal_14546, mcs1_mcs_mat1_1_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_15892, new_AGEMA_signal_15891, new_AGEMA_signal_15890, mcs1_mcs_mat1_1_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_10642, new_AGEMA_signal_10641, new_AGEMA_signal_10640, mcs1_mcs_mat1_1_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_13093, new_AGEMA_signal_13092, new_AGEMA_signal_13091, mcs1_mcs_mat1_1_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_14548, new_AGEMA_signal_14547, new_AGEMA_signal_14546, mcs1_mcs_mat1_1_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, new_AGEMA_signal_9509, mcs1_mcs_mat1_1_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_10642, new_AGEMA_signal_10641, new_AGEMA_signal_10640, mcs1_mcs_mat1_1_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_11656, new_AGEMA_signal_11655, new_AGEMA_signal_11654, mcs1_mcs_mat1_1_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .c ({new_AGEMA_signal_13090, new_AGEMA_signal_13089, new_AGEMA_signal_13088, mcs1_mcs_mat1_1_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_10645, new_AGEMA_signal_10644, new_AGEMA_signal_10643, mcs1_mcs_mat1_1_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8725, new_AGEMA_signal_8724, new_AGEMA_signal_8723, mcs1_mcs_mat1_1_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_11656, new_AGEMA_signal_11655, new_AGEMA_signal_11654, mcs1_mcs_mat1_1_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_13093, new_AGEMA_signal_13092, new_AGEMA_signal_13091, mcs1_mcs_mat1_1_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_11659, new_AGEMA_signal_11658, new_AGEMA_signal_11657, mcs1_mcs_mat1_1_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_14551, new_AGEMA_signal_14550, new_AGEMA_signal_14549, mcs1_mcs_mat1_1_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_10645, new_AGEMA_signal_10644, new_AGEMA_signal_10643, mcs1_mcs_mat1_1_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_11659, new_AGEMA_signal_11658, new_AGEMA_signal_11657, mcs1_mcs_mat1_1_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({new_AGEMA_signal_11662, new_AGEMA_signal_11661, new_AGEMA_signal_11660, mcs1_mcs_mat1_1_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_13093, new_AGEMA_signal_13092, new_AGEMA_signal_13091, mcs1_mcs_mat1_1_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .c ({new_AGEMA_signal_11662, new_AGEMA_signal_11661, new_AGEMA_signal_11660, mcs1_mcs_mat1_1_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396]}), .c ({new_AGEMA_signal_9511, new_AGEMA_signal_9510, new_AGEMA_signal_9509, mcs1_mcs_mat1_1_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402]}), .c ({new_AGEMA_signal_10645, new_AGEMA_signal_10644, new_AGEMA_signal_10643, mcs1_mcs_mat1_1_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_18871, new_AGEMA_signal_18870, new_AGEMA_signal_18869, mcs1_mcs_mat1_1_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .c ({new_AGEMA_signal_19600, new_AGEMA_signal_19599, new_AGEMA_signal_19598, mcs1_mcs_mat1_1_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({new_AGEMA_signal_18223, new_AGEMA_signal_18222, new_AGEMA_signal_18221, mcs1_mcs_mat1_1_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_18868, new_AGEMA_signal_18867, new_AGEMA_signal_18866, mcs1_mcs_mat1_1_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_19603, new_AGEMA_signal_19602, new_AGEMA_signal_19601, mcs1_mcs_mat1_1_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_16780, new_AGEMA_signal_16779, new_AGEMA_signal_16778, mcs1_mcs_mat1_1_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_20455, new_AGEMA_signal_20454, new_AGEMA_signal_20453, mcs1_mcs_mat1_1_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_18871, new_AGEMA_signal_18870, new_AGEMA_signal_18869, mcs1_mcs_mat1_1_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .c ({new_AGEMA_signal_19603, new_AGEMA_signal_19602, new_AGEMA_signal_19601, mcs1_mcs_mat1_1_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_14554, new_AGEMA_signal_14553, new_AGEMA_signal_14552, mcs1_mcs_mat1_1_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_18223, new_AGEMA_signal_18222, new_AGEMA_signal_18221, mcs1_mcs_mat1_1_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_18871, new_AGEMA_signal_18870, new_AGEMA_signal_18869, mcs1_mcs_mat1_1_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_13096, new_AGEMA_signal_13095, new_AGEMA_signal_13094, mcs1_mcs_mat1_1_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_17512, new_AGEMA_signal_17511, new_AGEMA_signal_17510, mcs1_mcs_mat1_1_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_18223, new_AGEMA_signal_18222, new_AGEMA_signal_18221, mcs1_mcs_mat1_1_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408]}), .c ({new_AGEMA_signal_17512, new_AGEMA_signal_17511, new_AGEMA_signal_17510, mcs1_mcs_mat1_1_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414]}), .c ({new_AGEMA_signal_14554, new_AGEMA_signal_14553, new_AGEMA_signal_14552, mcs1_mcs_mat1_1_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({new_AGEMA_signal_16780, new_AGEMA_signal_16779, new_AGEMA_signal_16778, mcs1_mcs_mat1_1_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_13105, new_AGEMA_signal_13104, new_AGEMA_signal_13103, mcs1_mcs_mat1_1_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_10648, new_AGEMA_signal_10647, new_AGEMA_signal_10646, mcs1_mcs_mat1_1_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_14557, new_AGEMA_signal_14556, new_AGEMA_signal_14555, mcs1_mcs_mat1_1_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_9514, new_AGEMA_signal_9513, new_AGEMA_signal_9512, mcs1_mcs_mat1_1_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_11665, new_AGEMA_signal_11664, new_AGEMA_signal_11663, mcs1_mcs_mat1_1_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_13099, new_AGEMA_signal_13098, new_AGEMA_signal_13097, mcs1_mcs_mat1_1_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({new_AGEMA_signal_11668, new_AGEMA_signal_11667, new_AGEMA_signal_11666, mcs1_mcs_mat1_1_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_13102, new_AGEMA_signal_13101, new_AGEMA_signal_13100, mcs1_mcs_mat1_1_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426]}), .c ({new_AGEMA_signal_11668, new_AGEMA_signal_11667, new_AGEMA_signal_11666, mcs1_mcs_mat1_1_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432]}), .c ({new_AGEMA_signal_9514, new_AGEMA_signal_9513, new_AGEMA_signal_9512, mcs1_mcs_mat1_1_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438]}), .c ({new_AGEMA_signal_10648, new_AGEMA_signal_10647, new_AGEMA_signal_10646, mcs1_mcs_mat1_1_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_9520, new_AGEMA_signal_9519, new_AGEMA_signal_9518, mcs1_mcs_mat1_1_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_10651, new_AGEMA_signal_10650, new_AGEMA_signal_10649, mcs1_mcs_mat1_1_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_11671, new_AGEMA_signal_11670, new_AGEMA_signal_11669, mcs1_mcs_mat1_1_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_9523, new_AGEMA_signal_9522, new_AGEMA_signal_9521, mcs1_mcs_mat1_1_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_11674, new_AGEMA_signal_11673, new_AGEMA_signal_11672, mcs1_mcs_mat1_1_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_13111, new_AGEMA_signal_13110, new_AGEMA_signal_13109, mcs1_mcs_mat1_1_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_13114, new_AGEMA_signal_13113, new_AGEMA_signal_13112, mcs1_mcs_mat1_1_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_11677, new_AGEMA_signal_11676, new_AGEMA_signal_11675, mcs1_mcs_mat1_1_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_14563, new_AGEMA_signal_14562, new_AGEMA_signal_14561, mcs1_mcs_mat1_1_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_11680, new_AGEMA_signal_11679, new_AGEMA_signal_11678, mcs1_mcs_mat1_1_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_13114, new_AGEMA_signal_13113, new_AGEMA_signal_13112, mcs1_mcs_mat1_1_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444]}), .c ({new_AGEMA_signal_11680, new_AGEMA_signal_11679, new_AGEMA_signal_11678, mcs1_mcs_mat1_1_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .c ({new_AGEMA_signal_9523, new_AGEMA_signal_9522, new_AGEMA_signal_9521, mcs1_mcs_mat1_1_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456]}), .c ({new_AGEMA_signal_10651, new_AGEMA_signal_10650, new_AGEMA_signal_10649, mcs1_mcs_mat1_1_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_11686, new_AGEMA_signal_11685, new_AGEMA_signal_11684, mcs1_mcs_mat1_1_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_13117, new_AGEMA_signal_13116, new_AGEMA_signal_13115, mcs1_mcs_mat1_1_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_14566, new_AGEMA_signal_14565, new_AGEMA_signal_14564, mcs1_mcs_mat1_1_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_14569, new_AGEMA_signal_14568, new_AGEMA_signal_14567, mcs1_mcs_mat1_1_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_11683, new_AGEMA_signal_11682, new_AGEMA_signal_11681, mcs1_mcs_mat1_1_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_15898, new_AGEMA_signal_15897, new_AGEMA_signal_15896, mcs1_mcs_mat1_1_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_10654, new_AGEMA_signal_10653, new_AGEMA_signal_10652, mcs1_mcs_mat1_1_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_11683, new_AGEMA_signal_11682, new_AGEMA_signal_11681, mcs1_mcs_mat1_1_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({new_AGEMA_signal_14569, new_AGEMA_signal_14568, new_AGEMA_signal_14567, mcs1_mcs_mat1_1_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_15901, new_AGEMA_signal_15900, new_AGEMA_signal_15899, mcs1_mcs_mat1_1_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_8734, new_AGEMA_signal_8733, new_AGEMA_signal_8732, mcs1_mcs_mat1_1_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_13117, new_AGEMA_signal_13116, new_AGEMA_signal_13115, mcs1_mcs_mat1_1_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_14569, new_AGEMA_signal_14568, new_AGEMA_signal_14567, mcs1_mcs_mat1_1_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_9526, new_AGEMA_signal_9525, new_AGEMA_signal_9524, mcs1_mcs_mat1_1_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_11692, new_AGEMA_signal_11691, new_AGEMA_signal_11690, mcs1_mcs_mat1_1_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_13117, new_AGEMA_signal_13116, new_AGEMA_signal_13115, mcs1_mcs_mat1_1_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_11689, new_AGEMA_signal_11688, new_AGEMA_signal_11687, mcs1_mcs_mat1_1_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_13120, new_AGEMA_signal_13119, new_AGEMA_signal_13118, mcs1_mcs_mat1_1_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_14572, new_AGEMA_signal_14571, new_AGEMA_signal_14570, mcs1_mcs_mat1_1_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_11686, new_AGEMA_signal_11685, new_AGEMA_signal_11684, mcs1_mcs_mat1_1_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_9526, new_AGEMA_signal_9525, new_AGEMA_signal_9524, mcs1_mcs_mat1_1_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_13120, new_AGEMA_signal_13119, new_AGEMA_signal_13118, mcs1_mcs_mat1_1_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_10654, new_AGEMA_signal_10653, new_AGEMA_signal_10652, mcs1_mcs_mat1_1_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_11686, new_AGEMA_signal_11685, new_AGEMA_signal_11684, mcs1_mcs_mat1_1_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462]}), .c ({new_AGEMA_signal_11692, new_AGEMA_signal_11691, new_AGEMA_signal_11690, mcs1_mcs_mat1_1_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468]}), .c ({new_AGEMA_signal_9526, new_AGEMA_signal_9525, new_AGEMA_signal_9524, mcs1_mcs_mat1_1_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474]}), .c ({new_AGEMA_signal_10654, new_AGEMA_signal_10653, new_AGEMA_signal_10652, mcs1_mcs_mat1_1_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_10660, new_AGEMA_signal_10659, new_AGEMA_signal_10658, mcs1_mcs_mat1_1_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_11695, new_AGEMA_signal_11694, new_AGEMA_signal_11693, mcs1_mcs_mat1_1_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_15904, new_AGEMA_signal_15903, new_AGEMA_signal_15902, mcs1_mcs_mat1_1_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_9529, new_AGEMA_signal_9528, new_AGEMA_signal_9527, mcs1_mcs_mat1_1_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_16783, new_AGEMA_signal_16782, new_AGEMA_signal_16781, mcs1_mcs_mat1_1_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_14575, new_AGEMA_signal_14574, new_AGEMA_signal_14573, mcs1_mcs_mat1_1_mcs_out[47]}), .b ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .c ({new_AGEMA_signal_15904, new_AGEMA_signal_15903, new_AGEMA_signal_15902, mcs1_mcs_mat1_1_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_13123, new_AGEMA_signal_13122, new_AGEMA_signal_13121, mcs1_mcs_mat1_1_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .c ({new_AGEMA_signal_14575, new_AGEMA_signal_14574, new_AGEMA_signal_14573, mcs1_mcs_mat1_1_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8736, new_AGEMA_signal_8735, mcs1_mcs_mat1_1_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_11698, new_AGEMA_signal_11697, new_AGEMA_signal_11696, mcs1_mcs_mat1_1_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_13123, new_AGEMA_signal_13122, new_AGEMA_signal_13121, mcs1_mcs_mat1_1_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({new_AGEMA_signal_11698, new_AGEMA_signal_11697, new_AGEMA_signal_11696, mcs1_mcs_mat1_1_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486]}), .c ({new_AGEMA_signal_9529, new_AGEMA_signal_9528, new_AGEMA_signal_9527, mcs1_mcs_mat1_1_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492]}), .c ({new_AGEMA_signal_10660, new_AGEMA_signal_10659, new_AGEMA_signal_10658, mcs1_mcs_mat1_1_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_13126, new_AGEMA_signal_13125, new_AGEMA_signal_13124, mcs1_mcs_mat1_1_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_10663, new_AGEMA_signal_10662, new_AGEMA_signal_10661, mcs1_mcs_mat1_1_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_14578, new_AGEMA_signal_14577, new_AGEMA_signal_14576, mcs1_mcs_mat1_1_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_11701, new_AGEMA_signal_11700, new_AGEMA_signal_11699, mcs1_mcs_mat1_1_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9532, new_AGEMA_signal_9531, new_AGEMA_signal_9530, mcs1_mcs_mat1_1_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_13126, new_AGEMA_signal_13125, new_AGEMA_signal_13124, mcs1_mcs_mat1_1_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_13129, new_AGEMA_signal_13128, new_AGEMA_signal_13127, mcs1_mcs_mat1_1_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_11707, new_AGEMA_signal_11706, new_AGEMA_signal_11705, mcs1_mcs_mat1_1_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_14581, new_AGEMA_signal_14580, new_AGEMA_signal_14579, mcs1_mcs_mat1_1_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_13132, new_AGEMA_signal_13131, new_AGEMA_signal_13130, mcs1_mcs_mat1_1_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_8740, new_AGEMA_signal_8739, new_AGEMA_signal_8738, mcs1_mcs_mat1_1_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_14584, new_AGEMA_signal_14583, new_AGEMA_signal_14582, mcs1_mcs_mat1_1_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_11701, new_AGEMA_signal_11700, new_AGEMA_signal_11699, mcs1_mcs_mat1_1_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_10666, new_AGEMA_signal_10665, new_AGEMA_signal_10664, mcs1_mcs_mat1_1_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_13132, new_AGEMA_signal_13131, new_AGEMA_signal_13130, mcs1_mcs_mat1_1_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_11704, new_AGEMA_signal_11703, new_AGEMA_signal_11702, mcs1_mcs_mat1_1_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_10666, new_AGEMA_signal_10665, new_AGEMA_signal_10664, mcs1_mcs_mat1_1_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_13135, new_AGEMA_signal_13134, new_AGEMA_signal_13133, mcs1_mcs_mat1_1_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498]}), .c ({new_AGEMA_signal_11707, new_AGEMA_signal_11706, new_AGEMA_signal_11705, mcs1_mcs_mat1_1_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504]}), .c ({new_AGEMA_signal_9532, new_AGEMA_signal_9531, new_AGEMA_signal_9530, mcs1_mcs_mat1_1_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .c ({new_AGEMA_signal_10666, new_AGEMA_signal_10665, new_AGEMA_signal_10664, mcs1_mcs_mat1_1_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_14587, new_AGEMA_signal_14586, new_AGEMA_signal_14585, mcs1_mcs_mat1_1_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_8743, new_AGEMA_signal_8742, new_AGEMA_signal_8741, mcs1_mcs_mat1_1_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_15907, new_AGEMA_signal_15906, new_AGEMA_signal_15905, mcs1_mcs_mat1_1_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_10672, new_AGEMA_signal_10671, new_AGEMA_signal_10670, mcs1_mcs_mat1_1_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_10669, new_AGEMA_signal_10668, new_AGEMA_signal_10667, mcs1_mcs_mat1_1_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_11710, new_AGEMA_signal_11709, new_AGEMA_signal_11708, mcs1_mcs_mat1_1_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({new_AGEMA_signal_14587, new_AGEMA_signal_14586, new_AGEMA_signal_14585, mcs1_mcs_mat1_1_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_15910, new_AGEMA_signal_15909, new_AGEMA_signal_15908, mcs1_mcs_mat1_1_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_11713, new_AGEMA_signal_11712, new_AGEMA_signal_11711, mcs1_mcs_mat1_1_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_13138, new_AGEMA_signal_13137, new_AGEMA_signal_13136, mcs1_mcs_mat1_1_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_14587, new_AGEMA_signal_14586, new_AGEMA_signal_14585, mcs1_mcs_mat1_1_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_11716, new_AGEMA_signal_11715, new_AGEMA_signal_11714, mcs1_mcs_mat1_1_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_10675, new_AGEMA_signal_10674, new_AGEMA_signal_10673, mcs1_mcs_mat1_1_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_13138, new_AGEMA_signal_13137, new_AGEMA_signal_13136, mcs1_mcs_mat1_1_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_11716, new_AGEMA_signal_11715, new_AGEMA_signal_11714, mcs1_mcs_mat1_1_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_10672, new_AGEMA_signal_10671, new_AGEMA_signal_10670, mcs1_mcs_mat1_1_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_13141, new_AGEMA_signal_13140, new_AGEMA_signal_13139, mcs1_mcs_mat1_1_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .b ({new_AGEMA_signal_10291, new_AGEMA_signal_10290, new_AGEMA_signal_10289, mcs1_mcs_mat1_1_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_10672, new_AGEMA_signal_10671, new_AGEMA_signal_10670, mcs1_mcs_mat1_1_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({new_AGEMA_signal_9535, new_AGEMA_signal_9534, new_AGEMA_signal_9533, mcs1_mcs_mat1_1_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_10291, new_AGEMA_signal_10290, new_AGEMA_signal_10289, mcs1_mcs_mat1_1_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516]}), .c ({new_AGEMA_signal_11716, new_AGEMA_signal_11715, new_AGEMA_signal_11714, mcs1_mcs_mat1_1_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522]}), .c ({new_AGEMA_signal_9535, new_AGEMA_signal_9534, new_AGEMA_signal_9533, mcs1_mcs_mat1_1_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528]}), .c ({new_AGEMA_signal_10675, new_AGEMA_signal_10674, new_AGEMA_signal_10673, mcs1_mcs_mat1_1_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_17518, new_AGEMA_signal_17517, new_AGEMA_signal_17516, mcs1_mcs_mat1_1_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_16786, new_AGEMA_signal_16785, new_AGEMA_signal_16784, mcs1_mcs_mat1_1_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_18229, new_AGEMA_signal_18228, new_AGEMA_signal_18227, mcs1_mcs_mat1_1_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_14590, new_AGEMA_signal_14589, new_AGEMA_signal_14588, mcs1_mcs_mat1_1_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_15913, new_AGEMA_signal_15912, new_AGEMA_signal_15911, mcs1_mcs_mat1_1_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_19606, new_AGEMA_signal_19605, new_AGEMA_signal_19604, mcs1_mcs_mat1_1_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_17521, new_AGEMA_signal_17520, new_AGEMA_signal_17519, mcs1_mcs_mat1_1_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_20458, new_AGEMA_signal_20457, new_AGEMA_signal_20456, mcs1_mcs_mat1_1_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534]}), .c ({new_AGEMA_signal_17521, new_AGEMA_signal_17520, new_AGEMA_signal_17519, mcs1_mcs_mat1_1_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({new_AGEMA_signal_14590, new_AGEMA_signal_14589, new_AGEMA_signal_14588, mcs1_mcs_mat1_1_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546]}), .c ({new_AGEMA_signal_16786, new_AGEMA_signal_16785, new_AGEMA_signal_16784, mcs1_mcs_mat1_1_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_14593, new_AGEMA_signal_14592, new_AGEMA_signal_14591, mcs1_mcs_mat1_1_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_13147, new_AGEMA_signal_13146, new_AGEMA_signal_13145, mcs1_mcs_mat1_1_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_15916, new_AGEMA_signal_15915, new_AGEMA_signal_15914, mcs1_mcs_mat1_1_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_9541, new_AGEMA_signal_9540, new_AGEMA_signal_9539, mcs1_mcs_mat1_1_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_13150, new_AGEMA_signal_13149, new_AGEMA_signal_13148, mcs1_mcs_mat1_1_mcs_out[29]}), .c ({new_AGEMA_signal_14593, new_AGEMA_signal_14592, new_AGEMA_signal_14591, mcs1_mcs_mat1_1_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_9538, new_AGEMA_signal_9537, new_AGEMA_signal_9536, mcs1_mcs_mat1_1_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_13147, new_AGEMA_signal_13146, new_AGEMA_signal_13145, mcs1_mcs_mat1_1_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_14596, new_AGEMA_signal_14595, new_AGEMA_signal_14594, mcs1_mcs_mat1_1_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_11725, new_AGEMA_signal_11724, new_AGEMA_signal_11723, mcs1_mcs_mat1_1_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .c ({new_AGEMA_signal_13147, new_AGEMA_signal_13146, new_AGEMA_signal_13145, mcs1_mcs_mat1_1_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_14599, new_AGEMA_signal_14598, new_AGEMA_signal_14597, mcs1_mcs_mat1_1_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_11719, new_AGEMA_signal_11718, new_AGEMA_signal_11717, mcs1_mcs_mat1_1_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_15919, new_AGEMA_signal_15918, new_AGEMA_signal_15917, mcs1_mcs_mat1_1_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_13153, new_AGEMA_signal_13152, new_AGEMA_signal_13151, mcs1_mcs_mat1_1_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_11722, new_AGEMA_signal_11721, new_AGEMA_signal_11720, mcs1_mcs_mat1_1_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_14599, new_AGEMA_signal_14598, new_AGEMA_signal_14597, mcs1_mcs_mat1_1_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_10678, new_AGEMA_signal_10677, new_AGEMA_signal_10676, mcs1_mcs_mat1_1_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_11722, new_AGEMA_signal_11721, new_AGEMA_signal_11720, mcs1_mcs_mat1_1_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_11725, new_AGEMA_signal_11724, new_AGEMA_signal_11723, mcs1_mcs_mat1_1_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_9541, new_AGEMA_signal_9540, new_AGEMA_signal_9539, mcs1_mcs_mat1_1_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_13153, new_AGEMA_signal_13152, new_AGEMA_signal_13151, mcs1_mcs_mat1_1_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552]}), .c ({new_AGEMA_signal_11725, new_AGEMA_signal_11724, new_AGEMA_signal_11723, mcs1_mcs_mat1_1_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558]}), .c ({new_AGEMA_signal_9541, new_AGEMA_signal_9540, new_AGEMA_signal_9539, mcs1_mcs_mat1_1_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564]}), .c ({new_AGEMA_signal_10678, new_AGEMA_signal_10677, new_AGEMA_signal_10676, mcs1_mcs_mat1_1_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_11728, new_AGEMA_signal_11727, new_AGEMA_signal_11726, mcs1_mcs_mat1_1_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_13156, new_AGEMA_signal_13155, new_AGEMA_signal_13154, mcs1_mcs_mat1_1_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_10681, new_AGEMA_signal_10680, new_AGEMA_signal_10679, mcs1_mcs_mat1_1_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_9544, new_AGEMA_signal_9543, new_AGEMA_signal_9542, mcs1_mcs_mat1_1_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_11728, new_AGEMA_signal_11727, new_AGEMA_signal_11726, mcs1_mcs_mat1_1_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_13159, new_AGEMA_signal_13158, new_AGEMA_signal_13157, mcs1_mcs_mat1_1_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_14602, new_AGEMA_signal_14601, new_AGEMA_signal_14600, mcs1_mcs_mat1_1_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_11734, new_AGEMA_signal_11733, new_AGEMA_signal_11732, mcs1_mcs_mat1_1_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_9544, new_AGEMA_signal_9543, new_AGEMA_signal_9542, mcs1_mcs_mat1_1_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_13159, new_AGEMA_signal_13158, new_AGEMA_signal_13157, mcs1_mcs_mat1_1_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_14605, new_AGEMA_signal_14604, new_AGEMA_signal_14603, mcs1_mcs_mat1_1_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .c ({new_AGEMA_signal_15922, new_AGEMA_signal_15921, new_AGEMA_signal_15920, mcs1_mcs_mat1_1_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_11734, new_AGEMA_signal_11733, new_AGEMA_signal_11732, mcs1_mcs_mat1_1_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_13162, new_AGEMA_signal_13161, new_AGEMA_signal_13160, mcs1_mcs_mat1_1_mcs_out[24]}), .c ({new_AGEMA_signal_14605, new_AGEMA_signal_14604, new_AGEMA_signal_14603, mcs1_mcs_mat1_1_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_11731, new_AGEMA_signal_11730, new_AGEMA_signal_11729, mcs1_mcs_mat1_1_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .c ({new_AGEMA_signal_13162, new_AGEMA_signal_13161, new_AGEMA_signal_13160, mcs1_mcs_mat1_1_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_10681, new_AGEMA_signal_10680, new_AGEMA_signal_10679, mcs1_mcs_mat1_1_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8749, new_AGEMA_signal_8748, new_AGEMA_signal_8747, mcs1_mcs_mat1_1_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_11731, new_AGEMA_signal_11730, new_AGEMA_signal_11729, mcs1_mcs_mat1_1_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .c ({new_AGEMA_signal_11734, new_AGEMA_signal_11733, new_AGEMA_signal_11732, mcs1_mcs_mat1_1_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576]}), .c ({new_AGEMA_signal_9544, new_AGEMA_signal_9543, new_AGEMA_signal_9542, mcs1_mcs_mat1_1_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582]}), .c ({new_AGEMA_signal_10681, new_AGEMA_signal_10680, new_AGEMA_signal_10679, mcs1_mcs_mat1_1_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_11737, new_AGEMA_signal_11736, new_AGEMA_signal_11735, mcs1_mcs_mat1_1_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .c ({new_AGEMA_signal_13165, new_AGEMA_signal_13164, new_AGEMA_signal_13163, mcs1_mcs_mat1_1_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_10684, new_AGEMA_signal_10683, new_AGEMA_signal_10682, mcs1_mcs_mat1_1_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_9547, new_AGEMA_signal_9546, new_AGEMA_signal_9545, mcs1_mcs_mat1_1_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_11737, new_AGEMA_signal_11736, new_AGEMA_signal_11735, mcs1_mcs_mat1_1_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_13168, new_AGEMA_signal_13167, new_AGEMA_signal_13166, mcs1_mcs_mat1_1_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .c ({new_AGEMA_signal_14608, new_AGEMA_signal_14607, new_AGEMA_signal_14606, mcs1_mcs_mat1_1_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_11743, new_AGEMA_signal_11742, new_AGEMA_signal_11741, mcs1_mcs_mat1_1_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_9547, new_AGEMA_signal_9546, new_AGEMA_signal_9545, mcs1_mcs_mat1_1_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_13168, new_AGEMA_signal_13167, new_AGEMA_signal_13166, mcs1_mcs_mat1_1_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_14611, new_AGEMA_signal_14610, new_AGEMA_signal_14609, mcs1_mcs_mat1_1_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_8410, new_AGEMA_signal_8409, new_AGEMA_signal_8408, mcs1_mcs_mat1_1_mcs_out[86]}), .c ({new_AGEMA_signal_15925, new_AGEMA_signal_15924, new_AGEMA_signal_15923, mcs1_mcs_mat1_1_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_11743, new_AGEMA_signal_11742, new_AGEMA_signal_11741, mcs1_mcs_mat1_1_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_13171, new_AGEMA_signal_13170, new_AGEMA_signal_13169, mcs1_mcs_mat1_1_mcs_out[20]}), .c ({new_AGEMA_signal_14611, new_AGEMA_signal_14610, new_AGEMA_signal_14609, mcs1_mcs_mat1_1_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_11740, new_AGEMA_signal_11739, new_AGEMA_signal_11738, mcs1_mcs_mat1_1_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .c ({new_AGEMA_signal_13171, new_AGEMA_signal_13170, new_AGEMA_signal_13169, mcs1_mcs_mat1_1_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_10684, new_AGEMA_signal_10683, new_AGEMA_signal_10682, mcs1_mcs_mat1_1_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8752, new_AGEMA_signal_8751, new_AGEMA_signal_8750, mcs1_mcs_mat1_1_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_11740, new_AGEMA_signal_11739, new_AGEMA_signal_11738, mcs1_mcs_mat1_1_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588]}), .c ({new_AGEMA_signal_11743, new_AGEMA_signal_11742, new_AGEMA_signal_11741, mcs1_mcs_mat1_1_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594]}), .c ({new_AGEMA_signal_9547, new_AGEMA_signal_9546, new_AGEMA_signal_9545, mcs1_mcs_mat1_1_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({new_AGEMA_signal_10684, new_AGEMA_signal_10683, new_AGEMA_signal_10682, mcs1_mcs_mat1_1_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_17524, new_AGEMA_signal_17523, new_AGEMA_signal_17522, mcs1_mcs_mat1_1_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_17533, new_AGEMA_signal_17532, new_AGEMA_signal_17531, mcs1_mcs_mat1_1_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_18235, new_AGEMA_signal_18234, new_AGEMA_signal_18233, mcs1_mcs_mat1_1_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_18238, new_AGEMA_signal_18237, new_AGEMA_signal_18236, mcs1_mcs_mat1_1_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_13174, new_AGEMA_signal_13173, new_AGEMA_signal_13172, mcs1_mcs_mat1_1_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_18877, new_AGEMA_signal_18876, new_AGEMA_signal_18875, mcs1_mcs_mat1_1_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_18880, new_AGEMA_signal_18879, new_AGEMA_signal_18878, mcs1_mcs_mat1_1_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_14614, new_AGEMA_signal_14613, new_AGEMA_signal_14612, mcs1_mcs_mat1_1_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_19609, new_AGEMA_signal_19608, new_AGEMA_signal_19607, mcs1_mcs_mat1_1_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11400, new_AGEMA_signal_11399, mcs1_mcs_mat1_1_mcs_out[50]}), .b ({new_AGEMA_signal_18238, new_AGEMA_signal_18237, new_AGEMA_signal_18236, mcs1_mcs_mat1_1_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_18880, new_AGEMA_signal_18879, new_AGEMA_signal_18878, mcs1_mcs_mat1_1_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_17527, new_AGEMA_signal_17526, new_AGEMA_signal_17525, mcs1_mcs_mat1_1_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .c ({new_AGEMA_signal_18238, new_AGEMA_signal_18237, new_AGEMA_signal_18236, mcs1_mcs_mat1_1_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_16789, new_AGEMA_signal_16788, new_AGEMA_signal_16787, mcs1_mcs_mat1_1_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_16792, new_AGEMA_signal_16791, new_AGEMA_signal_16790, mcs1_mcs_mat1_1_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_17527, new_AGEMA_signal_17526, new_AGEMA_signal_17525, mcs1_mcs_mat1_1_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_17530, new_AGEMA_signal_17529, new_AGEMA_signal_17528, mcs1_mcs_mat1_1_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_14614, new_AGEMA_signal_14613, new_AGEMA_signal_14612, mcs1_mcs_mat1_1_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_18241, new_AGEMA_signal_18240, new_AGEMA_signal_18239, mcs1_mcs_mat1_1_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606]}), .c ({new_AGEMA_signal_17533, new_AGEMA_signal_17532, new_AGEMA_signal_17531, mcs1_mcs_mat1_1_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612]}), .c ({new_AGEMA_signal_14614, new_AGEMA_signal_14613, new_AGEMA_signal_14612, mcs1_mcs_mat1_1_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618]}), .c ({new_AGEMA_signal_16792, new_AGEMA_signal_16791, new_AGEMA_signal_16790, mcs1_mcs_mat1_1_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_14623, new_AGEMA_signal_14622, new_AGEMA_signal_14621, mcs1_mcs_mat1_1_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, new_AGEMA_signal_10292, mcs1_mcs_mat1_1_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_15928, new_AGEMA_signal_15927, new_AGEMA_signal_15926, mcs1_mcs_mat1_1_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_13183, new_AGEMA_signal_13182, new_AGEMA_signal_13181, mcs1_mcs_mat1_1_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_13177, new_AGEMA_signal_13176, new_AGEMA_signal_13175, mcs1_mcs_mat1_1_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_14617, new_AGEMA_signal_14616, new_AGEMA_signal_14615, mcs1_mcs_mat1_1_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_11749, new_AGEMA_signal_11748, new_AGEMA_signal_11747, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_9550, new_AGEMA_signal_9549, new_AGEMA_signal_9548, mcs1_mcs_mat1_1_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_13177, new_AGEMA_signal_13176, new_AGEMA_signal_13175, mcs1_mcs_mat1_1_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, new_AGEMA_signal_10292, mcs1_mcs_mat1_1_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_13180, new_AGEMA_signal_13179, new_AGEMA_signal_13178, mcs1_mcs_mat1_1_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_14620, new_AGEMA_signal_14619, new_AGEMA_signal_14618, mcs1_mcs_mat1_1_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_11746, new_AGEMA_signal_11745, new_AGEMA_signal_11744, mcs1_mcs_mat1_1_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_11749, new_AGEMA_signal_11748, new_AGEMA_signal_11747, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_13180, new_AGEMA_signal_13179, new_AGEMA_signal_13178, mcs1_mcs_mat1_1_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_8755, new_AGEMA_signal_8754, new_AGEMA_signal_8753, mcs1_mcs_mat1_1_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_9550, new_AGEMA_signal_9549, new_AGEMA_signal_9548, mcs1_mcs_mat1_1_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_10294, new_AGEMA_signal_10293, new_AGEMA_signal_10292, mcs1_mcs_mat1_1_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_15931, new_AGEMA_signal_15930, new_AGEMA_signal_15929, mcs1_mcs_mat1_1_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .c ({new_AGEMA_signal_16795, new_AGEMA_signal_16794, new_AGEMA_signal_16793, mcs1_mcs_mat1_1_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_14623, new_AGEMA_signal_14622, new_AGEMA_signal_14621, mcs1_mcs_mat1_1_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_11749, new_AGEMA_signal_11748, new_AGEMA_signal_11747, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_15931, new_AGEMA_signal_15930, new_AGEMA_signal_15929, mcs1_mcs_mat1_1_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({new_AGEMA_signal_13183, new_AGEMA_signal_13182, new_AGEMA_signal_13181, mcs1_mcs_mat1_1_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_14623, new_AGEMA_signal_14622, new_AGEMA_signal_14621, mcs1_mcs_mat1_1_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({new_AGEMA_signal_11746, new_AGEMA_signal_11745, new_AGEMA_signal_11744, mcs1_mcs_mat1_1_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_13183, new_AGEMA_signal_13182, new_AGEMA_signal_13181, mcs1_mcs_mat1_1_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_8377, new_AGEMA_signal_8376, new_AGEMA_signal_8375, shiftr_out[120]}), .b ({new_AGEMA_signal_10687, new_AGEMA_signal_10686, new_AGEMA_signal_10685, mcs1_mcs_mat1_1_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_11746, new_AGEMA_signal_11745, new_AGEMA_signal_11744, mcs1_mcs_mat1_1_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10416, new_AGEMA_signal_10415, mcs1_mcs_mat1_1_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624]}), .c ({new_AGEMA_signal_11749, new_AGEMA_signal_11748, new_AGEMA_signal_11747, mcs1_mcs_mat1_1_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8580, new_AGEMA_signal_8579, mcs1_mcs_mat1_1_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .c ({new_AGEMA_signal_9550, new_AGEMA_signal_9549, new_AGEMA_signal_9548, mcs1_mcs_mat1_1_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10219, new_AGEMA_signal_10218, new_AGEMA_signal_10217, mcs1_mcs_mat1_1_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636]}), .c ({new_AGEMA_signal_10687, new_AGEMA_signal_10686, new_AGEMA_signal_10685, mcs1_mcs_mat1_1_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_10297, new_AGEMA_signal_10296, new_AGEMA_signal_10295, mcs1_mcs_mat1_1_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .c ({new_AGEMA_signal_10690, new_AGEMA_signal_10689, new_AGEMA_signal_10688, mcs1_mcs_mat1_1_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_13189, new_AGEMA_signal_13188, new_AGEMA_signal_13187, mcs1_mcs_mat1_1_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .c ({new_AGEMA_signal_14626, new_AGEMA_signal_14625, new_AGEMA_signal_14624, mcs1_mcs_mat1_1_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_11752, new_AGEMA_signal_11751, new_AGEMA_signal_11750, mcs1_mcs_mat1_1_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .c ({new_AGEMA_signal_13186, new_AGEMA_signal_13185, new_AGEMA_signal_13184, mcs1_mcs_mat1_1_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_10693, new_AGEMA_signal_10692, new_AGEMA_signal_10691, mcs1_mcs_mat1_1_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_10297, new_AGEMA_signal_10296, new_AGEMA_signal_10295, mcs1_mcs_mat1_1_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_11752, new_AGEMA_signal_11751, new_AGEMA_signal_11750, mcs1_mcs_mat1_1_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_8758, new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_1_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_9553, new_AGEMA_signal_9552, new_AGEMA_signal_9551, mcs1_mcs_mat1_1_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_10297, new_AGEMA_signal_10296, new_AGEMA_signal_10295, mcs1_mcs_mat1_1_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_14629, new_AGEMA_signal_14628, new_AGEMA_signal_14627, mcs1_mcs_mat1_1_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_8392, new_AGEMA_signal_8391, new_AGEMA_signal_8390, shiftr_out[88]}), .c ({new_AGEMA_signal_15934, new_AGEMA_signal_15933, new_AGEMA_signal_15932, mcs1_mcs_mat1_1_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_8758, new_AGEMA_signal_8757, new_AGEMA_signal_8756, mcs1_mcs_mat1_1_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_13189, new_AGEMA_signal_13188, new_AGEMA_signal_13187, mcs1_mcs_mat1_1_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_14629, new_AGEMA_signal_14628, new_AGEMA_signal_14627, mcs1_mcs_mat1_1_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_11755, new_AGEMA_signal_11754, new_AGEMA_signal_11753, mcs1_mcs_mat1_1_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_10693, new_AGEMA_signal_10692, new_AGEMA_signal_10691, mcs1_mcs_mat1_1_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_13189, new_AGEMA_signal_13188, new_AGEMA_signal_13187, mcs1_mcs_mat1_1_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10432, new_AGEMA_signal_10431, new_AGEMA_signal_10430, mcs1_mcs_mat1_1_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642]}), .c ({new_AGEMA_signal_11755, new_AGEMA_signal_11754, new_AGEMA_signal_11753, mcs1_mcs_mat1_1_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8596, new_AGEMA_signal_8595, new_AGEMA_signal_8594, mcs1_mcs_mat1_1_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648]}), .c ({new_AGEMA_signal_9553, new_AGEMA_signal_9552, new_AGEMA_signal_9551, mcs1_mcs_mat1_1_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10234, new_AGEMA_signal_10233, new_AGEMA_signal_10232, shiftr_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654]}), .c ({new_AGEMA_signal_10693, new_AGEMA_signal_10692, new_AGEMA_signal_10691, mcs1_mcs_mat1_1_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_16798, new_AGEMA_signal_16797, new_AGEMA_signal_16796, mcs1_mcs_mat1_1_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_10699, new_AGEMA_signal_10698, new_AGEMA_signal_10697, mcs1_mcs_mat1_1_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_17536, new_AGEMA_signal_17535, new_AGEMA_signal_17534, mcs1_mcs_mat1_1_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_15937, new_AGEMA_signal_15936, new_AGEMA_signal_15935, mcs1_mcs_mat1_1_mcs_out[7]}), .b ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .c ({new_AGEMA_signal_16798, new_AGEMA_signal_16797, new_AGEMA_signal_16796, mcs1_mcs_mat1_1_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_14632, new_AGEMA_signal_14631, new_AGEMA_signal_14630, mcs1_mcs_mat1_1_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .c ({new_AGEMA_signal_15937, new_AGEMA_signal_15936, new_AGEMA_signal_15935, mcs1_mcs_mat1_1_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_13192, new_AGEMA_signal_13191, new_AGEMA_signal_13190, mcs1_mcs_mat1_1_mcs_out[6]}), .b ({new_AGEMA_signal_9559, new_AGEMA_signal_9558, new_AGEMA_signal_9557, mcs1_mcs_mat1_1_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_14632, new_AGEMA_signal_14631, new_AGEMA_signal_14630, mcs1_mcs_mat1_1_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_9556, new_AGEMA_signal_9555, new_AGEMA_signal_9554, mcs1_mcs_mat1_1_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_11758, new_AGEMA_signal_11757, new_AGEMA_signal_11756, mcs1_mcs_mat1_1_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_13192, new_AGEMA_signal_13191, new_AGEMA_signal_13190, mcs1_mcs_mat1_1_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10449, new_AGEMA_signal_10448, shiftr_out[57]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({new_AGEMA_signal_11758, new_AGEMA_signal_11757, new_AGEMA_signal_11756, mcs1_mcs_mat1_1_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8614, new_AGEMA_signal_8613, new_AGEMA_signal_8612, shiftr_out[58]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666]}), .c ({new_AGEMA_signal_9559, new_AGEMA_signal_9558, new_AGEMA_signal_9557, mcs1_mcs_mat1_1_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10252, new_AGEMA_signal_10251, new_AGEMA_signal_10250, mcs1_mcs_mat1_1_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672]}), .c ({new_AGEMA_signal_10699, new_AGEMA_signal_10698, new_AGEMA_signal_10697, mcs1_mcs_mat1_1_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_16801, new_AGEMA_signal_16800, new_AGEMA_signal_16799, mcs1_mcs_mat1_1_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_17539, new_AGEMA_signal_17538, new_AGEMA_signal_17537, mcs1_mcs_mat1_1_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_18247, new_AGEMA_signal_18246, new_AGEMA_signal_18245, mcs1_mcs_mat1_1_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .b ({new_AGEMA_signal_16804, new_AGEMA_signal_16803, new_AGEMA_signal_16802, mcs1_mcs_mat1_1_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_17539, new_AGEMA_signal_17538, new_AGEMA_signal_17537, mcs1_mcs_mat1_1_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_18250, new_AGEMA_signal_18249, new_AGEMA_signal_18248, mcs1_mcs_mat1_1_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_14635, new_AGEMA_signal_14634, new_AGEMA_signal_14633, mcs1_mcs_mat1_1_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_18883, new_AGEMA_signal_18882, new_AGEMA_signal_18881, mcs1_mcs_mat1_1_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_18253, new_AGEMA_signal_18252, new_AGEMA_signal_18251, mcs1_mcs_mat1_1_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_17545, new_AGEMA_signal_17544, new_AGEMA_signal_17543, mcs1_mcs_mat1_1_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_18886, new_AGEMA_signal_18885, new_AGEMA_signal_18884, mcs1_mcs_mat1_1_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_17548, new_AGEMA_signal_17547, new_AGEMA_signal_17546, mcs1_mcs_mat1_1_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_13195, new_AGEMA_signal_13194, new_AGEMA_signal_13193, mcs1_mcs_mat1_1_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_18253, new_AGEMA_signal_18252, new_AGEMA_signal_18251, mcs1_mcs_mat1_1_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16627, new_AGEMA_signal_16626, new_AGEMA_signal_16625, shiftr_out[25]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678]}), .c ({new_AGEMA_signal_17548, new_AGEMA_signal_17547, new_AGEMA_signal_17546, mcs1_mcs_mat1_1_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12840, new_AGEMA_signal_12839, shiftr_out[26]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684]}), .c ({new_AGEMA_signal_14635, new_AGEMA_signal_14634, new_AGEMA_signal_14633, mcs1_mcs_mat1_1_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_1_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15715, new_AGEMA_signal_15714, new_AGEMA_signal_15713, mcs1_mcs_mat1_1_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .c ({new_AGEMA_signal_16804, new_AGEMA_signal_16803, new_AGEMA_signal_16802, mcs1_mcs_mat1_1_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U96 ( .a ({new_AGEMA_signal_20461, new_AGEMA_signal_20460, new_AGEMA_signal_20459, mcs1_mcs_mat1_2_n128}), .b ({new_AGEMA_signal_15940, new_AGEMA_signal_15939, new_AGEMA_signal_15938, mcs1_mcs_mat1_2_n127}), .c ({temp_next_s3[85], temp_next_s2[85], temp_next_s1[85], temp_next_s0[85]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U95 ( .a ({new_AGEMA_signal_14743, new_AGEMA_signal_14742, new_AGEMA_signal_14741, mcs1_mcs_mat1_2_mcs_out[41]}), .b ({new_AGEMA_signal_11854, new_AGEMA_signal_11853, new_AGEMA_signal_11852, mcs1_mcs_mat1_2_mcs_out[45]}), .c ({new_AGEMA_signal_15940, new_AGEMA_signal_15939, new_AGEMA_signal_15938, mcs1_mcs_mat1_2_n127}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U94 ( .a ({new_AGEMA_signal_10303, new_AGEMA_signal_10302, new_AGEMA_signal_10301, mcs1_mcs_mat1_2_mcs_out[33]}), .b ({new_AGEMA_signal_19678, new_AGEMA_signal_19677, new_AGEMA_signal_19676, mcs1_mcs_mat1_2_mcs_out[37]}), .c ({new_AGEMA_signal_20461, new_AGEMA_signal_20460, new_AGEMA_signal_20459, mcs1_mcs_mat1_2_n128}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U93 ( .a ({new_AGEMA_signal_18889, new_AGEMA_signal_18888, new_AGEMA_signal_18887, mcs1_mcs_mat1_2_n126}), .b ({new_AGEMA_signal_17551, new_AGEMA_signal_17550, new_AGEMA_signal_17549, mcs1_mcs_mat1_2_n125}), .c ({temp_next_s3[84], temp_next_s2[84], temp_next_s1[84], temp_next_s0[84]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U92 ( .a ({new_AGEMA_signal_13309, new_AGEMA_signal_13308, new_AGEMA_signal_13307, mcs1_mcs_mat1_2_mcs_out[40]}), .b ({new_AGEMA_signal_16879, new_AGEMA_signal_16878, new_AGEMA_signal_16877, mcs1_mcs_mat1_2_mcs_out[44]}), .c ({new_AGEMA_signal_17551, new_AGEMA_signal_17550, new_AGEMA_signal_17549, mcs1_mcs_mat1_2_n125}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U91 ( .a ({new_AGEMA_signal_16891, new_AGEMA_signal_16890, new_AGEMA_signal_16889, mcs1_mcs_mat1_2_mcs_out[32]}), .b ({new_AGEMA_signal_18304, new_AGEMA_signal_18303, new_AGEMA_signal_18302, mcs1_mcs_mat1_2_mcs_out[36]}), .c ({new_AGEMA_signal_18889, new_AGEMA_signal_18888, new_AGEMA_signal_18887, mcs1_mcs_mat1_2_n126}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U90 ( .a ({new_AGEMA_signal_18892, new_AGEMA_signal_18891, new_AGEMA_signal_18890, mcs1_mcs_mat1_2_n124}), .b ({new_AGEMA_signal_16807, new_AGEMA_signal_16806, new_AGEMA_signal_16805, mcs1_mcs_mat1_2_n123}), .c ({temp_next_s3[55], temp_next_s2[55], temp_next_s1[55], temp_next_s0[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U89 ( .a ({new_AGEMA_signal_13330, new_AGEMA_signal_13329, new_AGEMA_signal_13328, mcs1_mcs_mat1_2_mcs_out[27]}), .b ({new_AGEMA_signal_16030, new_AGEMA_signal_16029, new_AGEMA_signal_16028, mcs1_mcs_mat1_2_mcs_out[31]}), .c ({new_AGEMA_signal_16807, new_AGEMA_signal_16806, new_AGEMA_signal_16805, mcs1_mcs_mat1_2_n123}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U88 ( .a ({new_AGEMA_signal_13342, new_AGEMA_signal_13341, new_AGEMA_signal_13340, mcs1_mcs_mat1_2_mcs_out[19]}), .b ({new_AGEMA_signal_18307, new_AGEMA_signal_18306, new_AGEMA_signal_18305, mcs1_mcs_mat1_2_mcs_out[23]}), .c ({new_AGEMA_signal_18892, new_AGEMA_signal_18891, new_AGEMA_signal_18890, mcs1_mcs_mat1_2_n124}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U87 ( .a ({new_AGEMA_signal_19618, new_AGEMA_signal_19617, new_AGEMA_signal_19616, mcs1_mcs_mat1_2_n122}), .b ({new_AGEMA_signal_15943, new_AGEMA_signal_15942, new_AGEMA_signal_15941, mcs1_mcs_mat1_2_n121}), .c ({temp_next_s3[54], temp_next_s2[54], temp_next_s1[54], temp_next_s0[54]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U86 ( .a ({new_AGEMA_signal_14761, new_AGEMA_signal_14760, new_AGEMA_signal_14759, mcs1_mcs_mat1_2_mcs_out[26]}), .b ({new_AGEMA_signal_14755, new_AGEMA_signal_14754, new_AGEMA_signal_14753, mcs1_mcs_mat1_2_mcs_out[30]}), .c ({new_AGEMA_signal_15943, new_AGEMA_signal_15942, new_AGEMA_signal_15941, mcs1_mcs_mat1_2_n121}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U85 ( .a ({new_AGEMA_signal_14770, new_AGEMA_signal_14769, new_AGEMA_signal_14768, mcs1_mcs_mat1_2_mcs_out[18]}), .b ({new_AGEMA_signal_18955, new_AGEMA_signal_18954, new_AGEMA_signal_18953, mcs1_mcs_mat1_2_mcs_out[22]}), .c ({new_AGEMA_signal_19618, new_AGEMA_signal_19617, new_AGEMA_signal_19616, mcs1_mcs_mat1_2_n122}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U84 ( .a ({new_AGEMA_signal_20467, new_AGEMA_signal_20466, new_AGEMA_signal_20465, mcs1_mcs_mat1_2_n120}), .b ({new_AGEMA_signal_16810, new_AGEMA_signal_16809, new_AGEMA_signal_16808, mcs1_mcs_mat1_2_n119}), .c ({temp_next_s3[53], temp_next_s2[53], temp_next_s1[53], temp_next_s0[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U83 ( .a ({new_AGEMA_signal_16036, new_AGEMA_signal_16035, new_AGEMA_signal_16034, mcs1_mcs_mat1_2_mcs_out[25]}), .b ({new_AGEMA_signal_13324, new_AGEMA_signal_13323, new_AGEMA_signal_13322, mcs1_mcs_mat1_2_mcs_out[29]}), .c ({new_AGEMA_signal_16810, new_AGEMA_signal_16809, new_AGEMA_signal_16808, mcs1_mcs_mat1_2_n119}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U82 ( .a ({new_AGEMA_signal_16039, new_AGEMA_signal_16038, new_AGEMA_signal_16037, mcs1_mcs_mat1_2_mcs_out[17]}), .b ({new_AGEMA_signal_19681, new_AGEMA_signal_19680, new_AGEMA_signal_19679, mcs1_mcs_mat1_2_mcs_out[21]}), .c ({new_AGEMA_signal_20467, new_AGEMA_signal_20466, new_AGEMA_signal_20465, mcs1_mcs_mat1_2_n120}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U81 ( .a ({new_AGEMA_signal_18895, new_AGEMA_signal_18894, new_AGEMA_signal_18893, mcs1_mcs_mat1_2_n118}), .b ({new_AGEMA_signal_16813, new_AGEMA_signal_16812, new_AGEMA_signal_16811, mcs1_mcs_mat1_2_n117}), .c ({temp_next_s3[52], temp_next_s2[52], temp_next_s1[52], temp_next_s0[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U80 ( .a ({new_AGEMA_signal_13336, new_AGEMA_signal_13335, new_AGEMA_signal_13334, mcs1_mcs_mat1_2_mcs_out[24]}), .b ({new_AGEMA_signal_16033, new_AGEMA_signal_16032, new_AGEMA_signal_16031, mcs1_mcs_mat1_2_mcs_out[28]}), .c ({new_AGEMA_signal_16813, new_AGEMA_signal_16812, new_AGEMA_signal_16811, mcs1_mcs_mat1_2_n117}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U79 ( .a ({new_AGEMA_signal_13348, new_AGEMA_signal_13347, new_AGEMA_signal_13346, mcs1_mcs_mat1_2_mcs_out[16]}), .b ({new_AGEMA_signal_18313, new_AGEMA_signal_18312, new_AGEMA_signal_18311, mcs1_mcs_mat1_2_mcs_out[20]}), .c ({new_AGEMA_signal_18895, new_AGEMA_signal_18894, new_AGEMA_signal_18893, mcs1_mcs_mat1_2_n118}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U78 ( .a ({new_AGEMA_signal_16816, new_AGEMA_signal_16815, new_AGEMA_signal_16814, mcs1_mcs_mat1_2_n116}), .b ({new_AGEMA_signal_20470, new_AGEMA_signal_20469, new_AGEMA_signal_20468, mcs1_mcs_mat1_2_n115}), .c ({temp_next_s3[23], temp_next_s2[23], temp_next_s1[23], temp_next_s0[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U77 ( .a ({new_AGEMA_signal_13369, new_AGEMA_signal_13368, new_AGEMA_signal_13367, mcs1_mcs_mat1_2_mcs_out[3]}), .b ({new_AGEMA_signal_19684, new_AGEMA_signal_19683, new_AGEMA_signal_19682, mcs1_mcs_mat1_2_mcs_out[7]}), .c ({new_AGEMA_signal_20470, new_AGEMA_signal_20469, new_AGEMA_signal_20468, mcs1_mcs_mat1_2_n115}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U76 ( .a ({new_AGEMA_signal_10795, new_AGEMA_signal_10794, new_AGEMA_signal_10793, mcs1_mcs_mat1_2_mcs_out[11]}), .b ({new_AGEMA_signal_16042, new_AGEMA_signal_16041, new_AGEMA_signal_16040, mcs1_mcs_mat1_2_mcs_out[15]}), .c ({new_AGEMA_signal_16816, new_AGEMA_signal_16815, new_AGEMA_signal_16814, mcs1_mcs_mat1_2_n116}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U75 ( .a ({new_AGEMA_signal_20473, new_AGEMA_signal_20472, new_AGEMA_signal_20471, mcs1_mcs_mat1_2_n114}), .b ({new_AGEMA_signal_16819, new_AGEMA_signal_16818, new_AGEMA_signal_16817, mcs1_mcs_mat1_2_n113}), .c ({new_AGEMA_signal_21196, new_AGEMA_signal_21195, new_AGEMA_signal_21194, mcs_out[247]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U74 ( .a ({new_AGEMA_signal_15973, new_AGEMA_signal_15972, new_AGEMA_signal_15971, mcs1_mcs_mat1_2_mcs_out[123]}), .b ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_16819, new_AGEMA_signal_16818, new_AGEMA_signal_16817, mcs1_mcs_mat1_2_n113}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U73 ( .a ({new_AGEMA_signal_14662, new_AGEMA_signal_14661, new_AGEMA_signal_14660, mcs1_mcs_mat1_2_mcs_out[115]}), .b ({new_AGEMA_signal_19657, new_AGEMA_signal_19656, new_AGEMA_signal_19655, mcs1_mcs_mat1_2_mcs_out[119]}), .c ({new_AGEMA_signal_20473, new_AGEMA_signal_20472, new_AGEMA_signal_20471, mcs1_mcs_mat1_2_n114}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U72 ( .a ({new_AGEMA_signal_20476, new_AGEMA_signal_20475, new_AGEMA_signal_20474, mcs1_mcs_mat1_2_n112}), .b ({new_AGEMA_signal_13198, new_AGEMA_signal_13197, new_AGEMA_signal_13196, mcs1_mcs_mat1_2_n111}), .c ({new_AGEMA_signal_21199, new_AGEMA_signal_21198, new_AGEMA_signal_21197, mcs_out[246]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U71 ( .a ({new_AGEMA_signal_11761, new_AGEMA_signal_11760, new_AGEMA_signal_11759, mcs1_mcs_mat1_2_mcs_out[122]}), .b ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_13198, new_AGEMA_signal_13197, new_AGEMA_signal_13196, mcs1_mcs_mat1_2_n111}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U70 ( .a ({new_AGEMA_signal_13216, new_AGEMA_signal_13215, new_AGEMA_signal_13214, mcs1_mcs_mat1_2_mcs_out[114]}), .b ({new_AGEMA_signal_19660, new_AGEMA_signal_19659, new_AGEMA_signal_19658, mcs1_mcs_mat1_2_mcs_out[118]}), .c ({new_AGEMA_signal_20476, new_AGEMA_signal_20475, new_AGEMA_signal_20474, mcs1_mcs_mat1_2_n112}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U69 ( .a ({new_AGEMA_signal_15946, new_AGEMA_signal_15945, new_AGEMA_signal_15944, mcs1_mcs_mat1_2_n110}), .b ({new_AGEMA_signal_18898, new_AGEMA_signal_18897, new_AGEMA_signal_18896, mcs1_mcs_mat1_2_n109}), .c ({temp_next_s3[22], temp_next_s2[22], temp_next_s1[22], temp_next_s0[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U68 ( .a ({new_AGEMA_signal_13372, new_AGEMA_signal_13371, new_AGEMA_signal_13370, mcs1_mcs_mat1_2_mcs_out[2]}), .b ({new_AGEMA_signal_18316, new_AGEMA_signal_18315, new_AGEMA_signal_18314, mcs1_mcs_mat1_2_mcs_out[6]}), .c ({new_AGEMA_signal_18898, new_AGEMA_signal_18897, new_AGEMA_signal_18896, mcs1_mcs_mat1_2_n109}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U67 ( .a ({new_AGEMA_signal_14785, new_AGEMA_signal_14784, new_AGEMA_signal_14783, mcs1_mcs_mat1_2_mcs_out[10]}), .b ({new_AGEMA_signal_14776, new_AGEMA_signal_14775, new_AGEMA_signal_14774, mcs1_mcs_mat1_2_mcs_out[14]}), .c ({new_AGEMA_signal_15946, new_AGEMA_signal_15945, new_AGEMA_signal_15944, mcs1_mcs_mat1_2_n110}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U66 ( .a ({new_AGEMA_signal_19627, new_AGEMA_signal_19626, new_AGEMA_signal_19625, mcs1_mcs_mat1_2_n108}), .b ({new_AGEMA_signal_16822, new_AGEMA_signal_16821, new_AGEMA_signal_16820, mcs1_mcs_mat1_2_n107}), .c ({new_AGEMA_signal_20479, new_AGEMA_signal_20478, new_AGEMA_signal_20477, mcs_out[245]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U65 ( .a ({new_AGEMA_signal_15976, new_AGEMA_signal_15975, new_AGEMA_signal_15974, mcs1_mcs_mat1_2_mcs_out[121]}), .b ({new_AGEMA_signal_10702, new_AGEMA_signal_10701, new_AGEMA_signal_10700, mcs1_mcs_mat1_2_mcs_out[125]}), .c ({new_AGEMA_signal_16822, new_AGEMA_signal_16821, new_AGEMA_signal_16820, mcs1_mcs_mat1_2_n107}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U64 ( .a ({new_AGEMA_signal_11767, new_AGEMA_signal_11766, new_AGEMA_signal_11765, mcs1_mcs_mat1_2_mcs_out[113]}), .b ({new_AGEMA_signal_18925, new_AGEMA_signal_18924, new_AGEMA_signal_18923, mcs1_mcs_mat1_2_mcs_out[117]}), .c ({new_AGEMA_signal_19627, new_AGEMA_signal_19626, new_AGEMA_signal_19625, mcs1_mcs_mat1_2_n108}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U63 ( .a ({new_AGEMA_signal_18901, new_AGEMA_signal_18900, new_AGEMA_signal_18899, mcs1_mcs_mat1_2_n106}), .b ({new_AGEMA_signal_15949, new_AGEMA_signal_15948, new_AGEMA_signal_15947, mcs1_mcs_mat1_2_n105}), .c ({new_AGEMA_signal_19630, new_AGEMA_signal_19629, new_AGEMA_signal_19628, mcs_out[244]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U62 ( .a ({new_AGEMA_signal_14656, new_AGEMA_signal_14655, new_AGEMA_signal_14654, mcs1_mcs_mat1_2_mcs_out[120]}), .b ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_15949, new_AGEMA_signal_15948, new_AGEMA_signal_15947, mcs1_mcs_mat1_2_n105}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U61 ( .a ({new_AGEMA_signal_15979, new_AGEMA_signal_15978, new_AGEMA_signal_15977, mcs1_mcs_mat1_2_mcs_out[112]}), .b ({new_AGEMA_signal_18274, new_AGEMA_signal_18273, new_AGEMA_signal_18272, mcs1_mcs_mat1_2_mcs_out[116]}), .c ({new_AGEMA_signal_18901, new_AGEMA_signal_18900, new_AGEMA_signal_18899, mcs1_mcs_mat1_2_n106}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U60 ( .a ({new_AGEMA_signal_19633, new_AGEMA_signal_19632, new_AGEMA_signal_19631, mcs1_mcs_mat1_2_n104}), .b ({new_AGEMA_signal_16825, new_AGEMA_signal_16824, new_AGEMA_signal_16823, mcs1_mcs_mat1_2_n103}), .c ({new_AGEMA_signal_20482, new_AGEMA_signal_20481, new_AGEMA_signal_20480, mcs_out[215]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U59 ( .a ({new_AGEMA_signal_15982, new_AGEMA_signal_15981, new_AGEMA_signal_15980, mcs1_mcs_mat1_2_mcs_out[111]}), .b ({new_AGEMA_signal_15997, new_AGEMA_signal_15996, new_AGEMA_signal_15995, mcs1_mcs_mat1_2_mcs_out[99]}), .c ({new_AGEMA_signal_16825, new_AGEMA_signal_16824, new_AGEMA_signal_16823, mcs1_mcs_mat1_2_n103}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U58 ( .a ({new_AGEMA_signal_18928, new_AGEMA_signal_18927, new_AGEMA_signal_18926, mcs1_mcs_mat1_2_mcs_out[103]}), .b ({new_AGEMA_signal_14674, new_AGEMA_signal_14673, new_AGEMA_signal_14672, mcs1_mcs_mat1_2_mcs_out[107]}), .c ({new_AGEMA_signal_19633, new_AGEMA_signal_19632, new_AGEMA_signal_19631, mcs1_mcs_mat1_2_n104}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U57 ( .a ({new_AGEMA_signal_18256, new_AGEMA_signal_18255, new_AGEMA_signal_18254, mcs1_mcs_mat1_2_n102}), .b ({new_AGEMA_signal_16828, new_AGEMA_signal_16827, new_AGEMA_signal_16826, mcs1_mcs_mat1_2_n101}), .c ({new_AGEMA_signal_18904, new_AGEMA_signal_18903, new_AGEMA_signal_18902, mcs_out[214]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U56 ( .a ({new_AGEMA_signal_15985, new_AGEMA_signal_15984, new_AGEMA_signal_15983, mcs1_mcs_mat1_2_mcs_out[110]}), .b ({new_AGEMA_signal_13240, new_AGEMA_signal_13239, new_AGEMA_signal_13238, mcs1_mcs_mat1_2_mcs_out[98]}), .c ({new_AGEMA_signal_16828, new_AGEMA_signal_16827, new_AGEMA_signal_16826, mcs1_mcs_mat1_2_n101}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U55 ( .a ({new_AGEMA_signal_17572, new_AGEMA_signal_17571, new_AGEMA_signal_17570, mcs1_mcs_mat1_2_mcs_out[102]}), .b ({new_AGEMA_signal_14677, new_AGEMA_signal_14676, new_AGEMA_signal_14675, mcs1_mcs_mat1_2_mcs_out[106]}), .c ({new_AGEMA_signal_18256, new_AGEMA_signal_18255, new_AGEMA_signal_18254, mcs1_mcs_mat1_2_n102}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U54 ( .a ({new_AGEMA_signal_18907, new_AGEMA_signal_18906, new_AGEMA_signal_18905, mcs1_mcs_mat1_2_n100}), .b ({new_AGEMA_signal_16831, new_AGEMA_signal_16830, new_AGEMA_signal_16829, mcs1_mcs_mat1_2_n99}), .c ({new_AGEMA_signal_19636, new_AGEMA_signal_19635, new_AGEMA_signal_19634, mcs_out[213]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U53 ( .a ({new_AGEMA_signal_15988, new_AGEMA_signal_15987, new_AGEMA_signal_15986, mcs1_mcs_mat1_2_mcs_out[109]}), .b ({new_AGEMA_signal_10726, new_AGEMA_signal_10725, new_AGEMA_signal_10724, mcs1_mcs_mat1_2_mcs_out[97]}), .c ({new_AGEMA_signal_16831, new_AGEMA_signal_16830, new_AGEMA_signal_16829, mcs1_mcs_mat1_2_n99}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U52 ( .a ({new_AGEMA_signal_18280, new_AGEMA_signal_18279, new_AGEMA_signal_18278, mcs1_mcs_mat1_2_mcs_out[101]}), .b ({new_AGEMA_signal_14680, new_AGEMA_signal_14679, new_AGEMA_signal_14678, mcs1_mcs_mat1_2_mcs_out[105]}), .c ({new_AGEMA_signal_18907, new_AGEMA_signal_18906, new_AGEMA_signal_18905, mcs1_mcs_mat1_2_n100}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U51 ( .a ({new_AGEMA_signal_19639, new_AGEMA_signal_19638, new_AGEMA_signal_19637, mcs1_mcs_mat1_2_n98}), .b ({new_AGEMA_signal_18259, new_AGEMA_signal_18258, new_AGEMA_signal_18257, mcs1_mcs_mat1_2_n97}), .c ({new_AGEMA_signal_20485, new_AGEMA_signal_20484, new_AGEMA_signal_20483, mcs_out[212]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U50 ( .a ({new_AGEMA_signal_15991, new_AGEMA_signal_15990, new_AGEMA_signal_15989, mcs1_mcs_mat1_2_mcs_out[108]}), .b ({new_AGEMA_signal_17584, new_AGEMA_signal_17583, new_AGEMA_signal_17582, mcs1_mcs_mat1_2_mcs_out[96]}), .c ({new_AGEMA_signal_18259, new_AGEMA_signal_18258, new_AGEMA_signal_18257, mcs1_mcs_mat1_2_n97}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U49 ( .a ({new_AGEMA_signal_18931, new_AGEMA_signal_18930, new_AGEMA_signal_18929, mcs1_mcs_mat1_2_mcs_out[100]}), .b ({new_AGEMA_signal_15994, new_AGEMA_signal_15993, new_AGEMA_signal_15992, mcs1_mcs_mat1_2_mcs_out[104]}), .c ({new_AGEMA_signal_19639, new_AGEMA_signal_19638, new_AGEMA_signal_19637, mcs1_mcs_mat1_2_n98}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U48 ( .a ({new_AGEMA_signal_18262, new_AGEMA_signal_18261, new_AGEMA_signal_18260, mcs1_mcs_mat1_2_n96}), .b ({new_AGEMA_signal_15952, new_AGEMA_signal_15951, new_AGEMA_signal_15950, mcs1_mcs_mat1_2_n95}), .c ({new_AGEMA_signal_18910, new_AGEMA_signal_18909, new_AGEMA_signal_18908, mcs_out[183]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U47 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_14692, new_AGEMA_signal_14691, new_AGEMA_signal_14690, mcs1_mcs_mat1_2_mcs_out[95]}), .c ({new_AGEMA_signal_15952, new_AGEMA_signal_15951, new_AGEMA_signal_15950, mcs1_mcs_mat1_2_n95}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U46 ( .a ({new_AGEMA_signal_13246, new_AGEMA_signal_13245, new_AGEMA_signal_13244, mcs1_mcs_mat1_2_mcs_out[83]}), .b ({new_AGEMA_signal_17587, new_AGEMA_signal_17586, new_AGEMA_signal_17585, mcs1_mcs_mat1_2_mcs_out[87]}), .c ({new_AGEMA_signal_18262, new_AGEMA_signal_18261, new_AGEMA_signal_18260, mcs1_mcs_mat1_2_n96}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U45 ( .a ({new_AGEMA_signal_14638, new_AGEMA_signal_14637, new_AGEMA_signal_14636, mcs1_mcs_mat1_2_n94}), .b ({new_AGEMA_signal_13201, new_AGEMA_signal_13200, new_AGEMA_signal_13199, mcs1_mcs_mat1_2_n93}), .c ({new_AGEMA_signal_15955, new_AGEMA_signal_15954, new_AGEMA_signal_15953, mcs_out[182]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U43 ( .a ({new_AGEMA_signal_13249, new_AGEMA_signal_13248, new_AGEMA_signal_13247, mcs1_mcs_mat1_2_mcs_out[82]}), .b ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_14638, new_AGEMA_signal_14637, new_AGEMA_signal_14636, mcs1_mcs_mat1_2_n94}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U42 ( .a ({new_AGEMA_signal_16834, new_AGEMA_signal_16833, new_AGEMA_signal_16832, mcs1_mcs_mat1_2_n92}), .b ({new_AGEMA_signal_13204, new_AGEMA_signal_13203, new_AGEMA_signal_13202, mcs1_mcs_mat1_2_n91}), .c ({new_AGEMA_signal_17554, new_AGEMA_signal_17553, new_AGEMA_signal_17552, mcs_out[181]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U41 ( .a ({new_AGEMA_signal_10744, new_AGEMA_signal_10743, new_AGEMA_signal_10742, mcs1_mcs_mat1_2_mcs_out[89]}), .b ({new_AGEMA_signal_11794, new_AGEMA_signal_11793, new_AGEMA_signal_11792, mcs1_mcs_mat1_2_mcs_out[93]}), .c ({new_AGEMA_signal_13204, new_AGEMA_signal_13203, new_AGEMA_signal_13202, mcs1_mcs_mat1_2_n91}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U40 ( .a ({new_AGEMA_signal_13252, new_AGEMA_signal_13251, new_AGEMA_signal_13250, mcs1_mcs_mat1_2_mcs_out[81]}), .b ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_16834, new_AGEMA_signal_16833, new_AGEMA_signal_16832, mcs1_mcs_mat1_2_n92}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U39 ( .a ({new_AGEMA_signal_18913, new_AGEMA_signal_18912, new_AGEMA_signal_18911, mcs1_mcs_mat1_2_n90}), .b ({new_AGEMA_signal_16837, new_AGEMA_signal_16836, new_AGEMA_signal_16835, mcs1_mcs_mat1_2_n89}), .c ({new_AGEMA_signal_19642, new_AGEMA_signal_19641, new_AGEMA_signal_19640, mcs_out[180]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U38 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_16000, new_AGEMA_signal_15999, new_AGEMA_signal_15998, mcs1_mcs_mat1_2_mcs_out[92]}), .c ({new_AGEMA_signal_16837, new_AGEMA_signal_16836, new_AGEMA_signal_16835, mcs1_mcs_mat1_2_n89}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U37 ( .a ({new_AGEMA_signal_14698, new_AGEMA_signal_14697, new_AGEMA_signal_14696, mcs1_mcs_mat1_2_mcs_out[80]}), .b ({new_AGEMA_signal_18286, new_AGEMA_signal_18285, new_AGEMA_signal_18284, mcs1_mcs_mat1_2_mcs_out[84]}), .c ({new_AGEMA_signal_18913, new_AGEMA_signal_18912, new_AGEMA_signal_18911, mcs1_mcs_mat1_2_n90}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U36 ( .a ({new_AGEMA_signal_15958, new_AGEMA_signal_15957, new_AGEMA_signal_15956, mcs1_mcs_mat1_2_n88}), .b ({new_AGEMA_signal_17557, new_AGEMA_signal_17556, new_AGEMA_signal_17555, mcs1_mcs_mat1_2_n87}), .c ({temp_next_s3[21], temp_next_s2[21], temp_next_s1[21], temp_next_s0[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U35 ( .a ({new_AGEMA_signal_16900, new_AGEMA_signal_16899, new_AGEMA_signal_16898, mcs1_mcs_mat1_2_mcs_out[5]}), .b ({new_AGEMA_signal_13360, new_AGEMA_signal_13359, new_AGEMA_signal_13358, mcs1_mcs_mat1_2_mcs_out[9]}), .c ({new_AGEMA_signal_17557, new_AGEMA_signal_17556, new_AGEMA_signal_17555, mcs1_mcs_mat1_2_n87}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U34 ( .a ({new_AGEMA_signal_14779, new_AGEMA_signal_14778, new_AGEMA_signal_14777, mcs1_mcs_mat1_2_mcs_out[13]}), .b ({new_AGEMA_signal_14797, new_AGEMA_signal_14796, new_AGEMA_signal_14795, mcs1_mcs_mat1_2_mcs_out[1]}), .c ({new_AGEMA_signal_15958, new_AGEMA_signal_15957, new_AGEMA_signal_15956, mcs1_mcs_mat1_2_n88}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U33 ( .a ({new_AGEMA_signal_19645, new_AGEMA_signal_19644, new_AGEMA_signal_19643, mcs1_mcs_mat1_2_n86}), .b ({new_AGEMA_signal_15961, new_AGEMA_signal_15960, new_AGEMA_signal_15959, mcs1_mcs_mat1_2_n85}), .c ({new_AGEMA_signal_20488, new_AGEMA_signal_20487, new_AGEMA_signal_20486, mcs_out[151]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U32 ( .a ({new_AGEMA_signal_11818, new_AGEMA_signal_11817, new_AGEMA_signal_11816, mcs1_mcs_mat1_2_mcs_out[75]}), .b ({new_AGEMA_signal_14701, new_AGEMA_signal_14700, new_AGEMA_signal_14699, mcs1_mcs_mat1_2_mcs_out[79]}), .c ({new_AGEMA_signal_15961, new_AGEMA_signal_15960, new_AGEMA_signal_15959, mcs1_mcs_mat1_2_n85}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U31 ( .a ({new_AGEMA_signal_16012, new_AGEMA_signal_16011, new_AGEMA_signal_16010, mcs1_mcs_mat1_2_mcs_out[67]}), .b ({new_AGEMA_signal_18934, new_AGEMA_signal_18933, new_AGEMA_signal_18932, mcs1_mcs_mat1_2_mcs_out[71]}), .c ({new_AGEMA_signal_19645, new_AGEMA_signal_19644, new_AGEMA_signal_19643, mcs1_mcs_mat1_2_n86}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U30 ( .a ({new_AGEMA_signal_20491, new_AGEMA_signal_20490, new_AGEMA_signal_20489, mcs1_mcs_mat1_2_n84}), .b ({new_AGEMA_signal_16840, new_AGEMA_signal_16839, new_AGEMA_signal_16838, mcs1_mcs_mat1_2_n83}), .c ({new_AGEMA_signal_21202, new_AGEMA_signal_21201, new_AGEMA_signal_21200, mcs_out[150]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U29 ( .a ({new_AGEMA_signal_16006, new_AGEMA_signal_16005, new_AGEMA_signal_16004, mcs1_mcs_mat1_2_mcs_out[74]}), .b ({new_AGEMA_signal_9592, new_AGEMA_signal_9591, new_AGEMA_signal_9590, mcs1_mcs_mat1_2_mcs_out[78]}), .c ({new_AGEMA_signal_16840, new_AGEMA_signal_16839, new_AGEMA_signal_16838, mcs1_mcs_mat1_2_n83}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U28 ( .a ({new_AGEMA_signal_14716, new_AGEMA_signal_14715, new_AGEMA_signal_14714, mcs1_mcs_mat1_2_mcs_out[66]}), .b ({new_AGEMA_signal_19663, new_AGEMA_signal_19662, new_AGEMA_signal_19661, mcs1_mcs_mat1_2_mcs_out[70]}), .c ({new_AGEMA_signal_20491, new_AGEMA_signal_20490, new_AGEMA_signal_20489, mcs1_mcs_mat1_2_n84}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U27 ( .a ({new_AGEMA_signal_20494, new_AGEMA_signal_20493, new_AGEMA_signal_20492, mcs1_mcs_mat1_2_n82}), .b ({new_AGEMA_signal_14641, new_AGEMA_signal_14640, new_AGEMA_signal_14639, mcs1_mcs_mat1_2_n81}), .c ({new_AGEMA_signal_21205, new_AGEMA_signal_21204, new_AGEMA_signal_21203, mcs_out[149]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U26 ( .a ({new_AGEMA_signal_13261, new_AGEMA_signal_13260, new_AGEMA_signal_13259, mcs1_mcs_mat1_2_mcs_out[73]}), .b ({new_AGEMA_signal_11812, new_AGEMA_signal_11811, new_AGEMA_signal_11810, mcs1_mcs_mat1_2_mcs_out[77]}), .c ({new_AGEMA_signal_14641, new_AGEMA_signal_14640, new_AGEMA_signal_14639, mcs1_mcs_mat1_2_n81}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U25 ( .a ({new_AGEMA_signal_11827, new_AGEMA_signal_11826, new_AGEMA_signal_11825, mcs1_mcs_mat1_2_mcs_out[65]}), .b ({new_AGEMA_signal_19666, new_AGEMA_signal_19665, new_AGEMA_signal_19664, mcs1_mcs_mat1_2_mcs_out[69]}), .c ({new_AGEMA_signal_20494, new_AGEMA_signal_20493, new_AGEMA_signal_20492, mcs1_mcs_mat1_2_n82}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U24 ( .a ({new_AGEMA_signal_19648, new_AGEMA_signal_19647, new_AGEMA_signal_19646, mcs1_mcs_mat1_2_n80}), .b ({new_AGEMA_signal_16843, new_AGEMA_signal_16842, new_AGEMA_signal_16841, mcs1_mcs_mat1_2_n79}), .c ({new_AGEMA_signal_20497, new_AGEMA_signal_20496, new_AGEMA_signal_20495, mcs_out[148]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U23 ( .a ({new_AGEMA_signal_16009, new_AGEMA_signal_16008, new_AGEMA_signal_16007, mcs1_mcs_mat1_2_mcs_out[72]}), .b ({new_AGEMA_signal_16003, new_AGEMA_signal_16002, new_AGEMA_signal_16001, mcs1_mcs_mat1_2_mcs_out[76]}), .c ({new_AGEMA_signal_16843, new_AGEMA_signal_16842, new_AGEMA_signal_16841, mcs1_mcs_mat1_2_n79}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U22 ( .a ({new_AGEMA_signal_16873, new_AGEMA_signal_16872, new_AGEMA_signal_16871, mcs1_mcs_mat1_2_mcs_out[64]}), .b ({new_AGEMA_signal_18940, new_AGEMA_signal_18939, new_AGEMA_signal_18938, mcs1_mcs_mat1_2_mcs_out[68]}), .c ({new_AGEMA_signal_19648, new_AGEMA_signal_19647, new_AGEMA_signal_19646, mcs1_mcs_mat1_2_n80}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U21 ( .a ({new_AGEMA_signal_19651, new_AGEMA_signal_19650, new_AGEMA_signal_19649, mcs1_mcs_mat1_2_n78}), .b ({new_AGEMA_signal_15964, new_AGEMA_signal_15963, new_AGEMA_signal_15962, mcs1_mcs_mat1_2_n77}), .c ({temp_next_s3[119], temp_next_s2[119], temp_next_s1[119], temp_next_s0[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U20 ( .a ({new_AGEMA_signal_13282, new_AGEMA_signal_13281, new_AGEMA_signal_13280, mcs1_mcs_mat1_2_mcs_out[59]}), .b ({new_AGEMA_signal_14722, new_AGEMA_signal_14721, new_AGEMA_signal_14720, mcs1_mcs_mat1_2_mcs_out[63]}), .c ({new_AGEMA_signal_15964, new_AGEMA_signal_15963, new_AGEMA_signal_15962, mcs1_mcs_mat1_2_n77}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U19 ( .a ({new_AGEMA_signal_11851, new_AGEMA_signal_11850, new_AGEMA_signal_11849, mcs1_mcs_mat1_2_mcs_out[51]}), .b ({new_AGEMA_signal_18943, new_AGEMA_signal_18942, new_AGEMA_signal_18941, mcs1_mcs_mat1_2_mcs_out[55]}), .c ({new_AGEMA_signal_19651, new_AGEMA_signal_19650, new_AGEMA_signal_19649, mcs1_mcs_mat1_2_n78}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U18 ( .a ({new_AGEMA_signal_20503, new_AGEMA_signal_20502, new_AGEMA_signal_20501, mcs1_mcs_mat1_2_n76}), .b ({new_AGEMA_signal_14644, new_AGEMA_signal_14643, new_AGEMA_signal_14642, mcs1_mcs_mat1_2_n75}), .c ({temp_next_s3[118], temp_next_s2[118], temp_next_s1[118], temp_next_s0[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U17 ( .a ({new_AGEMA_signal_11839, new_AGEMA_signal_11838, new_AGEMA_signal_11837, mcs1_mcs_mat1_2_mcs_out[58]}), .b ({new_AGEMA_signal_13273, new_AGEMA_signal_13272, new_AGEMA_signal_13271, mcs1_mcs_mat1_2_mcs_out[62]}), .c ({new_AGEMA_signal_14644, new_AGEMA_signal_14643, new_AGEMA_signal_14642, mcs1_mcs_mat1_2_n75}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U16 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_19669, new_AGEMA_signal_19668, new_AGEMA_signal_19667, mcs1_mcs_mat1_2_mcs_out[54]}), .c ({new_AGEMA_signal_20503, new_AGEMA_signal_20502, new_AGEMA_signal_20501, mcs1_mcs_mat1_2_n76}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U15 ( .a ({new_AGEMA_signal_20506, new_AGEMA_signal_20505, new_AGEMA_signal_20504, mcs1_mcs_mat1_2_n74}), .b ({new_AGEMA_signal_14647, new_AGEMA_signal_14646, new_AGEMA_signal_14645, mcs1_mcs_mat1_2_n73}), .c ({temp_next_s3[117], temp_next_s2[117], temp_next_s1[117], temp_next_s0[117]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U14 ( .a ({new_AGEMA_signal_13285, new_AGEMA_signal_13284, new_AGEMA_signal_13283, mcs1_mcs_mat1_2_mcs_out[57]}), .b ({new_AGEMA_signal_13276, new_AGEMA_signal_13275, new_AGEMA_signal_13274, mcs1_mcs_mat1_2_mcs_out[61]}), .c ({new_AGEMA_signal_14647, new_AGEMA_signal_14646, new_AGEMA_signal_14645, mcs1_mcs_mat1_2_n73}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U13 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({new_AGEMA_signal_19672, new_AGEMA_signal_19671, new_AGEMA_signal_19670, mcs1_mcs_mat1_2_mcs_out[53]}), .c ({new_AGEMA_signal_20506, new_AGEMA_signal_20505, new_AGEMA_signal_20504, mcs1_mcs_mat1_2_n74}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U12 ( .a ({new_AGEMA_signal_19654, new_AGEMA_signal_19653, new_AGEMA_signal_19652, mcs1_mcs_mat1_2_n72}), .b ({new_AGEMA_signal_16846, new_AGEMA_signal_16845, new_AGEMA_signal_16844, mcs1_mcs_mat1_2_n71}), .c ({temp_next_s3[116], temp_next_s2[116], temp_next_s1[116], temp_next_s0[116]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U11 ( .a ({new_AGEMA_signal_14728, new_AGEMA_signal_14727, new_AGEMA_signal_14726, mcs1_mcs_mat1_2_mcs_out[56]}), .b ({new_AGEMA_signal_16018, new_AGEMA_signal_16017, new_AGEMA_signal_16016, mcs1_mcs_mat1_2_mcs_out[60]}), .c ({new_AGEMA_signal_16846, new_AGEMA_signal_16845, new_AGEMA_signal_16844, mcs1_mcs_mat1_2_n71}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U10 ( .a ({new_AGEMA_signal_13294, new_AGEMA_signal_13293, new_AGEMA_signal_13292, mcs1_mcs_mat1_2_mcs_out[48]}), .b ({new_AGEMA_signal_18949, new_AGEMA_signal_18948, new_AGEMA_signal_18947, mcs1_mcs_mat1_2_mcs_out[52]}), .c ({new_AGEMA_signal_19654, new_AGEMA_signal_19653, new_AGEMA_signal_19652, mcs1_mcs_mat1_2_n72}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U9 ( .a ({new_AGEMA_signal_20512, new_AGEMA_signal_20511, new_AGEMA_signal_20510, mcs1_mcs_mat1_2_n70}), .b ({new_AGEMA_signal_15967, new_AGEMA_signal_15966, new_AGEMA_signal_15965, mcs1_mcs_mat1_2_n69}), .c ({temp_next_s3[87], temp_next_s2[87], temp_next_s1[87], temp_next_s0[87]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U8 ( .a ({new_AGEMA_signal_14737, new_AGEMA_signal_14736, new_AGEMA_signal_14735, mcs1_mcs_mat1_2_mcs_out[43]}), .b ({new_AGEMA_signal_14734, new_AGEMA_signal_14733, new_AGEMA_signal_14732, mcs1_mcs_mat1_2_mcs_out[47]}), .c ({new_AGEMA_signal_15967, new_AGEMA_signal_15966, new_AGEMA_signal_15965, mcs1_mcs_mat1_2_n69}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U7 ( .a ({new_AGEMA_signal_14749, new_AGEMA_signal_14748, new_AGEMA_signal_14747, mcs1_mcs_mat1_2_mcs_out[35]}), .b ({new_AGEMA_signal_19675, new_AGEMA_signal_19674, new_AGEMA_signal_19673, mcs1_mcs_mat1_2_mcs_out[39]}), .c ({new_AGEMA_signal_20512, new_AGEMA_signal_20511, new_AGEMA_signal_20510, mcs1_mcs_mat1_2_n70}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U6 ( .a ({new_AGEMA_signal_18268, new_AGEMA_signal_18267, new_AGEMA_signal_18266, mcs1_mcs_mat1_2_n68}), .b ({new_AGEMA_signal_15970, new_AGEMA_signal_15969, new_AGEMA_signal_15968, mcs1_mcs_mat1_2_n67}), .c ({temp_next_s3[86], temp_next_s2[86], temp_next_s1[86], temp_next_s0[86]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U5 ( .a ({new_AGEMA_signal_14740, new_AGEMA_signal_14739, new_AGEMA_signal_14738, mcs1_mcs_mat1_2_mcs_out[42]}), .b ({new_AGEMA_signal_10765, new_AGEMA_signal_10764, new_AGEMA_signal_10763, mcs1_mcs_mat1_2_mcs_out[46]}), .c ({new_AGEMA_signal_15970, new_AGEMA_signal_15969, new_AGEMA_signal_15968, mcs1_mcs_mat1_2_n67}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U4 ( .a ({new_AGEMA_signal_13315, new_AGEMA_signal_13314, new_AGEMA_signal_13313, mcs1_mcs_mat1_2_mcs_out[34]}), .b ({new_AGEMA_signal_17611, new_AGEMA_signal_17610, new_AGEMA_signal_17609, mcs1_mcs_mat1_2_mcs_out[38]}), .c ({new_AGEMA_signal_18268, new_AGEMA_signal_18267, new_AGEMA_signal_18266, mcs1_mcs_mat1_2_n68}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U3 ( .a ({new_AGEMA_signal_17560, new_AGEMA_signal_17559, new_AGEMA_signal_17558, mcs1_mcs_mat1_2_n66}), .b ({new_AGEMA_signal_21685, new_AGEMA_signal_21684, new_AGEMA_signal_21683, mcs1_mcs_mat1_2_n65}), .c ({temp_next_s3[20], temp_next_s2[20], temp_next_s1[20], temp_next_s0[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U2 ( .a ({new_AGEMA_signal_21217, new_AGEMA_signal_21216, new_AGEMA_signal_21215, mcs1_mcs_mat1_2_mcs_out[4]}), .b ({new_AGEMA_signal_16048, new_AGEMA_signal_16047, new_AGEMA_signal_16046, mcs1_mcs_mat1_2_mcs_out[8]}), .c ({new_AGEMA_signal_21685, new_AGEMA_signal_21684, new_AGEMA_signal_21683, mcs1_mcs_mat1_2_n65}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_U1 ( .a ({new_AGEMA_signal_14800, new_AGEMA_signal_14799, new_AGEMA_signal_14798, mcs1_mcs_mat1_2_mcs_out[0]}), .b ({new_AGEMA_signal_16897, new_AGEMA_signal_16896, new_AGEMA_signal_16895, mcs1_mcs_mat1_2_mcs_out[12]}), .c ({new_AGEMA_signal_17560, new_AGEMA_signal_17559, new_AGEMA_signal_17558, mcs1_mcs_mat1_2_n66}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_14650, new_AGEMA_signal_14649, new_AGEMA_signal_14648, mcs1_mcs_mat1_2_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_15973, new_AGEMA_signal_15972, new_AGEMA_signal_15971, mcs1_mcs_mat1_2_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_13207, new_AGEMA_signal_13206, new_AGEMA_signal_13205, mcs1_mcs_mat1_2_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_8764, new_AGEMA_signal_8763, new_AGEMA_signal_8762, mcs1_mcs_mat1_2_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_14650, new_AGEMA_signal_14649, new_AGEMA_signal_14648, mcs1_mcs_mat1_2_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_9562, new_AGEMA_signal_9561, new_AGEMA_signal_9560, mcs1_mcs_mat1_2_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_10705, new_AGEMA_signal_10704, new_AGEMA_signal_10703, mcs1_mcs_mat1_2_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_11761, new_AGEMA_signal_11760, new_AGEMA_signal_11759, mcs1_mcs_mat1_2_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_9565, new_AGEMA_signal_9564, new_AGEMA_signal_9563, mcs1_mcs_mat1_2_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .c ({new_AGEMA_signal_10705, new_AGEMA_signal_10704, new_AGEMA_signal_10703, mcs1_mcs_mat1_2_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_14653, new_AGEMA_signal_14652, new_AGEMA_signal_14651, mcs1_mcs_mat1_2_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .c ({new_AGEMA_signal_15976, new_AGEMA_signal_15975, new_AGEMA_signal_15974, mcs1_mcs_mat1_2_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_13207, new_AGEMA_signal_13206, new_AGEMA_signal_13205, mcs1_mcs_mat1_2_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_14653, new_AGEMA_signal_14652, new_AGEMA_signal_14651, mcs1_mcs_mat1_2_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_11764, new_AGEMA_signal_11763, new_AGEMA_signal_11762, mcs1_mcs_mat1_2_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_10708, new_AGEMA_signal_10707, new_AGEMA_signal_10706, mcs1_mcs_mat1_2_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_13207, new_AGEMA_signal_13206, new_AGEMA_signal_13205, mcs1_mcs_mat1_2_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_13210, new_AGEMA_signal_13209, new_AGEMA_signal_13208, mcs1_mcs_mat1_2_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_14656, new_AGEMA_signal_14655, new_AGEMA_signal_14654, mcs1_mcs_mat1_2_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_11764, new_AGEMA_signal_11763, new_AGEMA_signal_11762, mcs1_mcs_mat1_2_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9565, new_AGEMA_signal_9564, new_AGEMA_signal_9563, mcs1_mcs_mat1_2_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_13210, new_AGEMA_signal_13209, new_AGEMA_signal_13208, mcs1_mcs_mat1_2_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696]}), .c ({new_AGEMA_signal_11764, new_AGEMA_signal_11763, new_AGEMA_signal_11762, mcs1_mcs_mat1_2_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702]}), .c ({new_AGEMA_signal_9565, new_AGEMA_signal_9564, new_AGEMA_signal_9563, mcs1_mcs_mat1_2_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708]}), .c ({new_AGEMA_signal_10708, new_AGEMA_signal_10707, new_AGEMA_signal_10706, mcs1_mcs_mat1_2_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_18919, new_AGEMA_signal_18918, new_AGEMA_signal_18917, mcs1_mcs_mat1_2_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .c ({new_AGEMA_signal_19657, new_AGEMA_signal_19656, new_AGEMA_signal_19655, mcs1_mcs_mat1_2_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_18271, new_AGEMA_signal_18270, new_AGEMA_signal_18269, mcs1_mcs_mat1_2_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_16855, new_AGEMA_signal_16854, new_AGEMA_signal_16853, mcs1_mcs_mat1_2_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_18919, new_AGEMA_signal_18918, new_AGEMA_signal_18917, mcs1_mcs_mat1_2_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_18922, new_AGEMA_signal_18921, new_AGEMA_signal_18920, mcs1_mcs_mat1_2_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_17566, new_AGEMA_signal_17565, new_AGEMA_signal_17564, mcs1_mcs_mat1_2_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_19660, new_AGEMA_signal_19659, new_AGEMA_signal_19658, mcs1_mcs_mat1_2_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_18271, new_AGEMA_signal_18270, new_AGEMA_signal_18269, mcs1_mcs_mat1_2_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .c ({new_AGEMA_signal_18922, new_AGEMA_signal_18921, new_AGEMA_signal_18920, mcs1_mcs_mat1_2_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_18271, new_AGEMA_signal_18270, new_AGEMA_signal_18269, mcs1_mcs_mat1_2_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_17563, new_AGEMA_signal_17562, new_AGEMA_signal_17561, mcs1_mcs_mat1_2_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_18925, new_AGEMA_signal_18924, new_AGEMA_signal_18923, mcs1_mcs_mat1_2_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_17569, new_AGEMA_signal_17568, new_AGEMA_signal_17567, mcs1_mcs_mat1_2_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_14659, new_AGEMA_signal_14658, new_AGEMA_signal_14657, mcs1_mcs_mat1_2_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_18271, new_AGEMA_signal_18270, new_AGEMA_signal_18269, mcs1_mcs_mat1_2_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_16852, new_AGEMA_signal_16851, new_AGEMA_signal_16850, mcs1_mcs_mat1_2_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_17566, new_AGEMA_signal_17565, new_AGEMA_signal_17564, mcs1_mcs_mat1_2_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_18274, new_AGEMA_signal_18273, new_AGEMA_signal_18272, mcs1_mcs_mat1_2_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_13213, new_AGEMA_signal_13212, new_AGEMA_signal_13211, mcs1_mcs_mat1_2_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_16855, new_AGEMA_signal_16854, new_AGEMA_signal_16853, mcs1_mcs_mat1_2_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_17566, new_AGEMA_signal_17565, new_AGEMA_signal_17564, mcs1_mcs_mat1_2_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_14659, new_AGEMA_signal_14658, new_AGEMA_signal_14657, mcs1_mcs_mat1_2_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_16852, new_AGEMA_signal_16851, new_AGEMA_signal_16850, mcs1_mcs_mat1_2_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714]}), .c ({new_AGEMA_signal_17569, new_AGEMA_signal_17568, new_AGEMA_signal_17567, mcs1_mcs_mat1_2_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({new_AGEMA_signal_14659, new_AGEMA_signal_14658, new_AGEMA_signal_14657, mcs1_mcs_mat1_2_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726]}), .c ({new_AGEMA_signal_16855, new_AGEMA_signal_16854, new_AGEMA_signal_16853, mcs1_mcs_mat1_2_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_13219, new_AGEMA_signal_13218, new_AGEMA_signal_13217, mcs1_mcs_mat1_2_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_9568, new_AGEMA_signal_9567, new_AGEMA_signal_9566, mcs1_mcs_mat1_2_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_14662, new_AGEMA_signal_14661, new_AGEMA_signal_14660, mcs1_mcs_mat1_2_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_10711, new_AGEMA_signal_10710, new_AGEMA_signal_10709, mcs1_mcs_mat1_2_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_10714, new_AGEMA_signal_10713, new_AGEMA_signal_10712, mcs1_mcs_mat1_2_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_11767, new_AGEMA_signal_11766, new_AGEMA_signal_11765, mcs1_mcs_mat1_2_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_13222, new_AGEMA_signal_13221, new_AGEMA_signal_13220, mcs1_mcs_mat1_2_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_14665, new_AGEMA_signal_14664, new_AGEMA_signal_14663, mcs1_mcs_mat1_2_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_15979, new_AGEMA_signal_15978, new_AGEMA_signal_15977, mcs1_mcs_mat1_2_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_13219, new_AGEMA_signal_13218, new_AGEMA_signal_13217, mcs1_mcs_mat1_2_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_14665, new_AGEMA_signal_14664, new_AGEMA_signal_14663, mcs1_mcs_mat1_2_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_8767, new_AGEMA_signal_8766, new_AGEMA_signal_8765, mcs1_mcs_mat1_2_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_11773, new_AGEMA_signal_11772, new_AGEMA_signal_11771, mcs1_mcs_mat1_2_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_13219, new_AGEMA_signal_13218, new_AGEMA_signal_13217, mcs1_mcs_mat1_2_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_9571, new_AGEMA_signal_9570, new_AGEMA_signal_9569, mcs1_mcs_mat1_2_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_11770, new_AGEMA_signal_11769, new_AGEMA_signal_11768, mcs1_mcs_mat1_2_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_13222, new_AGEMA_signal_13221, new_AGEMA_signal_13220, mcs1_mcs_mat1_2_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732]}), .c ({new_AGEMA_signal_11773, new_AGEMA_signal_11772, new_AGEMA_signal_11771, mcs1_mcs_mat1_2_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738]}), .c ({new_AGEMA_signal_9571, new_AGEMA_signal_9570, new_AGEMA_signal_9569, mcs1_mcs_mat1_2_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744]}), .c ({new_AGEMA_signal_10714, new_AGEMA_signal_10713, new_AGEMA_signal_10712, mcs1_mcs_mat1_2_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({new_AGEMA_signal_14668, new_AGEMA_signal_14667, new_AGEMA_signal_14666, mcs1_mcs_mat1_2_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_15982, new_AGEMA_signal_15981, new_AGEMA_signal_15980, mcs1_mcs_mat1_2_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({new_AGEMA_signal_14671, new_AGEMA_signal_14670, new_AGEMA_signal_14669, mcs1_mcs_mat1_2_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_15985, new_AGEMA_signal_15984, new_AGEMA_signal_15983, mcs1_mcs_mat1_2_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_10717, new_AGEMA_signal_10716, new_AGEMA_signal_10715, mcs1_mcs_mat1_2_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_14668, new_AGEMA_signal_14667, new_AGEMA_signal_14666, mcs1_mcs_mat1_2_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_15988, new_AGEMA_signal_15987, new_AGEMA_signal_15986, mcs1_mcs_mat1_2_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_9574, new_AGEMA_signal_9573, new_AGEMA_signal_9572, mcs1_mcs_mat1_2_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_13225, new_AGEMA_signal_13224, new_AGEMA_signal_13223, mcs1_mcs_mat1_2_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_14668, new_AGEMA_signal_14667, new_AGEMA_signal_14666, mcs1_mcs_mat1_2_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_11776, new_AGEMA_signal_11775, new_AGEMA_signal_11774, mcs1_mcs_mat1_2_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_14671, new_AGEMA_signal_14670, new_AGEMA_signal_14669, mcs1_mcs_mat1_2_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_15991, new_AGEMA_signal_15990, new_AGEMA_signal_15989, mcs1_mcs_mat1_2_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_13228, new_AGEMA_signal_13227, new_AGEMA_signal_13226, mcs1_mcs_mat1_2_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_14671, new_AGEMA_signal_14670, new_AGEMA_signal_14669, mcs1_mcs_mat1_2_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_10717, new_AGEMA_signal_10716, new_AGEMA_signal_10715, mcs1_mcs_mat1_2_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_11779, new_AGEMA_signal_11778, new_AGEMA_signal_11777, mcs1_mcs_mat1_2_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_13228, new_AGEMA_signal_13227, new_AGEMA_signal_13226, mcs1_mcs_mat1_2_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .c ({new_AGEMA_signal_11779, new_AGEMA_signal_11778, new_AGEMA_signal_11777, mcs1_mcs_mat1_2_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756]}), .c ({new_AGEMA_signal_9574, new_AGEMA_signal_9573, new_AGEMA_signal_9572, mcs1_mcs_mat1_2_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762]}), .c ({new_AGEMA_signal_10717, new_AGEMA_signal_10716, new_AGEMA_signal_10715, mcs1_mcs_mat1_2_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_13234, new_AGEMA_signal_13233, new_AGEMA_signal_13232, mcs1_mcs_mat1_2_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_13231, new_AGEMA_signal_13230, new_AGEMA_signal_13229, mcs1_mcs_mat1_2_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_14674, new_AGEMA_signal_14673, new_AGEMA_signal_14672, mcs1_mcs_mat1_2_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_13231, new_AGEMA_signal_13230, new_AGEMA_signal_13229, mcs1_mcs_mat1_2_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_10720, new_AGEMA_signal_10719, new_AGEMA_signal_10718, mcs1_mcs_mat1_2_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_14677, new_AGEMA_signal_14676, new_AGEMA_signal_14675, mcs1_mcs_mat1_2_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_9577, new_AGEMA_signal_9576, new_AGEMA_signal_9575, mcs1_mcs_mat1_2_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .c ({new_AGEMA_signal_10720, new_AGEMA_signal_10719, new_AGEMA_signal_10718, mcs1_mcs_mat1_2_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({new_AGEMA_signal_13231, new_AGEMA_signal_13230, new_AGEMA_signal_13229, mcs1_mcs_mat1_2_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_14680, new_AGEMA_signal_14679, new_AGEMA_signal_14678, mcs1_mcs_mat1_2_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_11785, new_AGEMA_signal_11784, new_AGEMA_signal_11783, mcs1_mcs_mat1_2_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_8773, new_AGEMA_signal_8772, new_AGEMA_signal_8771, mcs1_mcs_mat1_2_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_13231, new_AGEMA_signal_13230, new_AGEMA_signal_13229, mcs1_mcs_mat1_2_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_14683, new_AGEMA_signal_14682, new_AGEMA_signal_14681, mcs1_mcs_mat1_2_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_15994, new_AGEMA_signal_15993, new_AGEMA_signal_15992, mcs1_mcs_mat1_2_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_13234, new_AGEMA_signal_13233, new_AGEMA_signal_13232, mcs1_mcs_mat1_2_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_11785, new_AGEMA_signal_11784, new_AGEMA_signal_11783, mcs1_mcs_mat1_2_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_14683, new_AGEMA_signal_14682, new_AGEMA_signal_14681, mcs1_mcs_mat1_2_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_11782, new_AGEMA_signal_11781, new_AGEMA_signal_11780, mcs1_mcs_mat1_2_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .c ({new_AGEMA_signal_13234, new_AGEMA_signal_13233, new_AGEMA_signal_13232, mcs1_mcs_mat1_2_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_9577, new_AGEMA_signal_9576, new_AGEMA_signal_9575, mcs1_mcs_mat1_2_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_10723, new_AGEMA_signal_10722, new_AGEMA_signal_10721, mcs1_mcs_mat1_2_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_11782, new_AGEMA_signal_11781, new_AGEMA_signal_11780, mcs1_mcs_mat1_2_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768]}), .c ({new_AGEMA_signal_11785, new_AGEMA_signal_11784, new_AGEMA_signal_11783, mcs1_mcs_mat1_2_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774]}), .c ({new_AGEMA_signal_9577, new_AGEMA_signal_9576, new_AGEMA_signal_9575, mcs1_mcs_mat1_2_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({new_AGEMA_signal_10723, new_AGEMA_signal_10722, new_AGEMA_signal_10721, mcs1_mcs_mat1_2_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_16858, new_AGEMA_signal_16857, new_AGEMA_signal_16856, mcs1_mcs_mat1_2_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_18277, new_AGEMA_signal_18276, new_AGEMA_signal_18275, mcs1_mcs_mat1_2_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_18928, new_AGEMA_signal_18927, new_AGEMA_signal_18926, mcs1_mcs_mat1_2_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_17581, new_AGEMA_signal_17580, new_AGEMA_signal_17579, mcs1_mcs_mat1_2_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_18277, new_AGEMA_signal_18276, new_AGEMA_signal_18275, mcs1_mcs_mat1_2_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_17575, new_AGEMA_signal_17574, new_AGEMA_signal_17573, mcs1_mcs_mat1_2_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_16861, new_AGEMA_signal_16860, new_AGEMA_signal_16859, mcs1_mcs_mat1_2_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_18280, new_AGEMA_signal_18279, new_AGEMA_signal_18278, mcs1_mcs_mat1_2_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_17578, new_AGEMA_signal_17577, new_AGEMA_signal_17576, mcs1_mcs_mat1_2_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_18283, new_AGEMA_signal_18282, new_AGEMA_signal_18281, mcs1_mcs_mat1_2_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_18931, new_AGEMA_signal_18930, new_AGEMA_signal_18929, mcs1_mcs_mat1_2_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_13237, new_AGEMA_signal_13236, new_AGEMA_signal_13235, mcs1_mcs_mat1_2_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_17581, new_AGEMA_signal_17580, new_AGEMA_signal_17579, mcs1_mcs_mat1_2_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_18283, new_AGEMA_signal_18282, new_AGEMA_signal_18281, mcs1_mcs_mat1_2_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_14686, new_AGEMA_signal_14685, new_AGEMA_signal_14684, mcs1_mcs_mat1_2_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .c ({new_AGEMA_signal_17578, new_AGEMA_signal_17577, new_AGEMA_signal_17576, mcs1_mcs_mat1_2_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786]}), .c ({new_AGEMA_signal_17581, new_AGEMA_signal_17580, new_AGEMA_signal_17579, mcs1_mcs_mat1_2_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792]}), .c ({new_AGEMA_signal_14686, new_AGEMA_signal_14685, new_AGEMA_signal_14684, mcs1_mcs_mat1_2_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798]}), .c ({new_AGEMA_signal_16861, new_AGEMA_signal_16860, new_AGEMA_signal_16859, mcs1_mcs_mat1_2_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_16864, new_AGEMA_signal_16863, new_AGEMA_signal_16862, mcs1_mcs_mat1_2_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_10729, new_AGEMA_signal_10728, new_AGEMA_signal_10727, mcs1_mcs_mat1_2_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_17584, new_AGEMA_signal_17583, new_AGEMA_signal_17582, mcs1_mcs_mat1_2_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_15997, new_AGEMA_signal_15996, new_AGEMA_signal_15995, mcs1_mcs_mat1_2_mcs_out[99]}), .b ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .c ({new_AGEMA_signal_16864, new_AGEMA_signal_16863, new_AGEMA_signal_16862, mcs1_mcs_mat1_2_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_14689, new_AGEMA_signal_14688, new_AGEMA_signal_14687, mcs1_mcs_mat1_2_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .c ({new_AGEMA_signal_15997, new_AGEMA_signal_15996, new_AGEMA_signal_15995, mcs1_mcs_mat1_2_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_13240, new_AGEMA_signal_13239, new_AGEMA_signal_13238, mcs1_mcs_mat1_2_mcs_out[98]}), .b ({new_AGEMA_signal_9583, new_AGEMA_signal_9582, new_AGEMA_signal_9581, mcs1_mcs_mat1_2_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_14689, new_AGEMA_signal_14688, new_AGEMA_signal_14687, mcs1_mcs_mat1_2_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_9580, new_AGEMA_signal_9579, new_AGEMA_signal_9578, mcs1_mcs_mat1_2_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_11788, new_AGEMA_signal_11787, new_AGEMA_signal_11786, mcs1_mcs_mat1_2_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_13240, new_AGEMA_signal_13239, new_AGEMA_signal_13238, mcs1_mcs_mat1_2_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804]}), .c ({new_AGEMA_signal_11788, new_AGEMA_signal_11787, new_AGEMA_signal_11786, mcs1_mcs_mat1_2_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .c ({new_AGEMA_signal_9583, new_AGEMA_signal_9582, new_AGEMA_signal_9581, mcs1_mcs_mat1_2_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816]}), .c ({new_AGEMA_signal_10729, new_AGEMA_signal_10728, new_AGEMA_signal_10727, mcs1_mcs_mat1_2_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_13243, new_AGEMA_signal_13242, new_AGEMA_signal_13241, mcs1_mcs_mat1_2_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_14692, new_AGEMA_signal_14691, new_AGEMA_signal_14690, mcs1_mcs_mat1_2_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_10735, new_AGEMA_signal_10734, new_AGEMA_signal_10733, mcs1_mcs_mat1_2_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_10738, new_AGEMA_signal_10737, new_AGEMA_signal_10736, mcs1_mcs_mat1_2_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_11794, new_AGEMA_signal_11793, new_AGEMA_signal_11792, mcs1_mcs_mat1_2_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_14695, new_AGEMA_signal_14694, new_AGEMA_signal_14693, mcs1_mcs_mat1_2_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_9586, new_AGEMA_signal_9585, new_AGEMA_signal_9584, mcs1_mcs_mat1_2_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_16000, new_AGEMA_signal_15999, new_AGEMA_signal_15998, mcs1_mcs_mat1_2_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_13243, new_AGEMA_signal_13242, new_AGEMA_signal_13241, mcs1_mcs_mat1_2_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .c ({new_AGEMA_signal_14695, new_AGEMA_signal_14694, new_AGEMA_signal_14693, mcs1_mcs_mat1_2_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_8779, new_AGEMA_signal_8778, new_AGEMA_signal_8777, mcs1_mcs_mat1_2_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_11797, new_AGEMA_signal_11796, new_AGEMA_signal_11795, mcs1_mcs_mat1_2_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_13243, new_AGEMA_signal_13242, new_AGEMA_signal_13241, mcs1_mcs_mat1_2_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822]}), .c ({new_AGEMA_signal_11797, new_AGEMA_signal_11796, new_AGEMA_signal_11795, mcs1_mcs_mat1_2_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828]}), .c ({new_AGEMA_signal_9586, new_AGEMA_signal_9585, new_AGEMA_signal_9584, mcs1_mcs_mat1_2_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834]}), .c ({new_AGEMA_signal_10738, new_AGEMA_signal_10737, new_AGEMA_signal_10736, mcs1_mcs_mat1_2_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_11806, new_AGEMA_signal_11805, new_AGEMA_signal_11804, mcs1_mcs_mat1_2_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_11809, new_AGEMA_signal_11808, new_AGEMA_signal_11807, mcs1_mcs_mat1_2_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_13246, new_AGEMA_signal_13245, new_AGEMA_signal_13244, mcs1_mcs_mat1_2_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_11800, new_AGEMA_signal_11799, new_AGEMA_signal_11798, mcs1_mcs_mat1_2_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_8782, new_AGEMA_signal_8781, new_AGEMA_signal_8780, mcs1_mcs_mat1_2_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_13249, new_AGEMA_signal_13248, new_AGEMA_signal_13247, mcs1_mcs_mat1_2_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_10747, new_AGEMA_signal_10746, new_AGEMA_signal_10745, mcs1_mcs_mat1_2_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_11800, new_AGEMA_signal_11799, new_AGEMA_signal_11798, mcs1_mcs_mat1_2_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_11803, new_AGEMA_signal_11802, new_AGEMA_signal_11801, mcs1_mcs_mat1_2_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_13252, new_AGEMA_signal_13251, new_AGEMA_signal_13250, mcs1_mcs_mat1_2_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_9589, new_AGEMA_signal_9588, new_AGEMA_signal_9587, mcs1_mcs_mat1_2_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_10747, new_AGEMA_signal_10746, new_AGEMA_signal_10745, mcs1_mcs_mat1_2_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_11803, new_AGEMA_signal_11802, new_AGEMA_signal_11801, mcs1_mcs_mat1_2_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_13255, new_AGEMA_signal_13254, new_AGEMA_signal_13253, mcs1_mcs_mat1_2_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .c ({new_AGEMA_signal_14698, new_AGEMA_signal_14697, new_AGEMA_signal_14696, mcs1_mcs_mat1_2_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_11806, new_AGEMA_signal_11805, new_AGEMA_signal_11804, mcs1_mcs_mat1_2_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_9589, new_AGEMA_signal_9588, new_AGEMA_signal_9587, mcs1_mcs_mat1_2_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_13255, new_AGEMA_signal_13254, new_AGEMA_signal_13253, mcs1_mcs_mat1_2_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({new_AGEMA_signal_11809, new_AGEMA_signal_11808, new_AGEMA_signal_11807, mcs1_mcs_mat1_2_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846]}), .c ({new_AGEMA_signal_9589, new_AGEMA_signal_9588, new_AGEMA_signal_9587, mcs1_mcs_mat1_2_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852]}), .c ({new_AGEMA_signal_10747, new_AGEMA_signal_10746, new_AGEMA_signal_10745, mcs1_mcs_mat1_2_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_13258, new_AGEMA_signal_13257, new_AGEMA_signal_13256, mcs1_mcs_mat1_2_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_14701, new_AGEMA_signal_14700, new_AGEMA_signal_14699, mcs1_mcs_mat1_2_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_10750, new_AGEMA_signal_10749, new_AGEMA_signal_10748, mcs1_mcs_mat1_2_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_11812, new_AGEMA_signal_11811, new_AGEMA_signal_11810, mcs1_mcs_mat1_2_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_14704, new_AGEMA_signal_14703, new_AGEMA_signal_14702, mcs1_mcs_mat1_2_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_9595, new_AGEMA_signal_9594, new_AGEMA_signal_9593, mcs1_mcs_mat1_2_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_16003, new_AGEMA_signal_16002, new_AGEMA_signal_16001, mcs1_mcs_mat1_2_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_13258, new_AGEMA_signal_13257, new_AGEMA_signal_13256, mcs1_mcs_mat1_2_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .c ({new_AGEMA_signal_14704, new_AGEMA_signal_14703, new_AGEMA_signal_14702, mcs1_mcs_mat1_2_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_8785, new_AGEMA_signal_8784, new_AGEMA_signal_8783, mcs1_mcs_mat1_2_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_11815, new_AGEMA_signal_11814, new_AGEMA_signal_11813, mcs1_mcs_mat1_2_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_13258, new_AGEMA_signal_13257, new_AGEMA_signal_13256, mcs1_mcs_mat1_2_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858]}), .c ({new_AGEMA_signal_11815, new_AGEMA_signal_11814, new_AGEMA_signal_11813, mcs1_mcs_mat1_2_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864]}), .c ({new_AGEMA_signal_9595, new_AGEMA_signal_9594, new_AGEMA_signal_9593, mcs1_mcs_mat1_2_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .c ({new_AGEMA_signal_10750, new_AGEMA_signal_10749, new_AGEMA_signal_10748, mcs1_mcs_mat1_2_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_14707, new_AGEMA_signal_14706, new_AGEMA_signal_14705, mcs1_mcs_mat1_2_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_16006, new_AGEMA_signal_16005, new_AGEMA_signal_16004, mcs1_mcs_mat1_2_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_13264, new_AGEMA_signal_13263, new_AGEMA_signal_13262, mcs1_mcs_mat1_2_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_11821, new_AGEMA_signal_11820, new_AGEMA_signal_11819, mcs1_mcs_mat1_2_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_14707, new_AGEMA_signal_14706, new_AGEMA_signal_14705, mcs1_mcs_mat1_2_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, new_AGEMA_signal_10298, mcs1_mcs_mat1_2_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_11818, new_AGEMA_signal_11817, new_AGEMA_signal_11816, mcs1_mcs_mat1_2_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_11821, new_AGEMA_signal_11820, new_AGEMA_signal_11819, mcs1_mcs_mat1_2_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, new_AGEMA_signal_10298, mcs1_mcs_mat1_2_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_13261, new_AGEMA_signal_13260, new_AGEMA_signal_13259, mcs1_mcs_mat1_2_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_9598, new_AGEMA_signal_9597, new_AGEMA_signal_9596, mcs1_mcs_mat1_2_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_9601, new_AGEMA_signal_9600, new_AGEMA_signal_9599, mcs1_mcs_mat1_2_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_10300, new_AGEMA_signal_10299, new_AGEMA_signal_10298, mcs1_mcs_mat1_2_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_10753, new_AGEMA_signal_10752, new_AGEMA_signal_10751, mcs1_mcs_mat1_2_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .c ({new_AGEMA_signal_11821, new_AGEMA_signal_11820, new_AGEMA_signal_11819, mcs1_mcs_mat1_2_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_14710, new_AGEMA_signal_14709, new_AGEMA_signal_14708, mcs1_mcs_mat1_2_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_9598, new_AGEMA_signal_9597, new_AGEMA_signal_9596, mcs1_mcs_mat1_2_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_16009, new_AGEMA_signal_16008, new_AGEMA_signal_16007, mcs1_mcs_mat1_2_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_13264, new_AGEMA_signal_13263, new_AGEMA_signal_13262, mcs1_mcs_mat1_2_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_10753, new_AGEMA_signal_10752, new_AGEMA_signal_10751, mcs1_mcs_mat1_2_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_14710, new_AGEMA_signal_14709, new_AGEMA_signal_14708, mcs1_mcs_mat1_2_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .b ({new_AGEMA_signal_11824, new_AGEMA_signal_11823, new_AGEMA_signal_11822, mcs1_mcs_mat1_2_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_13264, new_AGEMA_signal_13263, new_AGEMA_signal_13262, mcs1_mcs_mat1_2_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876]}), .c ({new_AGEMA_signal_11824, new_AGEMA_signal_11823, new_AGEMA_signal_11822, mcs1_mcs_mat1_2_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882]}), .c ({new_AGEMA_signal_9601, new_AGEMA_signal_9600, new_AGEMA_signal_9599, mcs1_mcs_mat1_2_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888]}), .c ({new_AGEMA_signal_10753, new_AGEMA_signal_10752, new_AGEMA_signal_10751, mcs1_mcs_mat1_2_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_18289, new_AGEMA_signal_18288, new_AGEMA_signal_18287, mcs1_mcs_mat1_2_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_16867, new_AGEMA_signal_16866, new_AGEMA_signal_16865, mcs1_mcs_mat1_2_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_18934, new_AGEMA_signal_18933, new_AGEMA_signal_18932, mcs1_mcs_mat1_2_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_17593, new_AGEMA_signal_17592, new_AGEMA_signal_17591, mcs1_mcs_mat1_2_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_18937, new_AGEMA_signal_18936, new_AGEMA_signal_18935, mcs1_mcs_mat1_2_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_19663, new_AGEMA_signal_19662, new_AGEMA_signal_19661, mcs1_mcs_mat1_2_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_18289, new_AGEMA_signal_18288, new_AGEMA_signal_18287, mcs1_mcs_mat1_2_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_18937, new_AGEMA_signal_18936, new_AGEMA_signal_18935, mcs1_mcs_mat1_2_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_19666, new_AGEMA_signal_19665, new_AGEMA_signal_19664, mcs1_mcs_mat1_2_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_16867, new_AGEMA_signal_16866, new_AGEMA_signal_16865, mcs1_mcs_mat1_2_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_18292, new_AGEMA_signal_18291, new_AGEMA_signal_18290, mcs1_mcs_mat1_2_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_18937, new_AGEMA_signal_18936, new_AGEMA_signal_18935, mcs1_mcs_mat1_2_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({new_AGEMA_signal_14713, new_AGEMA_signal_14712, new_AGEMA_signal_14711, mcs1_mcs_mat1_2_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_16867, new_AGEMA_signal_16866, new_AGEMA_signal_16865, mcs1_mcs_mat1_2_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_17590, new_AGEMA_signal_17589, new_AGEMA_signal_17588, mcs1_mcs_mat1_2_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .c ({new_AGEMA_signal_18289, new_AGEMA_signal_18288, new_AGEMA_signal_18287, mcs1_mcs_mat1_2_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_16870, new_AGEMA_signal_16869, new_AGEMA_signal_16868, mcs1_mcs_mat1_2_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_13267, new_AGEMA_signal_13266, new_AGEMA_signal_13265, mcs1_mcs_mat1_2_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_17590, new_AGEMA_signal_17589, new_AGEMA_signal_17588, mcs1_mcs_mat1_2_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_18292, new_AGEMA_signal_18291, new_AGEMA_signal_18290, mcs1_mcs_mat1_2_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_17593, new_AGEMA_signal_17592, new_AGEMA_signal_17591, mcs1_mcs_mat1_2_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_18940, new_AGEMA_signal_18939, new_AGEMA_signal_18938, mcs1_mcs_mat1_2_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_16870, new_AGEMA_signal_16869, new_AGEMA_signal_16868, mcs1_mcs_mat1_2_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_17593, new_AGEMA_signal_17592, new_AGEMA_signal_17591, mcs1_mcs_mat1_2_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({new_AGEMA_signal_17596, new_AGEMA_signal_17595, new_AGEMA_signal_17594, mcs1_mcs_mat1_2_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_18292, new_AGEMA_signal_18291, new_AGEMA_signal_18290, mcs1_mcs_mat1_2_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894]}), .c ({new_AGEMA_signal_17596, new_AGEMA_signal_17595, new_AGEMA_signal_17594, mcs1_mcs_mat1_2_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({new_AGEMA_signal_14713, new_AGEMA_signal_14712, new_AGEMA_signal_14711, mcs1_mcs_mat1_2_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906]}), .c ({new_AGEMA_signal_16870, new_AGEMA_signal_16869, new_AGEMA_signal_16868, mcs1_mcs_mat1_2_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_14719, new_AGEMA_signal_14718, new_AGEMA_signal_14717, mcs1_mcs_mat1_2_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .c ({new_AGEMA_signal_16012, new_AGEMA_signal_16011, new_AGEMA_signal_16010, mcs1_mcs_mat1_2_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({new_AGEMA_signal_13270, new_AGEMA_signal_13269, new_AGEMA_signal_13268, mcs1_mcs_mat1_2_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_14716, new_AGEMA_signal_14715, new_AGEMA_signal_14714, mcs1_mcs_mat1_2_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_16015, new_AGEMA_signal_16014, new_AGEMA_signal_16013, mcs1_mcs_mat1_2_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_10756, new_AGEMA_signal_10755, new_AGEMA_signal_10754, mcs1_mcs_mat1_2_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_16873, new_AGEMA_signal_16872, new_AGEMA_signal_16871, mcs1_mcs_mat1_2_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_14719, new_AGEMA_signal_14718, new_AGEMA_signal_14717, mcs1_mcs_mat1_2_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .c ({new_AGEMA_signal_16015, new_AGEMA_signal_16014, new_AGEMA_signal_16013, mcs1_mcs_mat1_2_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_9604, new_AGEMA_signal_9603, new_AGEMA_signal_9602, mcs1_mcs_mat1_2_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_13270, new_AGEMA_signal_13269, new_AGEMA_signal_13268, mcs1_mcs_mat1_2_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_14719, new_AGEMA_signal_14718, new_AGEMA_signal_14717, mcs1_mcs_mat1_2_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_8791, new_AGEMA_signal_8790, new_AGEMA_signal_8789, mcs1_mcs_mat1_2_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_11830, new_AGEMA_signal_11829, new_AGEMA_signal_11828, mcs1_mcs_mat1_2_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_13270, new_AGEMA_signal_13269, new_AGEMA_signal_13268, mcs1_mcs_mat1_2_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912]}), .c ({new_AGEMA_signal_11830, new_AGEMA_signal_11829, new_AGEMA_signal_11828, mcs1_mcs_mat1_2_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918]}), .c ({new_AGEMA_signal_9604, new_AGEMA_signal_9603, new_AGEMA_signal_9602, mcs1_mcs_mat1_2_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924]}), .c ({new_AGEMA_signal_10756, new_AGEMA_signal_10755, new_AGEMA_signal_10754, mcs1_mcs_mat1_2_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_13279, new_AGEMA_signal_13278, new_AGEMA_signal_13277, mcs1_mcs_mat1_2_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_10759, new_AGEMA_signal_10758, new_AGEMA_signal_10757, mcs1_mcs_mat1_2_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_14722, new_AGEMA_signal_14721, new_AGEMA_signal_14720, mcs1_mcs_mat1_2_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_9607, new_AGEMA_signal_9606, new_AGEMA_signal_9605, mcs1_mcs_mat1_2_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_11833, new_AGEMA_signal_11832, new_AGEMA_signal_11831, mcs1_mcs_mat1_2_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_13273, new_AGEMA_signal_13272, new_AGEMA_signal_13271, mcs1_mcs_mat1_2_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({new_AGEMA_signal_11836, new_AGEMA_signal_11835, new_AGEMA_signal_11834, mcs1_mcs_mat1_2_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_13276, new_AGEMA_signal_13275, new_AGEMA_signal_13274, mcs1_mcs_mat1_2_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .c ({new_AGEMA_signal_11836, new_AGEMA_signal_11835, new_AGEMA_signal_11834, mcs1_mcs_mat1_2_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936]}), .c ({new_AGEMA_signal_9607, new_AGEMA_signal_9606, new_AGEMA_signal_9605, mcs1_mcs_mat1_2_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942]}), .c ({new_AGEMA_signal_10759, new_AGEMA_signal_10758, new_AGEMA_signal_10757, mcs1_mcs_mat1_2_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_9613, new_AGEMA_signal_9612, new_AGEMA_signal_9611, mcs1_mcs_mat1_2_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_10762, new_AGEMA_signal_10761, new_AGEMA_signal_10760, mcs1_mcs_mat1_2_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_11839, new_AGEMA_signal_11838, new_AGEMA_signal_11837, mcs1_mcs_mat1_2_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_9616, new_AGEMA_signal_9615, new_AGEMA_signal_9614, mcs1_mcs_mat1_2_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_11842, new_AGEMA_signal_11841, new_AGEMA_signal_11840, mcs1_mcs_mat1_2_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_13285, new_AGEMA_signal_13284, new_AGEMA_signal_13283, mcs1_mcs_mat1_2_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_13288, new_AGEMA_signal_13287, new_AGEMA_signal_13286, mcs1_mcs_mat1_2_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_11845, new_AGEMA_signal_11844, new_AGEMA_signal_11843, mcs1_mcs_mat1_2_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_14728, new_AGEMA_signal_14727, new_AGEMA_signal_14726, mcs1_mcs_mat1_2_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_11848, new_AGEMA_signal_11847, new_AGEMA_signal_11846, mcs1_mcs_mat1_2_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_13288, new_AGEMA_signal_13287, new_AGEMA_signal_13286, mcs1_mcs_mat1_2_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948]}), .c ({new_AGEMA_signal_11848, new_AGEMA_signal_11847, new_AGEMA_signal_11846, mcs1_mcs_mat1_2_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954]}), .c ({new_AGEMA_signal_9616, new_AGEMA_signal_9615, new_AGEMA_signal_9614, mcs1_mcs_mat1_2_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({new_AGEMA_signal_10762, new_AGEMA_signal_10761, new_AGEMA_signal_10760, mcs1_mcs_mat1_2_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_17602, new_AGEMA_signal_17601, new_AGEMA_signal_17600, mcs1_mcs_mat1_2_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_18295, new_AGEMA_signal_18294, new_AGEMA_signal_18293, mcs1_mcs_mat1_2_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_18943, new_AGEMA_signal_18942, new_AGEMA_signal_18941, mcs1_mcs_mat1_2_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_18946, new_AGEMA_signal_18945, new_AGEMA_signal_18944, mcs1_mcs_mat1_2_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_17599, new_AGEMA_signal_17598, new_AGEMA_signal_17597, mcs1_mcs_mat1_2_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_19669, new_AGEMA_signal_19668, new_AGEMA_signal_19667, mcs1_mcs_mat1_2_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_16876, new_AGEMA_signal_16875, new_AGEMA_signal_16874, mcs1_mcs_mat1_2_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_17599, new_AGEMA_signal_17598, new_AGEMA_signal_17597, mcs1_mcs_mat1_2_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({new_AGEMA_signal_18946, new_AGEMA_signal_18945, new_AGEMA_signal_18944, mcs1_mcs_mat1_2_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_19672, new_AGEMA_signal_19671, new_AGEMA_signal_19670, mcs1_mcs_mat1_2_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_13291, new_AGEMA_signal_13290, new_AGEMA_signal_13289, mcs1_mcs_mat1_2_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_18295, new_AGEMA_signal_18294, new_AGEMA_signal_18293, mcs1_mcs_mat1_2_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_18946, new_AGEMA_signal_18945, new_AGEMA_signal_18944, mcs1_mcs_mat1_2_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_14731, new_AGEMA_signal_14730, new_AGEMA_signal_14729, mcs1_mcs_mat1_2_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_17608, new_AGEMA_signal_17607, new_AGEMA_signal_17606, mcs1_mcs_mat1_2_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_18295, new_AGEMA_signal_18294, new_AGEMA_signal_18293, mcs1_mcs_mat1_2_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_17605, new_AGEMA_signal_17604, new_AGEMA_signal_17603, mcs1_mcs_mat1_2_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_18298, new_AGEMA_signal_18297, new_AGEMA_signal_18296, mcs1_mcs_mat1_2_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_18949, new_AGEMA_signal_18948, new_AGEMA_signal_18947, mcs1_mcs_mat1_2_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_17602, new_AGEMA_signal_17601, new_AGEMA_signal_17600, mcs1_mcs_mat1_2_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_14731, new_AGEMA_signal_14730, new_AGEMA_signal_14729, mcs1_mcs_mat1_2_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_18298, new_AGEMA_signal_18297, new_AGEMA_signal_18296, mcs1_mcs_mat1_2_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_16876, new_AGEMA_signal_16875, new_AGEMA_signal_16874, mcs1_mcs_mat1_2_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_17602, new_AGEMA_signal_17601, new_AGEMA_signal_17600, mcs1_mcs_mat1_2_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966]}), .c ({new_AGEMA_signal_17608, new_AGEMA_signal_17607, new_AGEMA_signal_17606, mcs1_mcs_mat1_2_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972]}), .c ({new_AGEMA_signal_14731, new_AGEMA_signal_14730, new_AGEMA_signal_14729, mcs1_mcs_mat1_2_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978]}), .c ({new_AGEMA_signal_16876, new_AGEMA_signal_16875, new_AGEMA_signal_16874, mcs1_mcs_mat1_2_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_10768, new_AGEMA_signal_10767, new_AGEMA_signal_10766, mcs1_mcs_mat1_2_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_11854, new_AGEMA_signal_11853, new_AGEMA_signal_11852, mcs1_mcs_mat1_2_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_16021, new_AGEMA_signal_16020, new_AGEMA_signal_16019, mcs1_mcs_mat1_2_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_9619, new_AGEMA_signal_9618, new_AGEMA_signal_9617, mcs1_mcs_mat1_2_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_16879, new_AGEMA_signal_16878, new_AGEMA_signal_16877, mcs1_mcs_mat1_2_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_14734, new_AGEMA_signal_14733, new_AGEMA_signal_14732, mcs1_mcs_mat1_2_mcs_out[47]}), .b ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .c ({new_AGEMA_signal_16021, new_AGEMA_signal_16020, new_AGEMA_signal_16019, mcs1_mcs_mat1_2_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_13297, new_AGEMA_signal_13296, new_AGEMA_signal_13295, mcs1_mcs_mat1_2_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .c ({new_AGEMA_signal_14734, new_AGEMA_signal_14733, new_AGEMA_signal_14732, mcs1_mcs_mat1_2_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_8800, new_AGEMA_signal_8799, new_AGEMA_signal_8798, mcs1_mcs_mat1_2_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_11857, new_AGEMA_signal_11856, new_AGEMA_signal_11855, mcs1_mcs_mat1_2_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_13297, new_AGEMA_signal_13296, new_AGEMA_signal_13295, mcs1_mcs_mat1_2_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984]}), .c ({new_AGEMA_signal_11857, new_AGEMA_signal_11856, new_AGEMA_signal_11855, mcs1_mcs_mat1_2_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .c ({new_AGEMA_signal_9619, new_AGEMA_signal_9618, new_AGEMA_signal_9617, mcs1_mcs_mat1_2_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996]}), .c ({new_AGEMA_signal_10768, new_AGEMA_signal_10767, new_AGEMA_signal_10766, mcs1_mcs_mat1_2_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_13300, new_AGEMA_signal_13299, new_AGEMA_signal_13298, mcs1_mcs_mat1_2_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_10771, new_AGEMA_signal_10770, new_AGEMA_signal_10769, mcs1_mcs_mat1_2_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_14737, new_AGEMA_signal_14736, new_AGEMA_signal_14735, mcs1_mcs_mat1_2_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_11860, new_AGEMA_signal_11859, new_AGEMA_signal_11858, mcs1_mcs_mat1_2_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9622, new_AGEMA_signal_9621, new_AGEMA_signal_9620, mcs1_mcs_mat1_2_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_13300, new_AGEMA_signal_13299, new_AGEMA_signal_13298, mcs1_mcs_mat1_2_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_13303, new_AGEMA_signal_13302, new_AGEMA_signal_13301, mcs1_mcs_mat1_2_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_11866, new_AGEMA_signal_11865, new_AGEMA_signal_11864, mcs1_mcs_mat1_2_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_14740, new_AGEMA_signal_14739, new_AGEMA_signal_14738, mcs1_mcs_mat1_2_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_13306, new_AGEMA_signal_13305, new_AGEMA_signal_13304, mcs1_mcs_mat1_2_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_8803, new_AGEMA_signal_8802, new_AGEMA_signal_8801, mcs1_mcs_mat1_2_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_14743, new_AGEMA_signal_14742, new_AGEMA_signal_14741, mcs1_mcs_mat1_2_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_11860, new_AGEMA_signal_11859, new_AGEMA_signal_11858, mcs1_mcs_mat1_2_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_10774, new_AGEMA_signal_10773, new_AGEMA_signal_10772, mcs1_mcs_mat1_2_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_13306, new_AGEMA_signal_13305, new_AGEMA_signal_13304, mcs1_mcs_mat1_2_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_11863, new_AGEMA_signal_11862, new_AGEMA_signal_11861, mcs1_mcs_mat1_2_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_10774, new_AGEMA_signal_10773, new_AGEMA_signal_10772, mcs1_mcs_mat1_2_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_13309, new_AGEMA_signal_13308, new_AGEMA_signal_13307, mcs1_mcs_mat1_2_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002]}), .c ({new_AGEMA_signal_11866, new_AGEMA_signal_11865, new_AGEMA_signal_11864, mcs1_mcs_mat1_2_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008]}), .c ({new_AGEMA_signal_9622, new_AGEMA_signal_9621, new_AGEMA_signal_9620, mcs1_mcs_mat1_2_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014]}), .c ({new_AGEMA_signal_10774, new_AGEMA_signal_10773, new_AGEMA_signal_10772, mcs1_mcs_mat1_2_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_18952, new_AGEMA_signal_18951, new_AGEMA_signal_18950, mcs1_mcs_mat1_2_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_13312, new_AGEMA_signal_13311, new_AGEMA_signal_13310, mcs1_mcs_mat1_2_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_19675, new_AGEMA_signal_19674, new_AGEMA_signal_19673, mcs1_mcs_mat1_2_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_16885, new_AGEMA_signal_16884, new_AGEMA_signal_16883, mcs1_mcs_mat1_2_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_16882, new_AGEMA_signal_16881, new_AGEMA_signal_16880, mcs1_mcs_mat1_2_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_17611, new_AGEMA_signal_17610, new_AGEMA_signal_17609, mcs1_mcs_mat1_2_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({new_AGEMA_signal_18952, new_AGEMA_signal_18951, new_AGEMA_signal_18950, mcs1_mcs_mat1_2_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_19678, new_AGEMA_signal_19677, new_AGEMA_signal_19676, mcs1_mcs_mat1_2_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_17614, new_AGEMA_signal_17613, new_AGEMA_signal_17612, mcs1_mcs_mat1_2_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_18301, new_AGEMA_signal_18300, new_AGEMA_signal_18299, mcs1_mcs_mat1_2_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_18952, new_AGEMA_signal_18951, new_AGEMA_signal_18950, mcs1_mcs_mat1_2_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_17617, new_AGEMA_signal_17616, new_AGEMA_signal_17615, mcs1_mcs_mat1_2_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_16888, new_AGEMA_signal_16887, new_AGEMA_signal_16886, mcs1_mcs_mat1_2_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_18301, new_AGEMA_signal_18300, new_AGEMA_signal_18299, mcs1_mcs_mat1_2_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_17617, new_AGEMA_signal_17616, new_AGEMA_signal_17615, mcs1_mcs_mat1_2_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_16885, new_AGEMA_signal_16884, new_AGEMA_signal_16883, mcs1_mcs_mat1_2_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_18304, new_AGEMA_signal_18303, new_AGEMA_signal_18302, mcs1_mcs_mat1_2_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .b ({new_AGEMA_signal_16024, new_AGEMA_signal_16023, new_AGEMA_signal_16022, mcs1_mcs_mat1_2_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_16885, new_AGEMA_signal_16884, new_AGEMA_signal_16883, mcs1_mcs_mat1_2_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({new_AGEMA_signal_14746, new_AGEMA_signal_14745, new_AGEMA_signal_14744, mcs1_mcs_mat1_2_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_16024, new_AGEMA_signal_16023, new_AGEMA_signal_16022, mcs1_mcs_mat1_2_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({new_AGEMA_signal_17617, new_AGEMA_signal_17616, new_AGEMA_signal_17615, mcs1_mcs_mat1_2_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026]}), .c ({new_AGEMA_signal_14746, new_AGEMA_signal_14745, new_AGEMA_signal_14744, mcs1_mcs_mat1_2_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032]}), .c ({new_AGEMA_signal_16888, new_AGEMA_signal_16887, new_AGEMA_signal_16886, mcs1_mcs_mat1_2_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_11869, new_AGEMA_signal_11868, new_AGEMA_signal_11867, mcs1_mcs_mat1_2_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_10777, new_AGEMA_signal_10776, new_AGEMA_signal_10775, mcs1_mcs_mat1_2_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_13315, new_AGEMA_signal_13314, new_AGEMA_signal_13313, mcs1_mcs_mat1_2_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_9625, new_AGEMA_signal_9624, new_AGEMA_signal_9623, mcs1_mcs_mat1_2_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_10303, new_AGEMA_signal_10302, new_AGEMA_signal_10301, mcs1_mcs_mat1_2_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_16027, new_AGEMA_signal_16026, new_AGEMA_signal_16025, mcs1_mcs_mat1_2_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_11872, new_AGEMA_signal_11871, new_AGEMA_signal_11870, mcs1_mcs_mat1_2_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_16891, new_AGEMA_signal_16890, new_AGEMA_signal_16889, mcs1_mcs_mat1_2_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038]}), .c ({new_AGEMA_signal_11872, new_AGEMA_signal_11871, new_AGEMA_signal_11870, mcs1_mcs_mat1_2_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044]}), .c ({new_AGEMA_signal_9625, new_AGEMA_signal_9624, new_AGEMA_signal_9623, mcs1_mcs_mat1_2_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .c ({new_AGEMA_signal_10777, new_AGEMA_signal_10776, new_AGEMA_signal_10775, mcs1_mcs_mat1_2_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_14752, new_AGEMA_signal_14751, new_AGEMA_signal_14750, mcs1_mcs_mat1_2_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_13321, new_AGEMA_signal_13320, new_AGEMA_signal_13319, mcs1_mcs_mat1_2_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_16030, new_AGEMA_signal_16029, new_AGEMA_signal_16028, mcs1_mcs_mat1_2_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_9631, new_AGEMA_signal_9630, new_AGEMA_signal_9629, mcs1_mcs_mat1_2_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_13324, new_AGEMA_signal_13323, new_AGEMA_signal_13322, mcs1_mcs_mat1_2_mcs_out[29]}), .c ({new_AGEMA_signal_14752, new_AGEMA_signal_14751, new_AGEMA_signal_14750, mcs1_mcs_mat1_2_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_9628, new_AGEMA_signal_9627, new_AGEMA_signal_9626, mcs1_mcs_mat1_2_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_13321, new_AGEMA_signal_13320, new_AGEMA_signal_13319, mcs1_mcs_mat1_2_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_14755, new_AGEMA_signal_14754, new_AGEMA_signal_14753, mcs1_mcs_mat1_2_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_11881, new_AGEMA_signal_11880, new_AGEMA_signal_11879, mcs1_mcs_mat1_2_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .c ({new_AGEMA_signal_13321, new_AGEMA_signal_13320, new_AGEMA_signal_13319, mcs1_mcs_mat1_2_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_14758, new_AGEMA_signal_14757, new_AGEMA_signal_14756, mcs1_mcs_mat1_2_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_11875, new_AGEMA_signal_11874, new_AGEMA_signal_11873, mcs1_mcs_mat1_2_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_16033, new_AGEMA_signal_16032, new_AGEMA_signal_16031, mcs1_mcs_mat1_2_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_13327, new_AGEMA_signal_13326, new_AGEMA_signal_13325, mcs1_mcs_mat1_2_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_11878, new_AGEMA_signal_11877, new_AGEMA_signal_11876, mcs1_mcs_mat1_2_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_14758, new_AGEMA_signal_14757, new_AGEMA_signal_14756, mcs1_mcs_mat1_2_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_10780, new_AGEMA_signal_10779, new_AGEMA_signal_10778, mcs1_mcs_mat1_2_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_11878, new_AGEMA_signal_11877, new_AGEMA_signal_11876, mcs1_mcs_mat1_2_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_11881, new_AGEMA_signal_11880, new_AGEMA_signal_11879, mcs1_mcs_mat1_2_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_9631, new_AGEMA_signal_9630, new_AGEMA_signal_9629, mcs1_mcs_mat1_2_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_13327, new_AGEMA_signal_13326, new_AGEMA_signal_13325, mcs1_mcs_mat1_2_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056]}), .c ({new_AGEMA_signal_11881, new_AGEMA_signal_11880, new_AGEMA_signal_11879, mcs1_mcs_mat1_2_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062]}), .c ({new_AGEMA_signal_9631, new_AGEMA_signal_9630, new_AGEMA_signal_9629, mcs1_mcs_mat1_2_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068]}), .c ({new_AGEMA_signal_10780, new_AGEMA_signal_10779, new_AGEMA_signal_10778, mcs1_mcs_mat1_2_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_11884, new_AGEMA_signal_11883, new_AGEMA_signal_11882, mcs1_mcs_mat1_2_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_13330, new_AGEMA_signal_13329, new_AGEMA_signal_13328, mcs1_mcs_mat1_2_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_10783, new_AGEMA_signal_10782, new_AGEMA_signal_10781, mcs1_mcs_mat1_2_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_9634, new_AGEMA_signal_9633, new_AGEMA_signal_9632, mcs1_mcs_mat1_2_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_11884, new_AGEMA_signal_11883, new_AGEMA_signal_11882, mcs1_mcs_mat1_2_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_13333, new_AGEMA_signal_13332, new_AGEMA_signal_13331, mcs1_mcs_mat1_2_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_14761, new_AGEMA_signal_14760, new_AGEMA_signal_14759, mcs1_mcs_mat1_2_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_11890, new_AGEMA_signal_11889, new_AGEMA_signal_11888, mcs1_mcs_mat1_2_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_9634, new_AGEMA_signal_9633, new_AGEMA_signal_9632, mcs1_mcs_mat1_2_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_13333, new_AGEMA_signal_13332, new_AGEMA_signal_13331, mcs1_mcs_mat1_2_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_14764, new_AGEMA_signal_14763, new_AGEMA_signal_14762, mcs1_mcs_mat1_2_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .c ({new_AGEMA_signal_16036, new_AGEMA_signal_16035, new_AGEMA_signal_16034, mcs1_mcs_mat1_2_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_11890, new_AGEMA_signal_11889, new_AGEMA_signal_11888, mcs1_mcs_mat1_2_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_13336, new_AGEMA_signal_13335, new_AGEMA_signal_13334, mcs1_mcs_mat1_2_mcs_out[24]}), .c ({new_AGEMA_signal_14764, new_AGEMA_signal_14763, new_AGEMA_signal_14762, mcs1_mcs_mat1_2_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_11887, new_AGEMA_signal_11886, new_AGEMA_signal_11885, mcs1_mcs_mat1_2_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .c ({new_AGEMA_signal_13336, new_AGEMA_signal_13335, new_AGEMA_signal_13334, mcs1_mcs_mat1_2_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_10783, new_AGEMA_signal_10782, new_AGEMA_signal_10781, mcs1_mcs_mat1_2_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8812, new_AGEMA_signal_8811, new_AGEMA_signal_8810, mcs1_mcs_mat1_2_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_11887, new_AGEMA_signal_11886, new_AGEMA_signal_11885, mcs1_mcs_mat1_2_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074]}), .c ({new_AGEMA_signal_11890, new_AGEMA_signal_11889, new_AGEMA_signal_11888, mcs1_mcs_mat1_2_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .c ({new_AGEMA_signal_9634, new_AGEMA_signal_9633, new_AGEMA_signal_9632, mcs1_mcs_mat1_2_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4091], Fresh[4090], Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086]}), .c ({new_AGEMA_signal_10783, new_AGEMA_signal_10782, new_AGEMA_signal_10781, mcs1_mcs_mat1_2_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_17620, new_AGEMA_signal_17619, new_AGEMA_signal_17618, mcs1_mcs_mat1_2_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .c ({new_AGEMA_signal_18307, new_AGEMA_signal_18306, new_AGEMA_signal_18305, mcs1_mcs_mat1_2_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_16894, new_AGEMA_signal_16893, new_AGEMA_signal_16892, mcs1_mcs_mat1_2_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_14767, new_AGEMA_signal_14766, new_AGEMA_signal_14765, mcs1_mcs_mat1_2_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_17620, new_AGEMA_signal_17619, new_AGEMA_signal_17618, mcs1_mcs_mat1_2_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_18310, new_AGEMA_signal_18309, new_AGEMA_signal_18308, mcs1_mcs_mat1_2_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .c ({new_AGEMA_signal_18955, new_AGEMA_signal_18954, new_AGEMA_signal_18953, mcs1_mcs_mat1_2_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_17626, new_AGEMA_signal_17625, new_AGEMA_signal_17624, mcs1_mcs_mat1_2_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_14767, new_AGEMA_signal_14766, new_AGEMA_signal_14765, mcs1_mcs_mat1_2_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_18310, new_AGEMA_signal_18309, new_AGEMA_signal_18308, mcs1_mcs_mat1_2_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_18958, new_AGEMA_signal_18957, new_AGEMA_signal_18956, mcs1_mcs_mat1_2_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_11395, new_AGEMA_signal_11394, new_AGEMA_signal_11393, mcs1_mcs_mat1_2_mcs_out[86]}), .c ({new_AGEMA_signal_19681, new_AGEMA_signal_19680, new_AGEMA_signal_19679, mcs1_mcs_mat1_2_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_17626, new_AGEMA_signal_17625, new_AGEMA_signal_17624, mcs1_mcs_mat1_2_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_18313, new_AGEMA_signal_18312, new_AGEMA_signal_18311, mcs1_mcs_mat1_2_mcs_out[20]}), .c ({new_AGEMA_signal_18958, new_AGEMA_signal_18957, new_AGEMA_signal_18956, mcs1_mcs_mat1_2_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_17623, new_AGEMA_signal_17622, new_AGEMA_signal_17621, mcs1_mcs_mat1_2_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .c ({new_AGEMA_signal_18313, new_AGEMA_signal_18312, new_AGEMA_signal_18311, mcs1_mcs_mat1_2_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_16894, new_AGEMA_signal_16893, new_AGEMA_signal_16892, mcs1_mcs_mat1_2_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_13339, new_AGEMA_signal_13338, new_AGEMA_signal_13337, mcs1_mcs_mat1_2_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_17623, new_AGEMA_signal_17622, new_AGEMA_signal_17621, mcs1_mcs_mat1_2_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092]}), .c ({new_AGEMA_signal_17626, new_AGEMA_signal_17625, new_AGEMA_signal_17624, mcs1_mcs_mat1_2_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100], Fresh[4099], Fresh[4098]}), .c ({new_AGEMA_signal_14767, new_AGEMA_signal_14766, new_AGEMA_signal_14765, mcs1_mcs_mat1_2_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104]}), .c ({new_AGEMA_signal_16894, new_AGEMA_signal_16893, new_AGEMA_signal_16892, mcs1_mcs_mat1_2_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_11893, new_AGEMA_signal_11892, new_AGEMA_signal_11891, mcs1_mcs_mat1_2_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_11902, new_AGEMA_signal_11901, new_AGEMA_signal_11900, mcs1_mcs_mat1_2_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_13342, new_AGEMA_signal_13341, new_AGEMA_signal_13340, mcs1_mcs_mat1_2_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_13345, new_AGEMA_signal_13344, new_AGEMA_signal_13343, mcs1_mcs_mat1_2_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_8815, new_AGEMA_signal_8814, new_AGEMA_signal_8813, mcs1_mcs_mat1_2_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_14770, new_AGEMA_signal_14769, new_AGEMA_signal_14768, mcs1_mcs_mat1_2_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_14773, new_AGEMA_signal_14772, new_AGEMA_signal_14771, mcs1_mcs_mat1_2_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_9637, new_AGEMA_signal_9636, new_AGEMA_signal_9635, mcs1_mcs_mat1_2_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_16039, new_AGEMA_signal_16038, new_AGEMA_signal_16037, mcs1_mcs_mat1_2_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_8428, new_AGEMA_signal_8427, new_AGEMA_signal_8426, mcs1_mcs_mat1_2_mcs_out[50]}), .b ({new_AGEMA_signal_13345, new_AGEMA_signal_13344, new_AGEMA_signal_13343, mcs1_mcs_mat1_2_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_14773, new_AGEMA_signal_14772, new_AGEMA_signal_14771, mcs1_mcs_mat1_2_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_11896, new_AGEMA_signal_11895, new_AGEMA_signal_11894, mcs1_mcs_mat1_2_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .c ({new_AGEMA_signal_13345, new_AGEMA_signal_13344, new_AGEMA_signal_13343, mcs1_mcs_mat1_2_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_10786, new_AGEMA_signal_10785, new_AGEMA_signal_10784, mcs1_mcs_mat1_2_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_10789, new_AGEMA_signal_10788, new_AGEMA_signal_10787, mcs1_mcs_mat1_2_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_11896, new_AGEMA_signal_11895, new_AGEMA_signal_11894, mcs1_mcs_mat1_2_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_11899, new_AGEMA_signal_11898, new_AGEMA_signal_11897, mcs1_mcs_mat1_2_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_9637, new_AGEMA_signal_9636, new_AGEMA_signal_9635, mcs1_mcs_mat1_2_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_13348, new_AGEMA_signal_13347, new_AGEMA_signal_13346, mcs1_mcs_mat1_2_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110]}), .c ({new_AGEMA_signal_11902, new_AGEMA_signal_11901, new_AGEMA_signal_11900, mcs1_mcs_mat1_2_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4121], Fresh[4120], Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116]}), .c ({new_AGEMA_signal_9637, new_AGEMA_signal_9636, new_AGEMA_signal_9635, mcs1_mcs_mat1_2_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122]}), .c ({new_AGEMA_signal_10789, new_AGEMA_signal_10788, new_AGEMA_signal_10787, mcs1_mcs_mat1_2_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_14782, new_AGEMA_signal_14781, new_AGEMA_signal_14780, mcs1_mcs_mat1_2_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, new_AGEMA_signal_10304, mcs1_mcs_mat1_2_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_16042, new_AGEMA_signal_16041, new_AGEMA_signal_16040, mcs1_mcs_mat1_2_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_13357, new_AGEMA_signal_13356, new_AGEMA_signal_13355, mcs1_mcs_mat1_2_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_13351, new_AGEMA_signal_13350, new_AGEMA_signal_13349, mcs1_mcs_mat1_2_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_14776, new_AGEMA_signal_14775, new_AGEMA_signal_14774, mcs1_mcs_mat1_2_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_11908, new_AGEMA_signal_11907, new_AGEMA_signal_11906, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_9640, new_AGEMA_signal_9639, new_AGEMA_signal_9638, mcs1_mcs_mat1_2_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_13351, new_AGEMA_signal_13350, new_AGEMA_signal_13349, mcs1_mcs_mat1_2_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, new_AGEMA_signal_10304, mcs1_mcs_mat1_2_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_13354, new_AGEMA_signal_13353, new_AGEMA_signal_13352, mcs1_mcs_mat1_2_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_14779, new_AGEMA_signal_14778, new_AGEMA_signal_14777, mcs1_mcs_mat1_2_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_11905, new_AGEMA_signal_11904, new_AGEMA_signal_11903, mcs1_mcs_mat1_2_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_11908, new_AGEMA_signal_11907, new_AGEMA_signal_11906, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_13354, new_AGEMA_signal_13353, new_AGEMA_signal_13352, mcs1_mcs_mat1_2_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_8818, new_AGEMA_signal_8817, new_AGEMA_signal_8816, mcs1_mcs_mat1_2_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_9640, new_AGEMA_signal_9639, new_AGEMA_signal_9638, mcs1_mcs_mat1_2_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_10306, new_AGEMA_signal_10305, new_AGEMA_signal_10304, mcs1_mcs_mat1_2_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_16045, new_AGEMA_signal_16044, new_AGEMA_signal_16043, mcs1_mcs_mat1_2_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .c ({new_AGEMA_signal_16897, new_AGEMA_signal_16896, new_AGEMA_signal_16895, mcs1_mcs_mat1_2_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_14782, new_AGEMA_signal_14781, new_AGEMA_signal_14780, mcs1_mcs_mat1_2_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_11908, new_AGEMA_signal_11907, new_AGEMA_signal_11906, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_16045, new_AGEMA_signal_16044, new_AGEMA_signal_16043, mcs1_mcs_mat1_2_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({new_AGEMA_signal_13357, new_AGEMA_signal_13356, new_AGEMA_signal_13355, mcs1_mcs_mat1_2_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_14782, new_AGEMA_signal_14781, new_AGEMA_signal_14780, mcs1_mcs_mat1_2_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({new_AGEMA_signal_11905, new_AGEMA_signal_11904, new_AGEMA_signal_11903, mcs1_mcs_mat1_2_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_13357, new_AGEMA_signal_13356, new_AGEMA_signal_13355, mcs1_mcs_mat1_2_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_8374, new_AGEMA_signal_8373, new_AGEMA_signal_8372, shiftr_out[116]}), .b ({new_AGEMA_signal_10792, new_AGEMA_signal_10791, new_AGEMA_signal_10790, mcs1_mcs_mat1_2_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_11905, new_AGEMA_signal_11904, new_AGEMA_signal_11903, mcs1_mcs_mat1_2_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10414, new_AGEMA_signal_10413, new_AGEMA_signal_10412, mcs1_mcs_mat1_2_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130], Fresh[4129], Fresh[4128]}), .c ({new_AGEMA_signal_11908, new_AGEMA_signal_11907, new_AGEMA_signal_11906, mcs1_mcs_mat1_2_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8578, new_AGEMA_signal_8577, new_AGEMA_signal_8576, mcs1_mcs_mat1_2_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134]}), .c ({new_AGEMA_signal_9640, new_AGEMA_signal_9639, new_AGEMA_signal_9638, mcs1_mcs_mat1_2_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10216, new_AGEMA_signal_10215, new_AGEMA_signal_10214, mcs1_mcs_mat1_2_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140]}), .c ({new_AGEMA_signal_10792, new_AGEMA_signal_10791, new_AGEMA_signal_10790, mcs1_mcs_mat1_2_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_10309, new_AGEMA_signal_10308, new_AGEMA_signal_10307, mcs1_mcs_mat1_2_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .c ({new_AGEMA_signal_10795, new_AGEMA_signal_10794, new_AGEMA_signal_10793, mcs1_mcs_mat1_2_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_13363, new_AGEMA_signal_13362, new_AGEMA_signal_13361, mcs1_mcs_mat1_2_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .c ({new_AGEMA_signal_14785, new_AGEMA_signal_14784, new_AGEMA_signal_14783, mcs1_mcs_mat1_2_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_11911, new_AGEMA_signal_11910, new_AGEMA_signal_11909, mcs1_mcs_mat1_2_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .c ({new_AGEMA_signal_13360, new_AGEMA_signal_13359, new_AGEMA_signal_13358, mcs1_mcs_mat1_2_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_10798, new_AGEMA_signal_10797, new_AGEMA_signal_10796, mcs1_mcs_mat1_2_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_10309, new_AGEMA_signal_10308, new_AGEMA_signal_10307, mcs1_mcs_mat1_2_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_11911, new_AGEMA_signal_11910, new_AGEMA_signal_11909, mcs1_mcs_mat1_2_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_8821, new_AGEMA_signal_8820, new_AGEMA_signal_8819, mcs1_mcs_mat1_2_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_9643, new_AGEMA_signal_9642, new_AGEMA_signal_9641, mcs1_mcs_mat1_2_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_10309, new_AGEMA_signal_10308, new_AGEMA_signal_10307, mcs1_mcs_mat1_2_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_14788, new_AGEMA_signal_14787, new_AGEMA_signal_14786, mcs1_mcs_mat1_2_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_8389, new_AGEMA_signal_8388, new_AGEMA_signal_8387, shiftr_out[84]}), .c ({new_AGEMA_signal_16048, new_AGEMA_signal_16047, new_AGEMA_signal_16046, mcs1_mcs_mat1_2_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_8821, new_AGEMA_signal_8820, new_AGEMA_signal_8819, mcs1_mcs_mat1_2_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_13363, new_AGEMA_signal_13362, new_AGEMA_signal_13361, mcs1_mcs_mat1_2_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_14788, new_AGEMA_signal_14787, new_AGEMA_signal_14786, mcs1_mcs_mat1_2_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_11914, new_AGEMA_signal_11913, new_AGEMA_signal_11912, mcs1_mcs_mat1_2_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_10798, new_AGEMA_signal_10797, new_AGEMA_signal_10796, mcs1_mcs_mat1_2_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_13363, new_AGEMA_signal_13362, new_AGEMA_signal_13361, mcs1_mcs_mat1_2_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10428, new_AGEMA_signal_10427, mcs1_mcs_mat1_2_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4151], Fresh[4150], Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146]}), .c ({new_AGEMA_signal_11914, new_AGEMA_signal_11913, new_AGEMA_signal_11912, mcs1_mcs_mat1_2_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8592, new_AGEMA_signal_8591, mcs1_mcs_mat1_2_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152]}), .c ({new_AGEMA_signal_9643, new_AGEMA_signal_9642, new_AGEMA_signal_9641, mcs1_mcs_mat1_2_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10231, new_AGEMA_signal_10230, new_AGEMA_signal_10229, shiftr_out[87]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160], Fresh[4159], Fresh[4158]}), .c ({new_AGEMA_signal_10798, new_AGEMA_signal_10797, new_AGEMA_signal_10796, mcs1_mcs_mat1_2_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_20515, new_AGEMA_signal_20514, new_AGEMA_signal_20513, mcs1_mcs_mat1_2_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_16903, new_AGEMA_signal_16902, new_AGEMA_signal_16901, mcs1_mcs_mat1_2_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_21217, new_AGEMA_signal_21216, new_AGEMA_signal_21215, mcs1_mcs_mat1_2_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_19684, new_AGEMA_signal_19683, new_AGEMA_signal_19682, mcs1_mcs_mat1_2_mcs_out[7]}), .b ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .c ({new_AGEMA_signal_20515, new_AGEMA_signal_20514, new_AGEMA_signal_20513, mcs1_mcs_mat1_2_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_18961, new_AGEMA_signal_18960, new_AGEMA_signal_18959, mcs1_mcs_mat1_2_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .c ({new_AGEMA_signal_19684, new_AGEMA_signal_19683, new_AGEMA_signal_19682, mcs1_mcs_mat1_2_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_18316, new_AGEMA_signal_18315, new_AGEMA_signal_18314, mcs1_mcs_mat1_2_mcs_out[6]}), .b ({new_AGEMA_signal_14794, new_AGEMA_signal_14793, new_AGEMA_signal_14792, mcs1_mcs_mat1_2_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_18961, new_AGEMA_signal_18960, new_AGEMA_signal_18959, mcs1_mcs_mat1_2_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_14791, new_AGEMA_signal_14790, new_AGEMA_signal_14789, mcs1_mcs_mat1_2_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_17629, new_AGEMA_signal_17628, new_AGEMA_signal_17627, mcs1_mcs_mat1_2_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_18316, new_AGEMA_signal_18315, new_AGEMA_signal_18314, mcs1_mcs_mat1_2_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16621, new_AGEMA_signal_16620, new_AGEMA_signal_16619, shiftr_out[53]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164]}), .c ({new_AGEMA_signal_17629, new_AGEMA_signal_17628, new_AGEMA_signal_17627, mcs1_mcs_mat1_2_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12835, new_AGEMA_signal_12834, new_AGEMA_signal_12833, shiftr_out[54]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170]}), .c ({new_AGEMA_signal_14794, new_AGEMA_signal_14793, new_AGEMA_signal_14792, mcs1_mcs_mat1_2_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15709, new_AGEMA_signal_15708, new_AGEMA_signal_15707, mcs1_mcs_mat1_2_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4181], Fresh[4180], Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176]}), .c ({new_AGEMA_signal_16903, new_AGEMA_signal_16902, new_AGEMA_signal_16901, mcs1_mcs_mat1_2_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_10801, new_AGEMA_signal_10800, new_AGEMA_signal_10799, mcs1_mcs_mat1_2_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_11917, new_AGEMA_signal_11916, new_AGEMA_signal_11915, mcs1_mcs_mat1_2_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_13372, new_AGEMA_signal_13371, new_AGEMA_signal_13370, mcs1_mcs_mat1_2_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .b ({new_AGEMA_signal_10804, new_AGEMA_signal_10803, new_AGEMA_signal_10802, mcs1_mcs_mat1_2_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_11917, new_AGEMA_signal_11916, new_AGEMA_signal_11915, mcs1_mcs_mat1_2_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_13375, new_AGEMA_signal_13374, new_AGEMA_signal_13373, mcs1_mcs_mat1_2_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_9646, new_AGEMA_signal_9645, new_AGEMA_signal_9644, mcs1_mcs_mat1_2_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_14797, new_AGEMA_signal_14796, new_AGEMA_signal_14795, mcs1_mcs_mat1_2_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_13378, new_AGEMA_signal_13377, new_AGEMA_signal_13376, mcs1_mcs_mat1_2_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_11923, new_AGEMA_signal_11922, new_AGEMA_signal_11921, mcs1_mcs_mat1_2_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_14800, new_AGEMA_signal_14799, new_AGEMA_signal_14798, mcs1_mcs_mat1_2_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_11926, new_AGEMA_signal_11925, new_AGEMA_signal_11924, mcs1_mcs_mat1_2_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_8824, new_AGEMA_signal_8823, new_AGEMA_signal_8822, mcs1_mcs_mat1_2_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_13378, new_AGEMA_signal_13377, new_AGEMA_signal_13376, mcs1_mcs_mat1_2_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10468, new_AGEMA_signal_10467, new_AGEMA_signal_10466, shiftr_out[21]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182]}), .c ({new_AGEMA_signal_11926, new_AGEMA_signal_11925, new_AGEMA_signal_11924, mcs1_mcs_mat1_2_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8632, new_AGEMA_signal_8631, new_AGEMA_signal_8630, shiftr_out[22]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190], Fresh[4189], Fresh[4188]}), .c ({new_AGEMA_signal_9646, new_AGEMA_signal_9645, new_AGEMA_signal_9644, mcs1_mcs_mat1_2_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_2_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10270, new_AGEMA_signal_10269, new_AGEMA_signal_10268, mcs1_mcs_mat1_2_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194]}), .c ({new_AGEMA_signal_10804, new_AGEMA_signal_10803, new_AGEMA_signal_10802, mcs1_mcs_mat1_2_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U96 ( .a ({new_AGEMA_signal_16906, new_AGEMA_signal_16905, new_AGEMA_signal_16904, mcs1_mcs_mat1_3_n128}), .b ({new_AGEMA_signal_19687, new_AGEMA_signal_19686, new_AGEMA_signal_19685, mcs1_mcs_mat1_3_n127}), .c ({temp_next_s3[81], temp_next_s2[81], temp_next_s1[81], temp_next_s0[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U95 ( .a ({new_AGEMA_signal_19030, new_AGEMA_signal_19029, new_AGEMA_signal_19028, mcs1_mcs_mat1_3_mcs_out[41]}), .b ({new_AGEMA_signal_12034, new_AGEMA_signal_12033, new_AGEMA_signal_12032, mcs1_mcs_mat1_3_mcs_out[45]}), .c ({new_AGEMA_signal_19687, new_AGEMA_signal_19686, new_AGEMA_signal_19685, mcs1_mcs_mat1_3_n127}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U94 ( .a ({new_AGEMA_signal_10315, new_AGEMA_signal_10314, new_AGEMA_signal_10313, mcs1_mcs_mat1_3_mcs_out[33]}), .b ({new_AGEMA_signal_16129, new_AGEMA_signal_16128, new_AGEMA_signal_16127, mcs1_mcs_mat1_3_mcs_out[37]}), .c ({new_AGEMA_signal_16906, new_AGEMA_signal_16905, new_AGEMA_signal_16904, mcs1_mcs_mat1_3_n128}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U93 ( .a ({new_AGEMA_signal_17632, new_AGEMA_signal_17631, new_AGEMA_signal_17630, mcs1_mcs_mat1_3_n126}), .b ({new_AGEMA_signal_18964, new_AGEMA_signal_18963, new_AGEMA_signal_18962, mcs1_mcs_mat1_3_n125}), .c ({temp_next_s3[80], temp_next_s2[80], temp_next_s1[80], temp_next_s0[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U92 ( .a ({new_AGEMA_signal_18379, new_AGEMA_signal_18378, new_AGEMA_signal_18377, mcs1_mcs_mat1_3_mcs_out[40]}), .b ({new_AGEMA_signal_16984, new_AGEMA_signal_16983, new_AGEMA_signal_16982, mcs1_mcs_mat1_3_mcs_out[44]}), .c ({new_AGEMA_signal_18964, new_AGEMA_signal_18963, new_AGEMA_signal_18962, mcs1_mcs_mat1_3_n125}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U91 ( .a ({new_AGEMA_signal_16993, new_AGEMA_signal_16992, new_AGEMA_signal_16991, mcs1_mcs_mat1_3_mcs_out[32]}), .b ({new_AGEMA_signal_13483, new_AGEMA_signal_13482, new_AGEMA_signal_13481, mcs1_mcs_mat1_3_mcs_out[36]}), .c ({new_AGEMA_signal_17632, new_AGEMA_signal_17631, new_AGEMA_signal_17630, mcs1_mcs_mat1_3_n126}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U90 ( .a ({new_AGEMA_signal_14803, new_AGEMA_signal_14802, new_AGEMA_signal_14801, mcs1_mcs_mat1_3_n124}), .b ({new_AGEMA_signal_18967, new_AGEMA_signal_18966, new_AGEMA_signal_18965, mcs1_mcs_mat1_3_n123}), .c ({temp_next_s3[51], temp_next_s2[51], temp_next_s1[51], temp_next_s0[51]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U89 ( .a ({new_AGEMA_signal_18382, new_AGEMA_signal_18381, new_AGEMA_signal_18380, mcs1_mcs_mat1_3_mcs_out[27]}), .b ({new_AGEMA_signal_16135, new_AGEMA_signal_16134, new_AGEMA_signal_16133, mcs1_mcs_mat1_3_mcs_out[31]}), .c ({new_AGEMA_signal_18967, new_AGEMA_signal_18966, new_AGEMA_signal_18965, mcs1_mcs_mat1_3_n123}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U88 ( .a ({new_AGEMA_signal_13513, new_AGEMA_signal_13512, new_AGEMA_signal_13511, mcs1_mcs_mat1_3_mcs_out[19]}), .b ({new_AGEMA_signal_13504, new_AGEMA_signal_13503, new_AGEMA_signal_13502, mcs1_mcs_mat1_3_mcs_out[23]}), .c ({new_AGEMA_signal_14803, new_AGEMA_signal_14802, new_AGEMA_signal_14801, mcs1_mcs_mat1_3_n124}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U87 ( .a ({new_AGEMA_signal_16051, new_AGEMA_signal_16050, new_AGEMA_signal_16049, mcs1_mcs_mat1_3_n122}), .b ({new_AGEMA_signal_19696, new_AGEMA_signal_19695, new_AGEMA_signal_19694, mcs1_mcs_mat1_3_n121}), .c ({temp_next_s3[50], temp_next_s2[50], temp_next_s1[50], temp_next_s0[50]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U86 ( .a ({new_AGEMA_signal_19033, new_AGEMA_signal_19032, new_AGEMA_signal_19031, mcs1_mcs_mat1_3_mcs_out[26]}), .b ({new_AGEMA_signal_14938, new_AGEMA_signal_14937, new_AGEMA_signal_14936, mcs1_mcs_mat1_3_mcs_out[30]}), .c ({new_AGEMA_signal_19696, new_AGEMA_signal_19695, new_AGEMA_signal_19694, mcs1_mcs_mat1_3_n121}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U85 ( .a ({new_AGEMA_signal_14953, new_AGEMA_signal_14952, new_AGEMA_signal_14951, mcs1_mcs_mat1_3_mcs_out[18]}), .b ({new_AGEMA_signal_14947, new_AGEMA_signal_14946, new_AGEMA_signal_14945, mcs1_mcs_mat1_3_mcs_out[22]}), .c ({new_AGEMA_signal_16051, new_AGEMA_signal_16050, new_AGEMA_signal_16049, mcs1_mcs_mat1_3_n122}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U84 ( .a ({new_AGEMA_signal_16909, new_AGEMA_signal_16908, new_AGEMA_signal_16907, mcs1_mcs_mat1_3_n120}), .b ({new_AGEMA_signal_20524, new_AGEMA_signal_20523, new_AGEMA_signal_20522, mcs1_mcs_mat1_3_n119}), .c ({temp_next_s3[49], temp_next_s2[49], temp_next_s1[49], temp_next_s0[49]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U83 ( .a ({new_AGEMA_signal_19753, new_AGEMA_signal_19752, new_AGEMA_signal_19751, mcs1_mcs_mat1_3_mcs_out[25]}), .b ({new_AGEMA_signal_13495, new_AGEMA_signal_13494, new_AGEMA_signal_13493, mcs1_mcs_mat1_3_mcs_out[29]}), .c ({new_AGEMA_signal_20524, new_AGEMA_signal_20523, new_AGEMA_signal_20522, mcs1_mcs_mat1_3_n119}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U82 ( .a ({new_AGEMA_signal_16144, new_AGEMA_signal_16143, new_AGEMA_signal_16142, mcs1_mcs_mat1_3_mcs_out[17]}), .b ({new_AGEMA_signal_16141, new_AGEMA_signal_16140, new_AGEMA_signal_16139, mcs1_mcs_mat1_3_mcs_out[21]}), .c ({new_AGEMA_signal_16909, new_AGEMA_signal_16908, new_AGEMA_signal_16907, mcs1_mcs_mat1_3_n120}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U81 ( .a ({new_AGEMA_signal_14806, new_AGEMA_signal_14805, new_AGEMA_signal_14804, mcs1_mcs_mat1_3_n118}), .b ({new_AGEMA_signal_18970, new_AGEMA_signal_18969, new_AGEMA_signal_18968, mcs1_mcs_mat1_3_n117}), .c ({temp_next_s3[48], temp_next_s2[48], temp_next_s1[48], temp_next_s0[48]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U80 ( .a ({new_AGEMA_signal_18388, new_AGEMA_signal_18387, new_AGEMA_signal_18386, mcs1_mcs_mat1_3_mcs_out[24]}), .b ({new_AGEMA_signal_16138, new_AGEMA_signal_16137, new_AGEMA_signal_16136, mcs1_mcs_mat1_3_mcs_out[28]}), .c ({new_AGEMA_signal_18970, new_AGEMA_signal_18969, new_AGEMA_signal_18968, mcs1_mcs_mat1_3_n117}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U79 ( .a ({new_AGEMA_signal_13519, new_AGEMA_signal_13518, new_AGEMA_signal_13517, mcs1_mcs_mat1_3_mcs_out[16]}), .b ({new_AGEMA_signal_13510, new_AGEMA_signal_13509, new_AGEMA_signal_13508, mcs1_mcs_mat1_3_mcs_out[20]}), .c ({new_AGEMA_signal_14806, new_AGEMA_signal_14805, new_AGEMA_signal_14804, mcs1_mcs_mat1_3_n118}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U78 ( .a ({new_AGEMA_signal_17635, new_AGEMA_signal_17634, new_AGEMA_signal_17633, mcs1_mcs_mat1_3_n116}), .b ({new_AGEMA_signal_16912, new_AGEMA_signal_16911, new_AGEMA_signal_16910, mcs1_mcs_mat1_3_n115}), .c ({temp_next_s3[19], temp_next_s2[19], temp_next_s1[19], temp_next_s0[19]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U77 ( .a ({new_AGEMA_signal_13537, new_AGEMA_signal_13536, new_AGEMA_signal_13535, mcs1_mcs_mat1_3_mcs_out[3]}), .b ({new_AGEMA_signal_16156, new_AGEMA_signal_16155, new_AGEMA_signal_16154, mcs1_mcs_mat1_3_mcs_out[7]}), .c ({new_AGEMA_signal_16912, new_AGEMA_signal_16911, new_AGEMA_signal_16910, mcs1_mcs_mat1_3_n115}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U76 ( .a ({new_AGEMA_signal_17002, new_AGEMA_signal_17001, new_AGEMA_signal_17000, mcs1_mcs_mat1_3_mcs_out[11]}), .b ({new_AGEMA_signal_16147, new_AGEMA_signal_16146, new_AGEMA_signal_16145, mcs1_mcs_mat1_3_mcs_out[15]}), .c ({new_AGEMA_signal_17635, new_AGEMA_signal_17634, new_AGEMA_signal_17633, mcs1_mcs_mat1_3_n116}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U75 ( .a ({new_AGEMA_signal_16915, new_AGEMA_signal_16914, new_AGEMA_signal_16913, mcs1_mcs_mat1_3_n114}), .b ({new_AGEMA_signal_20527, new_AGEMA_signal_20526, new_AGEMA_signal_20525, mcs1_mcs_mat1_3_n113}), .c ({new_AGEMA_signal_21223, new_AGEMA_signal_21222, new_AGEMA_signal_21221, mcs_out[243]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U74 ( .a ({new_AGEMA_signal_19738, new_AGEMA_signal_19737, new_AGEMA_signal_19736, mcs1_mcs_mat1_3_mcs_out[123]}), .b ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_20527, new_AGEMA_signal_20526, new_AGEMA_signal_20525, mcs1_mcs_mat1_3_n113}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U73 ( .a ({new_AGEMA_signal_14839, new_AGEMA_signal_14838, new_AGEMA_signal_14837, mcs1_mcs_mat1_3_mcs_out[115]}), .b ({new_AGEMA_signal_16069, new_AGEMA_signal_16068, new_AGEMA_signal_16067, mcs1_mcs_mat1_3_mcs_out[119]}), .c ({new_AGEMA_signal_16915, new_AGEMA_signal_16914, new_AGEMA_signal_16913, mcs1_mcs_mat1_3_n114}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U72 ( .a ({new_AGEMA_signal_16918, new_AGEMA_signal_16917, new_AGEMA_signal_16916, mcs1_mcs_mat1_3_n112}), .b ({new_AGEMA_signal_18322, new_AGEMA_signal_18321, new_AGEMA_signal_18320, mcs1_mcs_mat1_3_n111}), .c ({new_AGEMA_signal_18973, new_AGEMA_signal_18972, new_AGEMA_signal_18971, mcs_out[242]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U71 ( .a ({new_AGEMA_signal_17656, new_AGEMA_signal_17655, new_AGEMA_signal_17654, mcs1_mcs_mat1_3_mcs_out[122]}), .b ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_18322, new_AGEMA_signal_18321, new_AGEMA_signal_18320, mcs1_mcs_mat1_3_n111}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U70 ( .a ({new_AGEMA_signal_13390, new_AGEMA_signal_13389, new_AGEMA_signal_13388, mcs1_mcs_mat1_3_mcs_out[114]}), .b ({new_AGEMA_signal_16072, new_AGEMA_signal_16071, new_AGEMA_signal_16070, mcs1_mcs_mat1_3_mcs_out[118]}), .c ({new_AGEMA_signal_16918, new_AGEMA_signal_16917, new_AGEMA_signal_16916, mcs1_mcs_mat1_3_n112}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U69 ( .a ({new_AGEMA_signal_19702, new_AGEMA_signal_19701, new_AGEMA_signal_19700, mcs1_mcs_mat1_3_n110}), .b ({new_AGEMA_signal_14809, new_AGEMA_signal_14808, new_AGEMA_signal_14807, mcs1_mcs_mat1_3_n109}), .c ({temp_next_s3[18], temp_next_s2[18], temp_next_s1[18], temp_next_s0[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U68 ( .a ({new_AGEMA_signal_13540, new_AGEMA_signal_13539, new_AGEMA_signal_13538, mcs1_mcs_mat1_3_mcs_out[2]}), .b ({new_AGEMA_signal_13534, new_AGEMA_signal_13533, new_AGEMA_signal_13532, mcs1_mcs_mat1_3_mcs_out[6]}), .c ({new_AGEMA_signal_14809, new_AGEMA_signal_14808, new_AGEMA_signal_14807, mcs1_mcs_mat1_3_n109}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U67 ( .a ({new_AGEMA_signal_19039, new_AGEMA_signal_19038, new_AGEMA_signal_19037, mcs1_mcs_mat1_3_mcs_out[10]}), .b ({new_AGEMA_signal_14959, new_AGEMA_signal_14958, new_AGEMA_signal_14957, mcs1_mcs_mat1_3_mcs_out[14]}), .c ({new_AGEMA_signal_19702, new_AGEMA_signal_19701, new_AGEMA_signal_19700, mcs1_mcs_mat1_3_n110}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U66 ( .a ({new_AGEMA_signal_16054, new_AGEMA_signal_16053, new_AGEMA_signal_16052, mcs1_mcs_mat1_3_n108}), .b ({new_AGEMA_signal_20533, new_AGEMA_signal_20532, new_AGEMA_signal_20531, mcs1_mcs_mat1_3_n107}), .c ({new_AGEMA_signal_21226, new_AGEMA_signal_21225, new_AGEMA_signal_21224, mcs_out[241]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U65 ( .a ({new_AGEMA_signal_19741, new_AGEMA_signal_19740, new_AGEMA_signal_19739, mcs1_mcs_mat1_3_mcs_out[121]}), .b ({new_AGEMA_signal_10807, new_AGEMA_signal_10806, new_AGEMA_signal_10805, mcs1_mcs_mat1_3_mcs_out[125]}), .c ({new_AGEMA_signal_20533, new_AGEMA_signal_20532, new_AGEMA_signal_20531, mcs1_mcs_mat1_3_n107}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U64 ( .a ({new_AGEMA_signal_11938, new_AGEMA_signal_11937, new_AGEMA_signal_11936, mcs1_mcs_mat1_3_mcs_out[113]}), .b ({new_AGEMA_signal_14836, new_AGEMA_signal_14835, new_AGEMA_signal_14834, mcs1_mcs_mat1_3_mcs_out[117]}), .c ({new_AGEMA_signal_16054, new_AGEMA_signal_16053, new_AGEMA_signal_16052, mcs1_mcs_mat1_3_n108}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U63 ( .a ({new_AGEMA_signal_16921, new_AGEMA_signal_16920, new_AGEMA_signal_16919, mcs1_mcs_mat1_3_n106}), .b ({new_AGEMA_signal_19705, new_AGEMA_signal_19704, new_AGEMA_signal_19703, mcs1_mcs_mat1_3_n105}), .c ({new_AGEMA_signal_20536, new_AGEMA_signal_20535, new_AGEMA_signal_20534, mcs_out[240]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U62 ( .a ({new_AGEMA_signal_19000, new_AGEMA_signal_18999, new_AGEMA_signal_18998, mcs1_mcs_mat1_3_mcs_out[120]}), .b ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_19705, new_AGEMA_signal_19704, new_AGEMA_signal_19703, mcs1_mcs_mat1_3_n105}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U61 ( .a ({new_AGEMA_signal_16075, new_AGEMA_signal_16074, new_AGEMA_signal_16073, mcs1_mcs_mat1_3_mcs_out[112]}), .b ({new_AGEMA_signal_13387, new_AGEMA_signal_13386, new_AGEMA_signal_13385, mcs1_mcs_mat1_3_mcs_out[116]}), .c ({new_AGEMA_signal_16921, new_AGEMA_signal_16920, new_AGEMA_signal_16919, mcs1_mcs_mat1_3_n106}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U60 ( .a ({new_AGEMA_signal_19708, new_AGEMA_signal_19707, new_AGEMA_signal_19706, mcs1_mcs_mat1_3_n104}), .b ({new_AGEMA_signal_16924, new_AGEMA_signal_16923, new_AGEMA_signal_16922, mcs1_mcs_mat1_3_n103}), .c ({new_AGEMA_signal_20539, new_AGEMA_signal_20538, new_AGEMA_signal_20537, mcs_out[211]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U59 ( .a ({new_AGEMA_signal_16078, new_AGEMA_signal_16077, new_AGEMA_signal_16076, mcs1_mcs_mat1_3_mcs_out[111]}), .b ({new_AGEMA_signal_16090, new_AGEMA_signal_16089, new_AGEMA_signal_16088, mcs1_mcs_mat1_3_mcs_out[99]}), .c ({new_AGEMA_signal_16924, new_AGEMA_signal_16923, new_AGEMA_signal_16922, mcs1_mcs_mat1_3_n103}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U58 ( .a ({new_AGEMA_signal_14854, new_AGEMA_signal_14853, new_AGEMA_signal_14852, mcs1_mcs_mat1_3_mcs_out[103]}), .b ({new_AGEMA_signal_19003, new_AGEMA_signal_19002, new_AGEMA_signal_19001, mcs1_mcs_mat1_3_mcs_out[107]}), .c ({new_AGEMA_signal_19708, new_AGEMA_signal_19707, new_AGEMA_signal_19706, mcs1_mcs_mat1_3_n104}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U57 ( .a ({new_AGEMA_signal_19711, new_AGEMA_signal_19710, new_AGEMA_signal_19709, mcs1_mcs_mat1_3_n102}), .b ({new_AGEMA_signal_16927, new_AGEMA_signal_16926, new_AGEMA_signal_16925, mcs1_mcs_mat1_3_n101}), .c ({new_AGEMA_signal_20542, new_AGEMA_signal_20541, new_AGEMA_signal_20540, mcs_out[210]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U56 ( .a ({new_AGEMA_signal_16081, new_AGEMA_signal_16080, new_AGEMA_signal_16079, mcs1_mcs_mat1_3_mcs_out[110]}), .b ({new_AGEMA_signal_13417, new_AGEMA_signal_13416, new_AGEMA_signal_13415, mcs1_mcs_mat1_3_mcs_out[98]}), .c ({new_AGEMA_signal_16927, new_AGEMA_signal_16926, new_AGEMA_signal_16925, mcs1_mcs_mat1_3_n101}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U55 ( .a ({new_AGEMA_signal_11953, new_AGEMA_signal_11952, new_AGEMA_signal_11951, mcs1_mcs_mat1_3_mcs_out[102]}), .b ({new_AGEMA_signal_19006, new_AGEMA_signal_19005, new_AGEMA_signal_19004, mcs1_mcs_mat1_3_mcs_out[106]}), .c ({new_AGEMA_signal_19711, new_AGEMA_signal_19710, new_AGEMA_signal_19709, mcs1_mcs_mat1_3_n102}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U54 ( .a ({new_AGEMA_signal_19714, new_AGEMA_signal_19713, new_AGEMA_signal_19712, mcs1_mcs_mat1_3_n100}), .b ({new_AGEMA_signal_16930, new_AGEMA_signal_16929, new_AGEMA_signal_16928, mcs1_mcs_mat1_3_n99}), .c ({new_AGEMA_signal_20545, new_AGEMA_signal_20544, new_AGEMA_signal_20543, mcs_out[209]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U53 ( .a ({new_AGEMA_signal_16084, new_AGEMA_signal_16083, new_AGEMA_signal_16082, mcs1_mcs_mat1_3_mcs_out[109]}), .b ({new_AGEMA_signal_10834, new_AGEMA_signal_10833, new_AGEMA_signal_10832, mcs1_mcs_mat1_3_mcs_out[97]}), .c ({new_AGEMA_signal_16930, new_AGEMA_signal_16929, new_AGEMA_signal_16928, mcs1_mcs_mat1_3_n99}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U52 ( .a ({new_AGEMA_signal_13411, new_AGEMA_signal_13410, new_AGEMA_signal_13409, mcs1_mcs_mat1_3_mcs_out[101]}), .b ({new_AGEMA_signal_19009, new_AGEMA_signal_19008, new_AGEMA_signal_19007, mcs1_mcs_mat1_3_mcs_out[105]}), .c ({new_AGEMA_signal_19714, new_AGEMA_signal_19713, new_AGEMA_signal_19712, mcs1_mcs_mat1_3_n100}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U51 ( .a ({new_AGEMA_signal_20548, new_AGEMA_signal_20547, new_AGEMA_signal_20546, mcs1_mcs_mat1_3_n98}), .b ({new_AGEMA_signal_18325, new_AGEMA_signal_18324, new_AGEMA_signal_18323, mcs1_mcs_mat1_3_n97}), .c ({new_AGEMA_signal_21229, new_AGEMA_signal_21228, new_AGEMA_signal_21227, mcs_out[208]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U50 ( .a ({new_AGEMA_signal_16087, new_AGEMA_signal_16086, new_AGEMA_signal_16085, mcs1_mcs_mat1_3_mcs_out[108]}), .b ({new_AGEMA_signal_17668, new_AGEMA_signal_17667, new_AGEMA_signal_17666, mcs1_mcs_mat1_3_mcs_out[96]}), .c ({new_AGEMA_signal_18325, new_AGEMA_signal_18324, new_AGEMA_signal_18323, mcs1_mcs_mat1_3_n97}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U49 ( .a ({new_AGEMA_signal_14857, new_AGEMA_signal_14856, new_AGEMA_signal_14855, mcs1_mcs_mat1_3_mcs_out[100]}), .b ({new_AGEMA_signal_19744, new_AGEMA_signal_19743, new_AGEMA_signal_19742, mcs1_mcs_mat1_3_mcs_out[104]}), .c ({new_AGEMA_signal_20548, new_AGEMA_signal_20547, new_AGEMA_signal_20546, mcs1_mcs_mat1_3_n98}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U48 ( .a ({new_AGEMA_signal_14812, new_AGEMA_signal_14811, new_AGEMA_signal_14810, mcs1_mcs_mat1_3_n96}), .b ({new_AGEMA_signal_17638, new_AGEMA_signal_17637, new_AGEMA_signal_17636, mcs1_mcs_mat1_3_n95}), .c ({new_AGEMA_signal_18328, new_AGEMA_signal_18327, new_AGEMA_signal_18326, mcs_out[179]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U47 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_14863, new_AGEMA_signal_14862, new_AGEMA_signal_14861, mcs1_mcs_mat1_3_mcs_out[95]}), .c ({new_AGEMA_signal_17638, new_AGEMA_signal_17637, new_AGEMA_signal_17636, mcs1_mcs_mat1_3_n95}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U46 ( .a ({new_AGEMA_signal_13426, new_AGEMA_signal_13425, new_AGEMA_signal_13424, mcs1_mcs_mat1_3_mcs_out[83]}), .b ({new_AGEMA_signal_11977, new_AGEMA_signal_11976, new_AGEMA_signal_11975, mcs1_mcs_mat1_3_mcs_out[87]}), .c ({new_AGEMA_signal_14812, new_AGEMA_signal_14811, new_AGEMA_signal_14810, mcs1_mcs_mat1_3_n96}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U45 ( .a ({new_AGEMA_signal_14815, new_AGEMA_signal_14814, new_AGEMA_signal_14813, mcs1_mcs_mat1_3_n94}), .b ({new_AGEMA_signal_17641, new_AGEMA_signal_17640, new_AGEMA_signal_17639, mcs1_mcs_mat1_3_n93}), .c ({new_AGEMA_signal_18331, new_AGEMA_signal_18330, new_AGEMA_signal_18329, mcs_out[178]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U43 ( .a ({new_AGEMA_signal_13429, new_AGEMA_signal_13428, new_AGEMA_signal_13427, mcs1_mcs_mat1_3_mcs_out[82]}), .b ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_14815, new_AGEMA_signal_14814, new_AGEMA_signal_14813, mcs1_mcs_mat1_3_n94}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U42 ( .a ({new_AGEMA_signal_14818, new_AGEMA_signal_14817, new_AGEMA_signal_14816, mcs1_mcs_mat1_3_n92}), .b ({new_AGEMA_signal_17644, new_AGEMA_signal_17643, new_AGEMA_signal_17642, mcs1_mcs_mat1_3_n91}), .c ({new_AGEMA_signal_18334, new_AGEMA_signal_18333, new_AGEMA_signal_18332, mcs_out[177]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U41 ( .a ({new_AGEMA_signal_16972, new_AGEMA_signal_16971, new_AGEMA_signal_16970, mcs1_mcs_mat1_3_mcs_out[89]}), .b ({new_AGEMA_signal_11971, new_AGEMA_signal_11970, new_AGEMA_signal_11969, mcs1_mcs_mat1_3_mcs_out[93]}), .c ({new_AGEMA_signal_17644, new_AGEMA_signal_17643, new_AGEMA_signal_17642, mcs1_mcs_mat1_3_n91}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U40 ( .a ({new_AGEMA_signal_13432, new_AGEMA_signal_13431, new_AGEMA_signal_13430, mcs1_mcs_mat1_3_mcs_out[81]}), .b ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_14818, new_AGEMA_signal_14817, new_AGEMA_signal_14816, mcs1_mcs_mat1_3_n92}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U39 ( .a ({new_AGEMA_signal_16057, new_AGEMA_signal_16056, new_AGEMA_signal_16055, mcs1_mcs_mat1_3_n90}), .b ({new_AGEMA_signal_16933, new_AGEMA_signal_16932, new_AGEMA_signal_16931, mcs1_mcs_mat1_3_n89}), .c ({new_AGEMA_signal_17647, new_AGEMA_signal_17646, new_AGEMA_signal_17645, mcs_out[176]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U38 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_16093, new_AGEMA_signal_16092, new_AGEMA_signal_16091, mcs1_mcs_mat1_3_mcs_out[92]}), .c ({new_AGEMA_signal_16933, new_AGEMA_signal_16932, new_AGEMA_signal_16931, mcs1_mcs_mat1_3_n89}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U37 ( .a ({new_AGEMA_signal_14869, new_AGEMA_signal_14868, new_AGEMA_signal_14867, mcs1_mcs_mat1_3_mcs_out[80]}), .b ({new_AGEMA_signal_13423, new_AGEMA_signal_13422, new_AGEMA_signal_13421, mcs1_mcs_mat1_3_mcs_out[84]}), .c ({new_AGEMA_signal_16057, new_AGEMA_signal_16056, new_AGEMA_signal_16055, mcs1_mcs_mat1_3_n90}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U36 ( .a ({new_AGEMA_signal_16060, new_AGEMA_signal_16059, new_AGEMA_signal_16058, mcs1_mcs_mat1_3_n88}), .b ({new_AGEMA_signal_18976, new_AGEMA_signal_18975, new_AGEMA_signal_18974, mcs1_mcs_mat1_3_n87}), .c ({temp_next_s3[17], temp_next_s2[17], temp_next_s1[17], temp_next_s0[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U35 ( .a ({new_AGEMA_signal_10903, new_AGEMA_signal_10902, new_AGEMA_signal_10901, mcs1_mcs_mat1_3_mcs_out[5]}), .b ({new_AGEMA_signal_18391, new_AGEMA_signal_18390, new_AGEMA_signal_18389, mcs1_mcs_mat1_3_mcs_out[9]}), .c ({new_AGEMA_signal_18976, new_AGEMA_signal_18975, new_AGEMA_signal_18974, mcs1_mcs_mat1_3_n87}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U34 ( .a ({new_AGEMA_signal_14962, new_AGEMA_signal_14961, new_AGEMA_signal_14960, mcs1_mcs_mat1_3_mcs_out[13]}), .b ({new_AGEMA_signal_14974, new_AGEMA_signal_14973, new_AGEMA_signal_14972, mcs1_mcs_mat1_3_mcs_out[1]}), .c ({new_AGEMA_signal_16060, new_AGEMA_signal_16059, new_AGEMA_signal_16058, mcs1_mcs_mat1_3_n88}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U33 ( .a ({new_AGEMA_signal_16936, new_AGEMA_signal_16935, new_AGEMA_signal_16934, mcs1_mcs_mat1_3_n86}), .b ({new_AGEMA_signal_18337, new_AGEMA_signal_18336, new_AGEMA_signal_18335, mcs1_mcs_mat1_3_n85}), .c ({new_AGEMA_signal_18979, new_AGEMA_signal_18978, new_AGEMA_signal_18977, mcs_out[147]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U32 ( .a ({new_AGEMA_signal_17671, new_AGEMA_signal_17670, new_AGEMA_signal_17669, mcs1_mcs_mat1_3_mcs_out[75]}), .b ({new_AGEMA_signal_14872, new_AGEMA_signal_14871, new_AGEMA_signal_14870, mcs1_mcs_mat1_3_mcs_out[79]}), .c ({new_AGEMA_signal_18337, new_AGEMA_signal_18336, new_AGEMA_signal_18335, mcs1_mcs_mat1_3_n85}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U31 ( .a ({new_AGEMA_signal_16108, new_AGEMA_signal_16107, new_AGEMA_signal_16106, mcs1_mcs_mat1_3_mcs_out[67]}), .b ({new_AGEMA_signal_14884, new_AGEMA_signal_14883, new_AGEMA_signal_14882, mcs1_mcs_mat1_3_mcs_out[71]}), .c ({new_AGEMA_signal_16936, new_AGEMA_signal_16935, new_AGEMA_signal_16934, mcs1_mcs_mat1_3_n86}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U30 ( .a ({new_AGEMA_signal_16939, new_AGEMA_signal_16938, new_AGEMA_signal_16937, mcs1_mcs_mat1_3_n84}), .b ({new_AGEMA_signal_20551, new_AGEMA_signal_20550, new_AGEMA_signal_20549, mcs1_mcs_mat1_3_n83}), .c ({new_AGEMA_signal_21232, new_AGEMA_signal_21231, new_AGEMA_signal_21230, mcs_out[146]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U29 ( .a ({new_AGEMA_signal_19747, new_AGEMA_signal_19746, new_AGEMA_signal_19745, mcs1_mcs_mat1_3_mcs_out[74]}), .b ({new_AGEMA_signal_9676, new_AGEMA_signal_9675, new_AGEMA_signal_9674, mcs1_mcs_mat1_3_mcs_out[78]}), .c ({new_AGEMA_signal_20551, new_AGEMA_signal_20550, new_AGEMA_signal_20549, mcs1_mcs_mat1_3_n83}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U28 ( .a ({new_AGEMA_signal_14893, new_AGEMA_signal_14892, new_AGEMA_signal_14891, mcs1_mcs_mat1_3_mcs_out[66]}), .b ({new_AGEMA_signal_16102, new_AGEMA_signal_16101, new_AGEMA_signal_16100, mcs1_mcs_mat1_3_mcs_out[70]}), .c ({new_AGEMA_signal_16939, new_AGEMA_signal_16938, new_AGEMA_signal_16937, mcs1_mcs_mat1_3_n84}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U27 ( .a ({new_AGEMA_signal_16942, new_AGEMA_signal_16941, new_AGEMA_signal_16940, mcs1_mcs_mat1_3_n82}), .b ({new_AGEMA_signal_18982, new_AGEMA_signal_18981, new_AGEMA_signal_18980, mcs1_mcs_mat1_3_n81}), .c ({new_AGEMA_signal_19720, new_AGEMA_signal_19719, new_AGEMA_signal_19718, mcs_out[145]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U26 ( .a ({new_AGEMA_signal_18355, new_AGEMA_signal_18354, new_AGEMA_signal_18353, mcs1_mcs_mat1_3_mcs_out[73]}), .b ({new_AGEMA_signal_11992, new_AGEMA_signal_11991, new_AGEMA_signal_11990, mcs1_mcs_mat1_3_mcs_out[77]}), .c ({new_AGEMA_signal_18982, new_AGEMA_signal_18981, new_AGEMA_signal_18980, mcs1_mcs_mat1_3_n81}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U25 ( .a ({new_AGEMA_signal_12007, new_AGEMA_signal_12006, new_AGEMA_signal_12005, mcs1_mcs_mat1_3_mcs_out[65]}), .b ({new_AGEMA_signal_16105, new_AGEMA_signal_16104, new_AGEMA_signal_16103, mcs1_mcs_mat1_3_mcs_out[69]}), .c ({new_AGEMA_signal_16942, new_AGEMA_signal_16941, new_AGEMA_signal_16940, mcs1_mcs_mat1_3_n82}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U24 ( .a ({new_AGEMA_signal_17650, new_AGEMA_signal_17649, new_AGEMA_signal_17648, mcs1_mcs_mat1_3_n80}), .b ({new_AGEMA_signal_20554, new_AGEMA_signal_20553, new_AGEMA_signal_20552, mcs1_mcs_mat1_3_n79}), .c ({new_AGEMA_signal_21235, new_AGEMA_signal_21234, new_AGEMA_signal_21233, mcs_out[144]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U23 ( .a ({new_AGEMA_signal_19750, new_AGEMA_signal_19749, new_AGEMA_signal_19748, mcs1_mcs_mat1_3_mcs_out[72]}), .b ({new_AGEMA_signal_16096, new_AGEMA_signal_16095, new_AGEMA_signal_16094, mcs1_mcs_mat1_3_mcs_out[76]}), .c ({new_AGEMA_signal_20554, new_AGEMA_signal_20553, new_AGEMA_signal_20552, mcs1_mcs_mat1_3_n79}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U22 ( .a ({new_AGEMA_signal_16978, new_AGEMA_signal_16977, new_AGEMA_signal_16976, mcs1_mcs_mat1_3_mcs_out[64]}), .b ({new_AGEMA_signal_14890, new_AGEMA_signal_14889, new_AGEMA_signal_14888, mcs1_mcs_mat1_3_mcs_out[68]}), .c ({new_AGEMA_signal_17650, new_AGEMA_signal_17649, new_AGEMA_signal_17648, mcs1_mcs_mat1_3_n80}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U21 ( .a ({new_AGEMA_signal_16063, new_AGEMA_signal_16062, new_AGEMA_signal_16061, mcs1_mcs_mat1_3_n78}), .b ({new_AGEMA_signal_18985, new_AGEMA_signal_18984, new_AGEMA_signal_18983, mcs1_mcs_mat1_3_n77}), .c ({temp_next_s3[115], temp_next_s2[115], temp_next_s1[115], temp_next_s0[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U20 ( .a ({new_AGEMA_signal_18361, new_AGEMA_signal_18360, new_AGEMA_signal_18359, mcs1_mcs_mat1_3_mcs_out[59]}), .b ({new_AGEMA_signal_14899, new_AGEMA_signal_14898, new_AGEMA_signal_14897, mcs1_mcs_mat1_3_mcs_out[63]}), .c ({new_AGEMA_signal_18985, new_AGEMA_signal_18984, new_AGEMA_signal_18983, mcs1_mcs_mat1_3_n77}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U19 ( .a ({new_AGEMA_signal_12031, new_AGEMA_signal_12030, new_AGEMA_signal_12029, mcs1_mcs_mat1_3_mcs_out[51]}), .b ({new_AGEMA_signal_14914, new_AGEMA_signal_14913, new_AGEMA_signal_14912, mcs1_mcs_mat1_3_mcs_out[55]}), .c ({new_AGEMA_signal_16063, new_AGEMA_signal_16062, new_AGEMA_signal_16061, mcs1_mcs_mat1_3_n78}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U18 ( .a ({new_AGEMA_signal_16945, new_AGEMA_signal_16944, new_AGEMA_signal_16943, mcs1_mcs_mat1_3_n76}), .b ({new_AGEMA_signal_18340, new_AGEMA_signal_18339, new_AGEMA_signal_18338, mcs1_mcs_mat1_3_n75}), .c ({temp_next_s3[114], temp_next_s2[114], temp_next_s1[114], temp_next_s0[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U17 ( .a ({new_AGEMA_signal_17680, new_AGEMA_signal_17679, new_AGEMA_signal_17678, mcs1_mcs_mat1_3_mcs_out[58]}), .b ({new_AGEMA_signal_13453, new_AGEMA_signal_13452, new_AGEMA_signal_13451, mcs1_mcs_mat1_3_mcs_out[62]}), .c ({new_AGEMA_signal_18340, new_AGEMA_signal_18339, new_AGEMA_signal_18338, mcs1_mcs_mat1_3_n75}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U16 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_16117, new_AGEMA_signal_16116, new_AGEMA_signal_16115, mcs1_mcs_mat1_3_mcs_out[54]}), .c ({new_AGEMA_signal_16945, new_AGEMA_signal_16944, new_AGEMA_signal_16943, mcs1_mcs_mat1_3_n76}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U15 ( .a ({new_AGEMA_signal_16948, new_AGEMA_signal_16947, new_AGEMA_signal_16946, mcs1_mcs_mat1_3_n74}), .b ({new_AGEMA_signal_18991, new_AGEMA_signal_18990, new_AGEMA_signal_18989, mcs1_mcs_mat1_3_n73}), .c ({temp_next_s3[113], temp_next_s2[113], temp_next_s1[113], temp_next_s0[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U14 ( .a ({new_AGEMA_signal_18364, new_AGEMA_signal_18363, new_AGEMA_signal_18362, mcs1_mcs_mat1_3_mcs_out[57]}), .b ({new_AGEMA_signal_13456, new_AGEMA_signal_13455, new_AGEMA_signal_13454, mcs1_mcs_mat1_3_mcs_out[61]}), .c ({new_AGEMA_signal_18991, new_AGEMA_signal_18990, new_AGEMA_signal_18989, mcs1_mcs_mat1_3_n73}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U13 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({new_AGEMA_signal_16120, new_AGEMA_signal_16119, new_AGEMA_signal_16118, mcs1_mcs_mat1_3_mcs_out[53]}), .c ({new_AGEMA_signal_16948, new_AGEMA_signal_16947, new_AGEMA_signal_16946, mcs1_mcs_mat1_3_n74}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U12 ( .a ({new_AGEMA_signal_16066, new_AGEMA_signal_16065, new_AGEMA_signal_16064, mcs1_mcs_mat1_3_n72}), .b ({new_AGEMA_signal_19729, new_AGEMA_signal_19728, new_AGEMA_signal_19727, mcs1_mcs_mat1_3_n71}), .c ({temp_next_s3[112], temp_next_s2[112], temp_next_s1[112], temp_next_s0[112]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U11 ( .a ({new_AGEMA_signal_19021, new_AGEMA_signal_19020, new_AGEMA_signal_19019, mcs1_mcs_mat1_3_mcs_out[56]}), .b ({new_AGEMA_signal_16114, new_AGEMA_signal_16113, new_AGEMA_signal_16112, mcs1_mcs_mat1_3_mcs_out[60]}), .c ({new_AGEMA_signal_19729, new_AGEMA_signal_19728, new_AGEMA_signal_19727, mcs1_mcs_mat1_3_n71}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U10 ( .a ({new_AGEMA_signal_13471, new_AGEMA_signal_13470, new_AGEMA_signal_13469, mcs1_mcs_mat1_3_mcs_out[48]}), .b ({new_AGEMA_signal_14920, new_AGEMA_signal_14919, new_AGEMA_signal_14918, mcs1_mcs_mat1_3_mcs_out[52]}), .c ({new_AGEMA_signal_16066, new_AGEMA_signal_16065, new_AGEMA_signal_16064, mcs1_mcs_mat1_3_n72}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U9 ( .a ({new_AGEMA_signal_16951, new_AGEMA_signal_16950, new_AGEMA_signal_16949, mcs1_mcs_mat1_3_n70}), .b ({new_AGEMA_signal_19732, new_AGEMA_signal_19731, new_AGEMA_signal_19730, mcs1_mcs_mat1_3_n69}), .c ({temp_next_s3[83], temp_next_s2[83], temp_next_s1[83], temp_next_s0[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U8 ( .a ({new_AGEMA_signal_19024, new_AGEMA_signal_19023, new_AGEMA_signal_19022, mcs1_mcs_mat1_3_mcs_out[43]}), .b ({new_AGEMA_signal_14923, new_AGEMA_signal_14922, new_AGEMA_signal_14921, mcs1_mcs_mat1_3_mcs_out[47]}), .c ({new_AGEMA_signal_19732, new_AGEMA_signal_19731, new_AGEMA_signal_19730, mcs1_mcs_mat1_3_n69}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U7 ( .a ({new_AGEMA_signal_14932, new_AGEMA_signal_14931, new_AGEMA_signal_14930, mcs1_mcs_mat1_3_mcs_out[35]}), .b ({new_AGEMA_signal_16126, new_AGEMA_signal_16125, new_AGEMA_signal_16124, mcs1_mcs_mat1_3_mcs_out[39]}), .c ({new_AGEMA_signal_16951, new_AGEMA_signal_16950, new_AGEMA_signal_16949, mcs1_mcs_mat1_3_n70}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U6 ( .a ({new_AGEMA_signal_14821, new_AGEMA_signal_14820, new_AGEMA_signal_14819, mcs1_mcs_mat1_3_n68}), .b ({new_AGEMA_signal_19735, new_AGEMA_signal_19734, new_AGEMA_signal_19733, mcs1_mcs_mat1_3_n67}), .c ({temp_next_s3[82], temp_next_s2[82], temp_next_s1[82], temp_next_s0[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U5 ( .a ({new_AGEMA_signal_19027, new_AGEMA_signal_19026, new_AGEMA_signal_19025, mcs1_mcs_mat1_3_mcs_out[42]}), .b ({new_AGEMA_signal_10870, new_AGEMA_signal_10869, new_AGEMA_signal_10868, mcs1_mcs_mat1_3_mcs_out[46]}), .c ({new_AGEMA_signal_19735, new_AGEMA_signal_19734, new_AGEMA_signal_19733, mcs1_mcs_mat1_3_n67}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U4 ( .a ({new_AGEMA_signal_13486, new_AGEMA_signal_13485, new_AGEMA_signal_13484, mcs1_mcs_mat1_3_mcs_out[34]}), .b ({new_AGEMA_signal_12040, new_AGEMA_signal_12039, new_AGEMA_signal_12038, mcs1_mcs_mat1_3_mcs_out[38]}), .c ({new_AGEMA_signal_14821, new_AGEMA_signal_14820, new_AGEMA_signal_14819, mcs1_mcs_mat1_3_n68}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U3 ( .a ({new_AGEMA_signal_17653, new_AGEMA_signal_17652, new_AGEMA_signal_17651, mcs1_mcs_mat1_3_n66}), .b ({new_AGEMA_signal_20566, new_AGEMA_signal_20565, new_AGEMA_signal_20564, mcs1_mcs_mat1_3_n65}), .c ({temp_next_s3[16], temp_next_s2[16], temp_next_s1[16], temp_next_s0[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U2 ( .a ({new_AGEMA_signal_17716, new_AGEMA_signal_17715, new_AGEMA_signal_17714, mcs1_mcs_mat1_3_mcs_out[4]}), .b ({new_AGEMA_signal_19756, new_AGEMA_signal_19755, new_AGEMA_signal_19754, mcs1_mcs_mat1_3_mcs_out[8]}), .c ({new_AGEMA_signal_20566, new_AGEMA_signal_20565, new_AGEMA_signal_20564, mcs1_mcs_mat1_3_n65}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_U1 ( .a ({new_AGEMA_signal_14977, new_AGEMA_signal_14976, new_AGEMA_signal_14975, mcs1_mcs_mat1_3_mcs_out[0]}), .b ({new_AGEMA_signal_16999, new_AGEMA_signal_16998, new_AGEMA_signal_16997, mcs1_mcs_mat1_3_mcs_out[12]}), .c ({new_AGEMA_signal_17653, new_AGEMA_signal_17652, new_AGEMA_signal_17651, mcs1_mcs_mat1_3_n66}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_18994, new_AGEMA_signal_18993, new_AGEMA_signal_18992, mcs1_mcs_mat1_3_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_19738, new_AGEMA_signal_19737, new_AGEMA_signal_19736, mcs1_mcs_mat1_3_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_18343, new_AGEMA_signal_18342, new_AGEMA_signal_18341, mcs1_mcs_mat1_3_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_13381, new_AGEMA_signal_13380, new_AGEMA_signal_13379, mcs1_mcs_mat1_3_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_18994, new_AGEMA_signal_18993, new_AGEMA_signal_18992, mcs1_mcs_mat1_3_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_14824, new_AGEMA_signal_14823, new_AGEMA_signal_14822, mcs1_mcs_mat1_3_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_16954, new_AGEMA_signal_16953, new_AGEMA_signal_16952, mcs1_mcs_mat1_3_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_17656, new_AGEMA_signal_17655, new_AGEMA_signal_17654, mcs1_mcs_mat1_3_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_14827, new_AGEMA_signal_14826, new_AGEMA_signal_14825, mcs1_mcs_mat1_3_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .c ({new_AGEMA_signal_16954, new_AGEMA_signal_16953, new_AGEMA_signal_16952, mcs1_mcs_mat1_3_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_18997, new_AGEMA_signal_18996, new_AGEMA_signal_18995, mcs1_mcs_mat1_3_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .c ({new_AGEMA_signal_19741, new_AGEMA_signal_19740, new_AGEMA_signal_19739, mcs1_mcs_mat1_3_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_18343, new_AGEMA_signal_18342, new_AGEMA_signal_18341, mcs1_mcs_mat1_3_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_18997, new_AGEMA_signal_18996, new_AGEMA_signal_18995, mcs1_mcs_mat1_3_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_17659, new_AGEMA_signal_17658, new_AGEMA_signal_17657, mcs1_mcs_mat1_3_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_16957, new_AGEMA_signal_16956, new_AGEMA_signal_16955, mcs1_mcs_mat1_3_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_18343, new_AGEMA_signal_18342, new_AGEMA_signal_18341, mcs1_mcs_mat1_3_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_18346, new_AGEMA_signal_18345, new_AGEMA_signal_18344, mcs1_mcs_mat1_3_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_19000, new_AGEMA_signal_18999, new_AGEMA_signal_18998, mcs1_mcs_mat1_3_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_17659, new_AGEMA_signal_17658, new_AGEMA_signal_17657, mcs1_mcs_mat1_3_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_14827, new_AGEMA_signal_14826, new_AGEMA_signal_14825, mcs1_mcs_mat1_3_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_18346, new_AGEMA_signal_18345, new_AGEMA_signal_18344, mcs1_mcs_mat1_3_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200]}), .c ({new_AGEMA_signal_17659, new_AGEMA_signal_17658, new_AGEMA_signal_17657, mcs1_mcs_mat1_3_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4211], Fresh[4210], Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206]}), .c ({new_AGEMA_signal_14827, new_AGEMA_signal_14826, new_AGEMA_signal_14825, mcs1_mcs_mat1_3_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212]}), .c ({new_AGEMA_signal_16957, new_AGEMA_signal_16956, new_AGEMA_signal_16955, mcs1_mcs_mat1_3_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_14830, new_AGEMA_signal_14829, new_AGEMA_signal_14828, mcs1_mcs_mat1_3_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .c ({new_AGEMA_signal_16069, new_AGEMA_signal_16068, new_AGEMA_signal_16067, mcs1_mcs_mat1_3_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_13384, new_AGEMA_signal_13383, new_AGEMA_signal_13382, mcs1_mcs_mat1_3_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10816, new_AGEMA_signal_10815, new_AGEMA_signal_10814, mcs1_mcs_mat1_3_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_14830, new_AGEMA_signal_14829, new_AGEMA_signal_14828, mcs1_mcs_mat1_3_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_14833, new_AGEMA_signal_14832, new_AGEMA_signal_14831, mcs1_mcs_mat1_3_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_11932, new_AGEMA_signal_11931, new_AGEMA_signal_11930, mcs1_mcs_mat1_3_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_16072, new_AGEMA_signal_16071, new_AGEMA_signal_16070, mcs1_mcs_mat1_3_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_13384, new_AGEMA_signal_13383, new_AGEMA_signal_13382, mcs1_mcs_mat1_3_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .c ({new_AGEMA_signal_14833, new_AGEMA_signal_14832, new_AGEMA_signal_14831, mcs1_mcs_mat1_3_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_13384, new_AGEMA_signal_13383, new_AGEMA_signal_13382, mcs1_mcs_mat1_3_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_11929, new_AGEMA_signal_11928, new_AGEMA_signal_11927, mcs1_mcs_mat1_3_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_14836, new_AGEMA_signal_14835, new_AGEMA_signal_14834, mcs1_mcs_mat1_3_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_11935, new_AGEMA_signal_11934, new_AGEMA_signal_11933, mcs1_mcs_mat1_3_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_9649, new_AGEMA_signal_9648, new_AGEMA_signal_9647, mcs1_mcs_mat1_3_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_13384, new_AGEMA_signal_13383, new_AGEMA_signal_13382, mcs1_mcs_mat1_3_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_10813, new_AGEMA_signal_10812, new_AGEMA_signal_10811, mcs1_mcs_mat1_3_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_11932, new_AGEMA_signal_11931, new_AGEMA_signal_11930, mcs1_mcs_mat1_3_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_13387, new_AGEMA_signal_13386, new_AGEMA_signal_13385, mcs1_mcs_mat1_3_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_8827, new_AGEMA_signal_8826, new_AGEMA_signal_8825, mcs1_mcs_mat1_3_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_10816, new_AGEMA_signal_10815, new_AGEMA_signal_10814, mcs1_mcs_mat1_3_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_11932, new_AGEMA_signal_11931, new_AGEMA_signal_11930, mcs1_mcs_mat1_3_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_9649, new_AGEMA_signal_9648, new_AGEMA_signal_9647, mcs1_mcs_mat1_3_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_10813, new_AGEMA_signal_10812, new_AGEMA_signal_10811, mcs1_mcs_mat1_3_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220], Fresh[4219], Fresh[4218]}), .c ({new_AGEMA_signal_11935, new_AGEMA_signal_11934, new_AGEMA_signal_11933, mcs1_mcs_mat1_3_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224]}), .c ({new_AGEMA_signal_9649, new_AGEMA_signal_9648, new_AGEMA_signal_9647, mcs1_mcs_mat1_3_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230]}), .c ({new_AGEMA_signal_10816, new_AGEMA_signal_10815, new_AGEMA_signal_10814, mcs1_mcs_mat1_3_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_13393, new_AGEMA_signal_13392, new_AGEMA_signal_13391, mcs1_mcs_mat1_3_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_9652, new_AGEMA_signal_9651, new_AGEMA_signal_9650, mcs1_mcs_mat1_3_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_14839, new_AGEMA_signal_14838, new_AGEMA_signal_14837, mcs1_mcs_mat1_3_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_10819, new_AGEMA_signal_10818, new_AGEMA_signal_10817, mcs1_mcs_mat1_3_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_10822, new_AGEMA_signal_10821, new_AGEMA_signal_10820, mcs1_mcs_mat1_3_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_11938, new_AGEMA_signal_11937, new_AGEMA_signal_11936, mcs1_mcs_mat1_3_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_13396, new_AGEMA_signal_13395, new_AGEMA_signal_13394, mcs1_mcs_mat1_3_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_14842, new_AGEMA_signal_14841, new_AGEMA_signal_14840, mcs1_mcs_mat1_3_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_16075, new_AGEMA_signal_16074, new_AGEMA_signal_16073, mcs1_mcs_mat1_3_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_13393, new_AGEMA_signal_13392, new_AGEMA_signal_13391, mcs1_mcs_mat1_3_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_14842, new_AGEMA_signal_14841, new_AGEMA_signal_14840, mcs1_mcs_mat1_3_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_8830, new_AGEMA_signal_8829, new_AGEMA_signal_8828, mcs1_mcs_mat1_3_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_11944, new_AGEMA_signal_11943, new_AGEMA_signal_11942, mcs1_mcs_mat1_3_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_13393, new_AGEMA_signal_13392, new_AGEMA_signal_13391, mcs1_mcs_mat1_3_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_9655, new_AGEMA_signal_9654, new_AGEMA_signal_9653, mcs1_mcs_mat1_3_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_11941, new_AGEMA_signal_11940, new_AGEMA_signal_11939, mcs1_mcs_mat1_3_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_13396, new_AGEMA_signal_13395, new_AGEMA_signal_13394, mcs1_mcs_mat1_3_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4241], Fresh[4240], Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236]}), .c ({new_AGEMA_signal_11944, new_AGEMA_signal_11943, new_AGEMA_signal_11942, mcs1_mcs_mat1_3_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242]}), .c ({new_AGEMA_signal_9655, new_AGEMA_signal_9654, new_AGEMA_signal_9653, mcs1_mcs_mat1_3_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250], Fresh[4249], Fresh[4248]}), .c ({new_AGEMA_signal_10822, new_AGEMA_signal_10821, new_AGEMA_signal_10820, mcs1_mcs_mat1_3_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({new_AGEMA_signal_14845, new_AGEMA_signal_14844, new_AGEMA_signal_14843, mcs1_mcs_mat1_3_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_16078, new_AGEMA_signal_16077, new_AGEMA_signal_16076, mcs1_mcs_mat1_3_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({new_AGEMA_signal_14848, new_AGEMA_signal_14847, new_AGEMA_signal_14846, mcs1_mcs_mat1_3_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_16081, new_AGEMA_signal_16080, new_AGEMA_signal_16079, mcs1_mcs_mat1_3_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_10825, new_AGEMA_signal_10824, new_AGEMA_signal_10823, mcs1_mcs_mat1_3_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_14845, new_AGEMA_signal_14844, new_AGEMA_signal_14843, mcs1_mcs_mat1_3_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_16084, new_AGEMA_signal_16083, new_AGEMA_signal_16082, mcs1_mcs_mat1_3_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_9658, new_AGEMA_signal_9657, new_AGEMA_signal_9656, mcs1_mcs_mat1_3_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_13399, new_AGEMA_signal_13398, new_AGEMA_signal_13397, mcs1_mcs_mat1_3_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_14845, new_AGEMA_signal_14844, new_AGEMA_signal_14843, mcs1_mcs_mat1_3_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_11947, new_AGEMA_signal_11946, new_AGEMA_signal_11945, mcs1_mcs_mat1_3_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_14848, new_AGEMA_signal_14847, new_AGEMA_signal_14846, mcs1_mcs_mat1_3_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_16087, new_AGEMA_signal_16086, new_AGEMA_signal_16085, mcs1_mcs_mat1_3_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_13402, new_AGEMA_signal_13401, new_AGEMA_signal_13400, mcs1_mcs_mat1_3_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_14848, new_AGEMA_signal_14847, new_AGEMA_signal_14846, mcs1_mcs_mat1_3_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_10825, new_AGEMA_signal_10824, new_AGEMA_signal_10823, mcs1_mcs_mat1_3_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_11950, new_AGEMA_signal_11949, new_AGEMA_signal_11948, mcs1_mcs_mat1_3_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_13402, new_AGEMA_signal_13401, new_AGEMA_signal_13400, mcs1_mcs_mat1_3_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254]}), .c ({new_AGEMA_signal_11950, new_AGEMA_signal_11949, new_AGEMA_signal_11948, mcs1_mcs_mat1_3_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260]}), .c ({new_AGEMA_signal_9658, new_AGEMA_signal_9657, new_AGEMA_signal_9656, mcs1_mcs_mat1_3_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4271], Fresh[4270], Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266]}), .c ({new_AGEMA_signal_10825, new_AGEMA_signal_10824, new_AGEMA_signal_10823, mcs1_mcs_mat1_3_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_18352, new_AGEMA_signal_18351, new_AGEMA_signal_18350, mcs1_mcs_mat1_3_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_18349, new_AGEMA_signal_18348, new_AGEMA_signal_18347, mcs1_mcs_mat1_3_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_19003, new_AGEMA_signal_19002, new_AGEMA_signal_19001, mcs1_mcs_mat1_3_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_18349, new_AGEMA_signal_18348, new_AGEMA_signal_18347, mcs1_mcs_mat1_3_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_16960, new_AGEMA_signal_16959, new_AGEMA_signal_16958, mcs1_mcs_mat1_3_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_19006, new_AGEMA_signal_19005, new_AGEMA_signal_19004, mcs1_mcs_mat1_3_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_14851, new_AGEMA_signal_14850, new_AGEMA_signal_14849, mcs1_mcs_mat1_3_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .c ({new_AGEMA_signal_16960, new_AGEMA_signal_16959, new_AGEMA_signal_16958, mcs1_mcs_mat1_3_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({new_AGEMA_signal_18349, new_AGEMA_signal_18348, new_AGEMA_signal_18347, mcs1_mcs_mat1_3_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_19009, new_AGEMA_signal_19008, new_AGEMA_signal_19007, mcs1_mcs_mat1_3_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_17665, new_AGEMA_signal_17664, new_AGEMA_signal_17663, mcs1_mcs_mat1_3_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_13405, new_AGEMA_signal_13404, new_AGEMA_signal_13403, mcs1_mcs_mat1_3_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_18349, new_AGEMA_signal_18348, new_AGEMA_signal_18347, mcs1_mcs_mat1_3_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_19012, new_AGEMA_signal_19011, new_AGEMA_signal_19010, mcs1_mcs_mat1_3_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_19744, new_AGEMA_signal_19743, new_AGEMA_signal_19742, mcs1_mcs_mat1_3_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_18352, new_AGEMA_signal_18351, new_AGEMA_signal_18350, mcs1_mcs_mat1_3_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_17665, new_AGEMA_signal_17664, new_AGEMA_signal_17663, mcs1_mcs_mat1_3_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_19012, new_AGEMA_signal_19011, new_AGEMA_signal_19010, mcs1_mcs_mat1_3_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_17662, new_AGEMA_signal_17661, new_AGEMA_signal_17660, mcs1_mcs_mat1_3_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .c ({new_AGEMA_signal_18352, new_AGEMA_signal_18351, new_AGEMA_signal_18350, mcs1_mcs_mat1_3_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_14851, new_AGEMA_signal_14850, new_AGEMA_signal_14849, mcs1_mcs_mat1_3_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_16963, new_AGEMA_signal_16962, new_AGEMA_signal_16961, mcs1_mcs_mat1_3_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_17662, new_AGEMA_signal_17661, new_AGEMA_signal_17660, mcs1_mcs_mat1_3_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272]}), .c ({new_AGEMA_signal_17665, new_AGEMA_signal_17664, new_AGEMA_signal_17663, mcs1_mcs_mat1_3_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280], Fresh[4279], Fresh[4278]}), .c ({new_AGEMA_signal_14851, new_AGEMA_signal_14850, new_AGEMA_signal_14849, mcs1_mcs_mat1_3_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284]}), .c ({new_AGEMA_signal_16963, new_AGEMA_signal_16962, new_AGEMA_signal_16961, mcs1_mcs_mat1_3_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_10828, new_AGEMA_signal_10827, new_AGEMA_signal_10826, mcs1_mcs_mat1_3_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_13408, new_AGEMA_signal_13407, new_AGEMA_signal_13406, mcs1_mcs_mat1_3_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_14854, new_AGEMA_signal_14853, new_AGEMA_signal_14852, mcs1_mcs_mat1_3_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_11962, new_AGEMA_signal_11961, new_AGEMA_signal_11960, mcs1_mcs_mat1_3_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_13408, new_AGEMA_signal_13407, new_AGEMA_signal_13406, mcs1_mcs_mat1_3_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_11956, new_AGEMA_signal_11955, new_AGEMA_signal_11954, mcs1_mcs_mat1_3_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_10831, new_AGEMA_signal_10830, new_AGEMA_signal_10829, mcs1_mcs_mat1_3_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_13411, new_AGEMA_signal_13410, new_AGEMA_signal_13409, mcs1_mcs_mat1_3_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_11959, new_AGEMA_signal_11958, new_AGEMA_signal_11957, mcs1_mcs_mat1_3_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_13414, new_AGEMA_signal_13413, new_AGEMA_signal_13412, mcs1_mcs_mat1_3_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_14857, new_AGEMA_signal_14856, new_AGEMA_signal_14855, mcs1_mcs_mat1_3_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_8836, new_AGEMA_signal_8835, new_AGEMA_signal_8834, mcs1_mcs_mat1_3_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_11962, new_AGEMA_signal_11961, new_AGEMA_signal_11960, mcs1_mcs_mat1_3_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_13414, new_AGEMA_signal_13413, new_AGEMA_signal_13412, mcs1_mcs_mat1_3_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_9661, new_AGEMA_signal_9660, new_AGEMA_signal_9659, mcs1_mcs_mat1_3_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .c ({new_AGEMA_signal_11959, new_AGEMA_signal_11958, new_AGEMA_signal_11957, mcs1_mcs_mat1_3_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290]}), .c ({new_AGEMA_signal_11962, new_AGEMA_signal_11961, new_AGEMA_signal_11960, mcs1_mcs_mat1_3_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4301], Fresh[4300], Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296]}), .c ({new_AGEMA_signal_9661, new_AGEMA_signal_9660, new_AGEMA_signal_9659, mcs1_mcs_mat1_3_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4307], Fresh[4306], Fresh[4305], Fresh[4304], Fresh[4303], Fresh[4302]}), .c ({new_AGEMA_signal_10831, new_AGEMA_signal_10830, new_AGEMA_signal_10829, mcs1_mcs_mat1_3_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_16966, new_AGEMA_signal_16965, new_AGEMA_signal_16964, mcs1_mcs_mat1_3_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_10837, new_AGEMA_signal_10836, new_AGEMA_signal_10835, mcs1_mcs_mat1_3_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_17668, new_AGEMA_signal_17667, new_AGEMA_signal_17666, mcs1_mcs_mat1_3_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_16090, new_AGEMA_signal_16089, new_AGEMA_signal_16088, mcs1_mcs_mat1_3_mcs_out[99]}), .b ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .c ({new_AGEMA_signal_16966, new_AGEMA_signal_16965, new_AGEMA_signal_16964, mcs1_mcs_mat1_3_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_14860, new_AGEMA_signal_14859, new_AGEMA_signal_14858, mcs1_mcs_mat1_3_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .c ({new_AGEMA_signal_16090, new_AGEMA_signal_16089, new_AGEMA_signal_16088, mcs1_mcs_mat1_3_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_13417, new_AGEMA_signal_13416, new_AGEMA_signal_13415, mcs1_mcs_mat1_3_mcs_out[98]}), .b ({new_AGEMA_signal_9667, new_AGEMA_signal_9666, new_AGEMA_signal_9665, mcs1_mcs_mat1_3_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_14860, new_AGEMA_signal_14859, new_AGEMA_signal_14858, mcs1_mcs_mat1_3_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_9664, new_AGEMA_signal_9663, new_AGEMA_signal_9662, mcs1_mcs_mat1_3_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_11965, new_AGEMA_signal_11964, new_AGEMA_signal_11963, mcs1_mcs_mat1_3_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_13417, new_AGEMA_signal_13416, new_AGEMA_signal_13415, mcs1_mcs_mat1_3_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310], Fresh[4309], Fresh[4308]}), .c ({new_AGEMA_signal_11965, new_AGEMA_signal_11964, new_AGEMA_signal_11963, mcs1_mcs_mat1_3_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314]}), .c ({new_AGEMA_signal_9667, new_AGEMA_signal_9666, new_AGEMA_signal_9665, mcs1_mcs_mat1_3_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320]}), .c ({new_AGEMA_signal_10837, new_AGEMA_signal_10836, new_AGEMA_signal_10835, mcs1_mcs_mat1_3_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_13420, new_AGEMA_signal_13419, new_AGEMA_signal_13418, mcs1_mcs_mat1_3_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_14863, new_AGEMA_signal_14862, new_AGEMA_signal_14861, mcs1_mcs_mat1_3_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_10843, new_AGEMA_signal_10842, new_AGEMA_signal_10841, mcs1_mcs_mat1_3_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_10846, new_AGEMA_signal_10845, new_AGEMA_signal_10844, mcs1_mcs_mat1_3_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_11971, new_AGEMA_signal_11970, new_AGEMA_signal_11969, mcs1_mcs_mat1_3_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_14866, new_AGEMA_signal_14865, new_AGEMA_signal_14864, mcs1_mcs_mat1_3_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_9670, new_AGEMA_signal_9669, new_AGEMA_signal_9668, mcs1_mcs_mat1_3_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_16093, new_AGEMA_signal_16092, new_AGEMA_signal_16091, mcs1_mcs_mat1_3_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_13420, new_AGEMA_signal_13419, new_AGEMA_signal_13418, mcs1_mcs_mat1_3_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .c ({new_AGEMA_signal_14866, new_AGEMA_signal_14865, new_AGEMA_signal_14864, mcs1_mcs_mat1_3_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_8842, new_AGEMA_signal_8841, new_AGEMA_signal_8840, mcs1_mcs_mat1_3_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_11974, new_AGEMA_signal_11973, new_AGEMA_signal_11972, mcs1_mcs_mat1_3_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_13420, new_AGEMA_signal_13419, new_AGEMA_signal_13418, mcs1_mcs_mat1_3_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4331], Fresh[4330], Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326]}), .c ({new_AGEMA_signal_11974, new_AGEMA_signal_11973, new_AGEMA_signal_11972, mcs1_mcs_mat1_3_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4337], Fresh[4336], Fresh[4335], Fresh[4334], Fresh[4333], Fresh[4332]}), .c ({new_AGEMA_signal_9670, new_AGEMA_signal_9669, new_AGEMA_signal_9668, mcs1_mcs_mat1_3_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340], Fresh[4339], Fresh[4338]}), .c ({new_AGEMA_signal_10846, new_AGEMA_signal_10845, new_AGEMA_signal_10844, mcs1_mcs_mat1_3_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_11986, new_AGEMA_signal_11985, new_AGEMA_signal_11984, mcs1_mcs_mat1_3_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_11989, new_AGEMA_signal_11988, new_AGEMA_signal_11987, mcs1_mcs_mat1_3_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_13426, new_AGEMA_signal_13425, new_AGEMA_signal_13424, mcs1_mcs_mat1_3_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_11980, new_AGEMA_signal_11979, new_AGEMA_signal_11978, mcs1_mcs_mat1_3_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_8845, new_AGEMA_signal_8844, new_AGEMA_signal_8843, mcs1_mcs_mat1_3_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_13429, new_AGEMA_signal_13428, new_AGEMA_signal_13427, mcs1_mcs_mat1_3_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_10849, new_AGEMA_signal_10848, new_AGEMA_signal_10847, mcs1_mcs_mat1_3_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_11980, new_AGEMA_signal_11979, new_AGEMA_signal_11978, mcs1_mcs_mat1_3_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_11983, new_AGEMA_signal_11982, new_AGEMA_signal_11981, mcs1_mcs_mat1_3_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_13432, new_AGEMA_signal_13431, new_AGEMA_signal_13430, mcs1_mcs_mat1_3_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_9673, new_AGEMA_signal_9672, new_AGEMA_signal_9671, mcs1_mcs_mat1_3_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_10849, new_AGEMA_signal_10848, new_AGEMA_signal_10847, mcs1_mcs_mat1_3_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_11983, new_AGEMA_signal_11982, new_AGEMA_signal_11981, mcs1_mcs_mat1_3_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_13435, new_AGEMA_signal_13434, new_AGEMA_signal_13433, mcs1_mcs_mat1_3_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .c ({new_AGEMA_signal_14869, new_AGEMA_signal_14868, new_AGEMA_signal_14867, mcs1_mcs_mat1_3_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_11986, new_AGEMA_signal_11985, new_AGEMA_signal_11984, mcs1_mcs_mat1_3_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_9673, new_AGEMA_signal_9672, new_AGEMA_signal_9671, mcs1_mcs_mat1_3_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_13435, new_AGEMA_signal_13434, new_AGEMA_signal_13433, mcs1_mcs_mat1_3_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344]}), .c ({new_AGEMA_signal_11989, new_AGEMA_signal_11988, new_AGEMA_signal_11987, mcs1_mcs_mat1_3_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350]}), .c ({new_AGEMA_signal_9673, new_AGEMA_signal_9672, new_AGEMA_signal_9671, mcs1_mcs_mat1_3_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4361], Fresh[4360], Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356]}), .c ({new_AGEMA_signal_10849, new_AGEMA_signal_10848, new_AGEMA_signal_10847, mcs1_mcs_mat1_3_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_13438, new_AGEMA_signal_13437, new_AGEMA_signal_13436, mcs1_mcs_mat1_3_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_14872, new_AGEMA_signal_14871, new_AGEMA_signal_14870, mcs1_mcs_mat1_3_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_10852, new_AGEMA_signal_10851, new_AGEMA_signal_10850, mcs1_mcs_mat1_3_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_11992, new_AGEMA_signal_11991, new_AGEMA_signal_11990, mcs1_mcs_mat1_3_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_14875, new_AGEMA_signal_14874, new_AGEMA_signal_14873, mcs1_mcs_mat1_3_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_9679, new_AGEMA_signal_9678, new_AGEMA_signal_9677, mcs1_mcs_mat1_3_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_16096, new_AGEMA_signal_16095, new_AGEMA_signal_16094, mcs1_mcs_mat1_3_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_13438, new_AGEMA_signal_13437, new_AGEMA_signal_13436, mcs1_mcs_mat1_3_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .c ({new_AGEMA_signal_14875, new_AGEMA_signal_14874, new_AGEMA_signal_14873, mcs1_mcs_mat1_3_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_8848, new_AGEMA_signal_8847, new_AGEMA_signal_8846, mcs1_mcs_mat1_3_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_11995, new_AGEMA_signal_11994, new_AGEMA_signal_11993, mcs1_mcs_mat1_3_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_13438, new_AGEMA_signal_13437, new_AGEMA_signal_13436, mcs1_mcs_mat1_3_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4367], Fresh[4366], Fresh[4365], Fresh[4364], Fresh[4363], Fresh[4362]}), .c ({new_AGEMA_signal_11995, new_AGEMA_signal_11994, new_AGEMA_signal_11993, mcs1_mcs_mat1_3_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370], Fresh[4369], Fresh[4368]}), .c ({new_AGEMA_signal_9679, new_AGEMA_signal_9678, new_AGEMA_signal_9677, mcs1_mcs_mat1_3_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374]}), .c ({new_AGEMA_signal_10852, new_AGEMA_signal_10851, new_AGEMA_signal_10850, mcs1_mcs_mat1_3_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_19015, new_AGEMA_signal_19014, new_AGEMA_signal_19013, mcs1_mcs_mat1_3_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_19747, new_AGEMA_signal_19746, new_AGEMA_signal_19745, mcs1_mcs_mat1_3_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_18358, new_AGEMA_signal_18357, new_AGEMA_signal_18356, mcs1_mcs_mat1_3_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_17674, new_AGEMA_signal_17673, new_AGEMA_signal_17672, mcs1_mcs_mat1_3_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_19015, new_AGEMA_signal_19014, new_AGEMA_signal_19013, mcs1_mcs_mat1_3_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({new_AGEMA_signal_16099, new_AGEMA_signal_16098, new_AGEMA_signal_16097, mcs1_mcs_mat1_3_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_17671, new_AGEMA_signal_17670, new_AGEMA_signal_17669, mcs1_mcs_mat1_3_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_17674, new_AGEMA_signal_17673, new_AGEMA_signal_17672, mcs1_mcs_mat1_3_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_16099, new_AGEMA_signal_16098, new_AGEMA_signal_16097, mcs1_mcs_mat1_3_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_18355, new_AGEMA_signal_18354, new_AGEMA_signal_18353, mcs1_mcs_mat1_3_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_14878, new_AGEMA_signal_14877, new_AGEMA_signal_14876, mcs1_mcs_mat1_3_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_14881, new_AGEMA_signal_14880, new_AGEMA_signal_14879, mcs1_mcs_mat1_3_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_16099, new_AGEMA_signal_16098, new_AGEMA_signal_16097, mcs1_mcs_mat1_3_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_16975, new_AGEMA_signal_16974, new_AGEMA_signal_16973, mcs1_mcs_mat1_3_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .c ({new_AGEMA_signal_17674, new_AGEMA_signal_17673, new_AGEMA_signal_17672, mcs1_mcs_mat1_3_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_19018, new_AGEMA_signal_19017, new_AGEMA_signal_19016, mcs1_mcs_mat1_3_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_14878, new_AGEMA_signal_14877, new_AGEMA_signal_14876, mcs1_mcs_mat1_3_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_19750, new_AGEMA_signal_19749, new_AGEMA_signal_19748, mcs1_mcs_mat1_3_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_18358, new_AGEMA_signal_18357, new_AGEMA_signal_18356, mcs1_mcs_mat1_3_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_16975, new_AGEMA_signal_16974, new_AGEMA_signal_16973, mcs1_mcs_mat1_3_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_19018, new_AGEMA_signal_19017, new_AGEMA_signal_19016, mcs1_mcs_mat1_3_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .b ({new_AGEMA_signal_17677, new_AGEMA_signal_17676, new_AGEMA_signal_17675, mcs1_mcs_mat1_3_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_18358, new_AGEMA_signal_18357, new_AGEMA_signal_18356, mcs1_mcs_mat1_3_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380]}), .c ({new_AGEMA_signal_17677, new_AGEMA_signal_17676, new_AGEMA_signal_17675, mcs1_mcs_mat1_3_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4391], Fresh[4390], Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386]}), .c ({new_AGEMA_signal_14881, new_AGEMA_signal_14880, new_AGEMA_signal_14879, mcs1_mcs_mat1_3_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4397], Fresh[4396], Fresh[4395], Fresh[4394], Fresh[4393], Fresh[4392]}), .c ({new_AGEMA_signal_16975, new_AGEMA_signal_16974, new_AGEMA_signal_16973, mcs1_mcs_mat1_3_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_13444, new_AGEMA_signal_13443, new_AGEMA_signal_13442, mcs1_mcs_mat1_3_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_10855, new_AGEMA_signal_10854, new_AGEMA_signal_10853, mcs1_mcs_mat1_3_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_14884, new_AGEMA_signal_14883, new_AGEMA_signal_14882, mcs1_mcs_mat1_3_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_12001, new_AGEMA_signal_12000, new_AGEMA_signal_11999, mcs1_mcs_mat1_3_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_14887, new_AGEMA_signal_14886, new_AGEMA_signal_14885, mcs1_mcs_mat1_3_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_16102, new_AGEMA_signal_16101, new_AGEMA_signal_16100, mcs1_mcs_mat1_3_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_13444, new_AGEMA_signal_13443, new_AGEMA_signal_13442, mcs1_mcs_mat1_3_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_14887, new_AGEMA_signal_14886, new_AGEMA_signal_14885, mcs1_mcs_mat1_3_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_16105, new_AGEMA_signal_16104, new_AGEMA_signal_16103, mcs1_mcs_mat1_3_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_10855, new_AGEMA_signal_10854, new_AGEMA_signal_10853, mcs1_mcs_mat1_3_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_13447, new_AGEMA_signal_13446, new_AGEMA_signal_13445, mcs1_mcs_mat1_3_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_14887, new_AGEMA_signal_14886, new_AGEMA_signal_14885, mcs1_mcs_mat1_3_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({new_AGEMA_signal_9682, new_AGEMA_signal_9681, new_AGEMA_signal_9680, mcs1_mcs_mat1_3_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_10855, new_AGEMA_signal_10854, new_AGEMA_signal_10853, mcs1_mcs_mat1_3_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_11998, new_AGEMA_signal_11997, new_AGEMA_signal_11996, mcs1_mcs_mat1_3_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .c ({new_AGEMA_signal_13444, new_AGEMA_signal_13443, new_AGEMA_signal_13442, mcs1_mcs_mat1_3_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_10858, new_AGEMA_signal_10857, new_AGEMA_signal_10856, mcs1_mcs_mat1_3_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8851, new_AGEMA_signal_8850, new_AGEMA_signal_8849, mcs1_mcs_mat1_3_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_11998, new_AGEMA_signal_11997, new_AGEMA_signal_11996, mcs1_mcs_mat1_3_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_13447, new_AGEMA_signal_13446, new_AGEMA_signal_13445, mcs1_mcs_mat1_3_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_12001, new_AGEMA_signal_12000, new_AGEMA_signal_11999, mcs1_mcs_mat1_3_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_14890, new_AGEMA_signal_14889, new_AGEMA_signal_14888, mcs1_mcs_mat1_3_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_10858, new_AGEMA_signal_10857, new_AGEMA_signal_10856, mcs1_mcs_mat1_3_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_12001, new_AGEMA_signal_12000, new_AGEMA_signal_11999, mcs1_mcs_mat1_3_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({new_AGEMA_signal_12004, new_AGEMA_signal_12003, new_AGEMA_signal_12002, mcs1_mcs_mat1_3_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_13447, new_AGEMA_signal_13446, new_AGEMA_signal_13445, mcs1_mcs_mat1_3_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400], Fresh[4399], Fresh[4398]}), .c ({new_AGEMA_signal_12004, new_AGEMA_signal_12003, new_AGEMA_signal_12002, mcs1_mcs_mat1_3_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404]}), .c ({new_AGEMA_signal_9682, new_AGEMA_signal_9681, new_AGEMA_signal_9680, mcs1_mcs_mat1_3_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410]}), .c ({new_AGEMA_signal_10858, new_AGEMA_signal_10857, new_AGEMA_signal_10856, mcs1_mcs_mat1_3_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_14896, new_AGEMA_signal_14895, new_AGEMA_signal_14894, mcs1_mcs_mat1_3_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .c ({new_AGEMA_signal_16108, new_AGEMA_signal_16107, new_AGEMA_signal_16106, mcs1_mcs_mat1_3_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({new_AGEMA_signal_13450, new_AGEMA_signal_13449, new_AGEMA_signal_13448, mcs1_mcs_mat1_3_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_14893, new_AGEMA_signal_14892, new_AGEMA_signal_14891, mcs1_mcs_mat1_3_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_16111, new_AGEMA_signal_16110, new_AGEMA_signal_16109, mcs1_mcs_mat1_3_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_10861, new_AGEMA_signal_10860, new_AGEMA_signal_10859, mcs1_mcs_mat1_3_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_16978, new_AGEMA_signal_16977, new_AGEMA_signal_16976, mcs1_mcs_mat1_3_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_14896, new_AGEMA_signal_14895, new_AGEMA_signal_14894, mcs1_mcs_mat1_3_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .c ({new_AGEMA_signal_16111, new_AGEMA_signal_16110, new_AGEMA_signal_16109, mcs1_mcs_mat1_3_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_9685, new_AGEMA_signal_9684, new_AGEMA_signal_9683, mcs1_mcs_mat1_3_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_13450, new_AGEMA_signal_13449, new_AGEMA_signal_13448, mcs1_mcs_mat1_3_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_14896, new_AGEMA_signal_14895, new_AGEMA_signal_14894, mcs1_mcs_mat1_3_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_8854, new_AGEMA_signal_8853, new_AGEMA_signal_8852, mcs1_mcs_mat1_3_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_12010, new_AGEMA_signal_12009, new_AGEMA_signal_12008, mcs1_mcs_mat1_3_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_13450, new_AGEMA_signal_13449, new_AGEMA_signal_13448, mcs1_mcs_mat1_3_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4421], Fresh[4420], Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416]}), .c ({new_AGEMA_signal_12010, new_AGEMA_signal_12009, new_AGEMA_signal_12008, mcs1_mcs_mat1_3_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4427], Fresh[4426], Fresh[4425], Fresh[4424], Fresh[4423], Fresh[4422]}), .c ({new_AGEMA_signal_9685, new_AGEMA_signal_9684, new_AGEMA_signal_9683, mcs1_mcs_mat1_3_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430], Fresh[4429], Fresh[4428]}), .c ({new_AGEMA_signal_10861, new_AGEMA_signal_10860, new_AGEMA_signal_10859, mcs1_mcs_mat1_3_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_13459, new_AGEMA_signal_13458, new_AGEMA_signal_13457, mcs1_mcs_mat1_3_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_10864, new_AGEMA_signal_10863, new_AGEMA_signal_10862, mcs1_mcs_mat1_3_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_14899, new_AGEMA_signal_14898, new_AGEMA_signal_14897, mcs1_mcs_mat1_3_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_9688, new_AGEMA_signal_9687, new_AGEMA_signal_9686, mcs1_mcs_mat1_3_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_12013, new_AGEMA_signal_12012, new_AGEMA_signal_12011, mcs1_mcs_mat1_3_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_13453, new_AGEMA_signal_13452, new_AGEMA_signal_13451, mcs1_mcs_mat1_3_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({new_AGEMA_signal_12016, new_AGEMA_signal_12015, new_AGEMA_signal_12014, mcs1_mcs_mat1_3_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_13456, new_AGEMA_signal_13455, new_AGEMA_signal_13454, mcs1_mcs_mat1_3_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434]}), .c ({new_AGEMA_signal_12016, new_AGEMA_signal_12015, new_AGEMA_signal_12014, mcs1_mcs_mat1_3_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440]}), .c ({new_AGEMA_signal_9688, new_AGEMA_signal_9687, new_AGEMA_signal_9686, mcs1_mcs_mat1_3_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4451], Fresh[4450], Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446]}), .c ({new_AGEMA_signal_10864, new_AGEMA_signal_10863, new_AGEMA_signal_10862, mcs1_mcs_mat1_3_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_14908, new_AGEMA_signal_14907, new_AGEMA_signal_14906, mcs1_mcs_mat1_3_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_16981, new_AGEMA_signal_16980, new_AGEMA_signal_16979, mcs1_mcs_mat1_3_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_17680, new_AGEMA_signal_17679, new_AGEMA_signal_17678, mcs1_mcs_mat1_3_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_14911, new_AGEMA_signal_14910, new_AGEMA_signal_14909, mcs1_mcs_mat1_3_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_17683, new_AGEMA_signal_17682, new_AGEMA_signal_17681, mcs1_mcs_mat1_3_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_18364, new_AGEMA_signal_18363, new_AGEMA_signal_18362, mcs1_mcs_mat1_3_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_18367, new_AGEMA_signal_18366, new_AGEMA_signal_18365, mcs1_mcs_mat1_3_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_17686, new_AGEMA_signal_17685, new_AGEMA_signal_17684, mcs1_mcs_mat1_3_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_19021, new_AGEMA_signal_19020, new_AGEMA_signal_19019, mcs1_mcs_mat1_3_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_17689, new_AGEMA_signal_17688, new_AGEMA_signal_17687, mcs1_mcs_mat1_3_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_18367, new_AGEMA_signal_18366, new_AGEMA_signal_18365, mcs1_mcs_mat1_3_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4457], Fresh[4456], Fresh[4455], Fresh[4454], Fresh[4453], Fresh[4452]}), .c ({new_AGEMA_signal_17689, new_AGEMA_signal_17688, new_AGEMA_signal_17687, mcs1_mcs_mat1_3_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460], Fresh[4459], Fresh[4458]}), .c ({new_AGEMA_signal_14911, new_AGEMA_signal_14910, new_AGEMA_signal_14909, mcs1_mcs_mat1_3_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464]}), .c ({new_AGEMA_signal_16981, new_AGEMA_signal_16980, new_AGEMA_signal_16979, mcs1_mcs_mat1_3_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_12022, new_AGEMA_signal_12021, new_AGEMA_signal_12020, mcs1_mcs_mat1_3_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_13465, new_AGEMA_signal_13464, new_AGEMA_signal_13463, mcs1_mcs_mat1_3_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_14914, new_AGEMA_signal_14913, new_AGEMA_signal_14912, mcs1_mcs_mat1_3_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_14917, new_AGEMA_signal_14916, new_AGEMA_signal_14915, mcs1_mcs_mat1_3_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_12019, new_AGEMA_signal_12018, new_AGEMA_signal_12017, mcs1_mcs_mat1_3_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_16117, new_AGEMA_signal_16116, new_AGEMA_signal_16115, mcs1_mcs_mat1_3_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_10867, new_AGEMA_signal_10866, new_AGEMA_signal_10865, mcs1_mcs_mat1_3_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_12019, new_AGEMA_signal_12018, new_AGEMA_signal_12017, mcs1_mcs_mat1_3_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({new_AGEMA_signal_14917, new_AGEMA_signal_14916, new_AGEMA_signal_14915, mcs1_mcs_mat1_3_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_16120, new_AGEMA_signal_16119, new_AGEMA_signal_16118, mcs1_mcs_mat1_3_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_8860, new_AGEMA_signal_8859, new_AGEMA_signal_8858, mcs1_mcs_mat1_3_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_13465, new_AGEMA_signal_13464, new_AGEMA_signal_13463, mcs1_mcs_mat1_3_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_14917, new_AGEMA_signal_14916, new_AGEMA_signal_14915, mcs1_mcs_mat1_3_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_9691, new_AGEMA_signal_9690, new_AGEMA_signal_9689, mcs1_mcs_mat1_3_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_12028, new_AGEMA_signal_12027, new_AGEMA_signal_12026, mcs1_mcs_mat1_3_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_13465, new_AGEMA_signal_13464, new_AGEMA_signal_13463, mcs1_mcs_mat1_3_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_12025, new_AGEMA_signal_12024, new_AGEMA_signal_12023, mcs1_mcs_mat1_3_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_13468, new_AGEMA_signal_13467, new_AGEMA_signal_13466, mcs1_mcs_mat1_3_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_14920, new_AGEMA_signal_14919, new_AGEMA_signal_14918, mcs1_mcs_mat1_3_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_12022, new_AGEMA_signal_12021, new_AGEMA_signal_12020, mcs1_mcs_mat1_3_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_9691, new_AGEMA_signal_9690, new_AGEMA_signal_9689, mcs1_mcs_mat1_3_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_13468, new_AGEMA_signal_13467, new_AGEMA_signal_13466, mcs1_mcs_mat1_3_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_10867, new_AGEMA_signal_10866, new_AGEMA_signal_10865, mcs1_mcs_mat1_3_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_12022, new_AGEMA_signal_12021, new_AGEMA_signal_12020, mcs1_mcs_mat1_3_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470]}), .c ({new_AGEMA_signal_12028, new_AGEMA_signal_12027, new_AGEMA_signal_12026, mcs1_mcs_mat1_3_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4481], Fresh[4480], Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476]}), .c ({new_AGEMA_signal_9691, new_AGEMA_signal_9690, new_AGEMA_signal_9689, mcs1_mcs_mat1_3_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4487], Fresh[4486], Fresh[4485], Fresh[4484], Fresh[4483], Fresh[4482]}), .c ({new_AGEMA_signal_10867, new_AGEMA_signal_10866, new_AGEMA_signal_10865, mcs1_mcs_mat1_3_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_10873, new_AGEMA_signal_10872, new_AGEMA_signal_10871, mcs1_mcs_mat1_3_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_12034, new_AGEMA_signal_12033, new_AGEMA_signal_12032, mcs1_mcs_mat1_3_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_16123, new_AGEMA_signal_16122, new_AGEMA_signal_16121, mcs1_mcs_mat1_3_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_9694, new_AGEMA_signal_9693, new_AGEMA_signal_9692, mcs1_mcs_mat1_3_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_16984, new_AGEMA_signal_16983, new_AGEMA_signal_16982, mcs1_mcs_mat1_3_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_14923, new_AGEMA_signal_14922, new_AGEMA_signal_14921, mcs1_mcs_mat1_3_mcs_out[47]}), .b ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .c ({new_AGEMA_signal_16123, new_AGEMA_signal_16122, new_AGEMA_signal_16121, mcs1_mcs_mat1_3_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_13474, new_AGEMA_signal_13473, new_AGEMA_signal_13472, mcs1_mcs_mat1_3_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .c ({new_AGEMA_signal_14923, new_AGEMA_signal_14922, new_AGEMA_signal_14921, mcs1_mcs_mat1_3_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_8863, new_AGEMA_signal_8862, new_AGEMA_signal_8861, mcs1_mcs_mat1_3_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_12037, new_AGEMA_signal_12036, new_AGEMA_signal_12035, mcs1_mcs_mat1_3_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_13474, new_AGEMA_signal_13473, new_AGEMA_signal_13472, mcs1_mcs_mat1_3_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490], Fresh[4489], Fresh[4488]}), .c ({new_AGEMA_signal_12037, new_AGEMA_signal_12036, new_AGEMA_signal_12035, mcs1_mcs_mat1_3_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494]}), .c ({new_AGEMA_signal_9694, new_AGEMA_signal_9693, new_AGEMA_signal_9692, mcs1_mcs_mat1_3_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500]}), .c ({new_AGEMA_signal_10873, new_AGEMA_signal_10872, new_AGEMA_signal_10871, mcs1_mcs_mat1_3_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_18370, new_AGEMA_signal_18369, new_AGEMA_signal_18368, mcs1_mcs_mat1_3_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_16987, new_AGEMA_signal_16986, new_AGEMA_signal_16985, mcs1_mcs_mat1_3_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_19024, new_AGEMA_signal_19023, new_AGEMA_signal_19022, mcs1_mcs_mat1_3_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_17692, new_AGEMA_signal_17691, new_AGEMA_signal_17690, mcs1_mcs_mat1_3_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_14926, new_AGEMA_signal_14925, new_AGEMA_signal_14924, mcs1_mcs_mat1_3_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_18370, new_AGEMA_signal_18369, new_AGEMA_signal_18368, mcs1_mcs_mat1_3_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_18373, new_AGEMA_signal_18372, new_AGEMA_signal_18371, mcs1_mcs_mat1_3_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_17698, new_AGEMA_signal_17697, new_AGEMA_signal_17696, mcs1_mcs_mat1_3_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_19027, new_AGEMA_signal_19026, new_AGEMA_signal_19025, mcs1_mcs_mat1_3_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_18376, new_AGEMA_signal_18375, new_AGEMA_signal_18374, mcs1_mcs_mat1_3_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_13477, new_AGEMA_signal_13476, new_AGEMA_signal_13475, mcs1_mcs_mat1_3_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_19030, new_AGEMA_signal_19029, new_AGEMA_signal_19028, mcs1_mcs_mat1_3_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_17692, new_AGEMA_signal_17691, new_AGEMA_signal_17690, mcs1_mcs_mat1_3_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_16990, new_AGEMA_signal_16989, new_AGEMA_signal_16988, mcs1_mcs_mat1_3_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_18376, new_AGEMA_signal_18375, new_AGEMA_signal_18374, mcs1_mcs_mat1_3_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_17695, new_AGEMA_signal_17694, new_AGEMA_signal_17693, mcs1_mcs_mat1_3_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_16990, new_AGEMA_signal_16989, new_AGEMA_signal_16988, mcs1_mcs_mat1_3_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_18379, new_AGEMA_signal_18378, new_AGEMA_signal_18377, mcs1_mcs_mat1_3_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4511], Fresh[4510], Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506]}), .c ({new_AGEMA_signal_17698, new_AGEMA_signal_17697, new_AGEMA_signal_17696, mcs1_mcs_mat1_3_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4517], Fresh[4516], Fresh[4515], Fresh[4514], Fresh[4513], Fresh[4512]}), .c ({new_AGEMA_signal_14926, new_AGEMA_signal_14925, new_AGEMA_signal_14924, mcs1_mcs_mat1_3_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520], Fresh[4519], Fresh[4518]}), .c ({new_AGEMA_signal_16990, new_AGEMA_signal_16989, new_AGEMA_signal_16988, mcs1_mcs_mat1_3_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_14929, new_AGEMA_signal_14928, new_AGEMA_signal_14927, mcs1_mcs_mat1_3_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_8866, new_AGEMA_signal_8865, new_AGEMA_signal_8864, mcs1_mcs_mat1_3_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_16126, new_AGEMA_signal_16125, new_AGEMA_signal_16124, mcs1_mcs_mat1_3_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_10879, new_AGEMA_signal_10878, new_AGEMA_signal_10877, mcs1_mcs_mat1_3_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_10876, new_AGEMA_signal_10875, new_AGEMA_signal_10874, mcs1_mcs_mat1_3_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_12040, new_AGEMA_signal_12039, new_AGEMA_signal_12038, mcs1_mcs_mat1_3_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({new_AGEMA_signal_14929, new_AGEMA_signal_14928, new_AGEMA_signal_14927, mcs1_mcs_mat1_3_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_16129, new_AGEMA_signal_16128, new_AGEMA_signal_16127, mcs1_mcs_mat1_3_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_12043, new_AGEMA_signal_12042, new_AGEMA_signal_12041, mcs1_mcs_mat1_3_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_13480, new_AGEMA_signal_13479, new_AGEMA_signal_13478, mcs1_mcs_mat1_3_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_14929, new_AGEMA_signal_14928, new_AGEMA_signal_14927, mcs1_mcs_mat1_3_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_12046, new_AGEMA_signal_12045, new_AGEMA_signal_12044, mcs1_mcs_mat1_3_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_10882, new_AGEMA_signal_10881, new_AGEMA_signal_10880, mcs1_mcs_mat1_3_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_13480, new_AGEMA_signal_13479, new_AGEMA_signal_13478, mcs1_mcs_mat1_3_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_12046, new_AGEMA_signal_12045, new_AGEMA_signal_12044, mcs1_mcs_mat1_3_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_10879, new_AGEMA_signal_10878, new_AGEMA_signal_10877, mcs1_mcs_mat1_3_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_13483, new_AGEMA_signal_13482, new_AGEMA_signal_13481, mcs1_mcs_mat1_3_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .b ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, new_AGEMA_signal_10310, mcs1_mcs_mat1_3_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_10879, new_AGEMA_signal_10878, new_AGEMA_signal_10877, mcs1_mcs_mat1_3_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({new_AGEMA_signal_9697, new_AGEMA_signal_9696, new_AGEMA_signal_9695, mcs1_mcs_mat1_3_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_10312, new_AGEMA_signal_10311, new_AGEMA_signal_10310, mcs1_mcs_mat1_3_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524]}), .c ({new_AGEMA_signal_12046, new_AGEMA_signal_12045, new_AGEMA_signal_12044, mcs1_mcs_mat1_3_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530]}), .c ({new_AGEMA_signal_9697, new_AGEMA_signal_9696, new_AGEMA_signal_9695, mcs1_mcs_mat1_3_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4541], Fresh[4540], Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536]}), .c ({new_AGEMA_signal_10882, new_AGEMA_signal_10881, new_AGEMA_signal_10880, mcs1_mcs_mat1_3_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_12049, new_AGEMA_signal_12048, new_AGEMA_signal_12047, mcs1_mcs_mat1_3_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_10885, new_AGEMA_signal_10884, new_AGEMA_signal_10883, mcs1_mcs_mat1_3_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_13486, new_AGEMA_signal_13485, new_AGEMA_signal_13484, mcs1_mcs_mat1_3_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_9700, new_AGEMA_signal_9699, new_AGEMA_signal_9698, mcs1_mcs_mat1_3_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_10315, new_AGEMA_signal_10314, new_AGEMA_signal_10313, mcs1_mcs_mat1_3_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_16132, new_AGEMA_signal_16131, new_AGEMA_signal_16130, mcs1_mcs_mat1_3_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_12052, new_AGEMA_signal_12051, new_AGEMA_signal_12050, mcs1_mcs_mat1_3_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_16993, new_AGEMA_signal_16992, new_AGEMA_signal_16991, mcs1_mcs_mat1_3_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4547], Fresh[4546], Fresh[4545], Fresh[4544], Fresh[4543], Fresh[4542]}), .c ({new_AGEMA_signal_12052, new_AGEMA_signal_12051, new_AGEMA_signal_12050, mcs1_mcs_mat1_3_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550], Fresh[4549], Fresh[4548]}), .c ({new_AGEMA_signal_9700, new_AGEMA_signal_9699, new_AGEMA_signal_9698, mcs1_mcs_mat1_3_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554]}), .c ({new_AGEMA_signal_10885, new_AGEMA_signal_10884, new_AGEMA_signal_10883, mcs1_mcs_mat1_3_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_14935, new_AGEMA_signal_14934, new_AGEMA_signal_14933, mcs1_mcs_mat1_3_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_13492, new_AGEMA_signal_13491, new_AGEMA_signal_13490, mcs1_mcs_mat1_3_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_16135, new_AGEMA_signal_16134, new_AGEMA_signal_16133, mcs1_mcs_mat1_3_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_9706, new_AGEMA_signal_9705, new_AGEMA_signal_9704, mcs1_mcs_mat1_3_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_13495, new_AGEMA_signal_13494, new_AGEMA_signal_13493, mcs1_mcs_mat1_3_mcs_out[29]}), .c ({new_AGEMA_signal_14935, new_AGEMA_signal_14934, new_AGEMA_signal_14933, mcs1_mcs_mat1_3_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_9703, new_AGEMA_signal_9702, new_AGEMA_signal_9701, mcs1_mcs_mat1_3_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_13492, new_AGEMA_signal_13491, new_AGEMA_signal_13490, mcs1_mcs_mat1_3_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_14938, new_AGEMA_signal_14937, new_AGEMA_signal_14936, mcs1_mcs_mat1_3_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_12061, new_AGEMA_signal_12060, new_AGEMA_signal_12059, mcs1_mcs_mat1_3_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .c ({new_AGEMA_signal_13492, new_AGEMA_signal_13491, new_AGEMA_signal_13490, mcs1_mcs_mat1_3_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_14941, new_AGEMA_signal_14940, new_AGEMA_signal_14939, mcs1_mcs_mat1_3_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_12055, new_AGEMA_signal_12054, new_AGEMA_signal_12053, mcs1_mcs_mat1_3_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_16138, new_AGEMA_signal_16137, new_AGEMA_signal_16136, mcs1_mcs_mat1_3_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_13498, new_AGEMA_signal_13497, new_AGEMA_signal_13496, mcs1_mcs_mat1_3_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_12058, new_AGEMA_signal_12057, new_AGEMA_signal_12056, mcs1_mcs_mat1_3_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_14941, new_AGEMA_signal_14940, new_AGEMA_signal_14939, mcs1_mcs_mat1_3_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_10888, new_AGEMA_signal_10887, new_AGEMA_signal_10886, mcs1_mcs_mat1_3_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_12058, new_AGEMA_signal_12057, new_AGEMA_signal_12056, mcs1_mcs_mat1_3_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_12061, new_AGEMA_signal_12060, new_AGEMA_signal_12059, mcs1_mcs_mat1_3_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_9706, new_AGEMA_signal_9705, new_AGEMA_signal_9704, mcs1_mcs_mat1_3_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_13498, new_AGEMA_signal_13497, new_AGEMA_signal_13496, mcs1_mcs_mat1_3_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560]}), .c ({new_AGEMA_signal_12061, new_AGEMA_signal_12060, new_AGEMA_signal_12059, mcs1_mcs_mat1_3_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4571], Fresh[4570], Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566]}), .c ({new_AGEMA_signal_9706, new_AGEMA_signal_9705, new_AGEMA_signal_9704, mcs1_mcs_mat1_3_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4577], Fresh[4576], Fresh[4575], Fresh[4574], Fresh[4573], Fresh[4572]}), .c ({new_AGEMA_signal_10888, new_AGEMA_signal_10887, new_AGEMA_signal_10886, mcs1_mcs_mat1_3_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_17701, new_AGEMA_signal_17700, new_AGEMA_signal_17699, mcs1_mcs_mat1_3_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_18382, new_AGEMA_signal_18381, new_AGEMA_signal_18380, mcs1_mcs_mat1_3_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_16996, new_AGEMA_signal_16995, new_AGEMA_signal_16994, mcs1_mcs_mat1_3_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_14944, new_AGEMA_signal_14943, new_AGEMA_signal_14942, mcs1_mcs_mat1_3_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_17701, new_AGEMA_signal_17700, new_AGEMA_signal_17699, mcs1_mcs_mat1_3_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_18385, new_AGEMA_signal_18384, new_AGEMA_signal_18383, mcs1_mcs_mat1_3_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_19033, new_AGEMA_signal_19032, new_AGEMA_signal_19031, mcs1_mcs_mat1_3_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_17707, new_AGEMA_signal_17706, new_AGEMA_signal_17705, mcs1_mcs_mat1_3_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_14944, new_AGEMA_signal_14943, new_AGEMA_signal_14942, mcs1_mcs_mat1_3_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_18385, new_AGEMA_signal_18384, new_AGEMA_signal_18383, mcs1_mcs_mat1_3_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_19036, new_AGEMA_signal_19035, new_AGEMA_signal_19034, mcs1_mcs_mat1_3_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .c ({new_AGEMA_signal_19753, new_AGEMA_signal_19752, new_AGEMA_signal_19751, mcs1_mcs_mat1_3_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_17707, new_AGEMA_signal_17706, new_AGEMA_signal_17705, mcs1_mcs_mat1_3_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_18388, new_AGEMA_signal_18387, new_AGEMA_signal_18386, mcs1_mcs_mat1_3_mcs_out[24]}), .c ({new_AGEMA_signal_19036, new_AGEMA_signal_19035, new_AGEMA_signal_19034, mcs1_mcs_mat1_3_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_17704, new_AGEMA_signal_17703, new_AGEMA_signal_17702, mcs1_mcs_mat1_3_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .c ({new_AGEMA_signal_18388, new_AGEMA_signal_18387, new_AGEMA_signal_18386, mcs1_mcs_mat1_3_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_16996, new_AGEMA_signal_16995, new_AGEMA_signal_16994, mcs1_mcs_mat1_3_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_13501, new_AGEMA_signal_13500, new_AGEMA_signal_13499, mcs1_mcs_mat1_3_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_17704, new_AGEMA_signal_17703, new_AGEMA_signal_17702, mcs1_mcs_mat1_3_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580], Fresh[4579], Fresh[4578]}), .c ({new_AGEMA_signal_17707, new_AGEMA_signal_17706, new_AGEMA_signal_17705, mcs1_mcs_mat1_3_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584]}), .c ({new_AGEMA_signal_14944, new_AGEMA_signal_14943, new_AGEMA_signal_14942, mcs1_mcs_mat1_3_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590]}), .c ({new_AGEMA_signal_16996, new_AGEMA_signal_16995, new_AGEMA_signal_16994, mcs1_mcs_mat1_3_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_12064, new_AGEMA_signal_12063, new_AGEMA_signal_12062, mcs1_mcs_mat1_3_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .c ({new_AGEMA_signal_13504, new_AGEMA_signal_13503, new_AGEMA_signal_13502, mcs1_mcs_mat1_3_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_10891, new_AGEMA_signal_10890, new_AGEMA_signal_10889, mcs1_mcs_mat1_3_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_9709, new_AGEMA_signal_9708, new_AGEMA_signal_9707, mcs1_mcs_mat1_3_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_12064, new_AGEMA_signal_12063, new_AGEMA_signal_12062, mcs1_mcs_mat1_3_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_13507, new_AGEMA_signal_13506, new_AGEMA_signal_13505, mcs1_mcs_mat1_3_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .c ({new_AGEMA_signal_14947, new_AGEMA_signal_14946, new_AGEMA_signal_14945, mcs1_mcs_mat1_3_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_12070, new_AGEMA_signal_12069, new_AGEMA_signal_12068, mcs1_mcs_mat1_3_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_9709, new_AGEMA_signal_9708, new_AGEMA_signal_9707, mcs1_mcs_mat1_3_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_13507, new_AGEMA_signal_13506, new_AGEMA_signal_13505, mcs1_mcs_mat1_3_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_14950, new_AGEMA_signal_14949, new_AGEMA_signal_14948, mcs1_mcs_mat1_3_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_8407, new_AGEMA_signal_8406, new_AGEMA_signal_8405, mcs1_mcs_mat1_3_mcs_out[86]}), .c ({new_AGEMA_signal_16141, new_AGEMA_signal_16140, new_AGEMA_signal_16139, mcs1_mcs_mat1_3_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_12070, new_AGEMA_signal_12069, new_AGEMA_signal_12068, mcs1_mcs_mat1_3_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_13510, new_AGEMA_signal_13509, new_AGEMA_signal_13508, mcs1_mcs_mat1_3_mcs_out[20]}), .c ({new_AGEMA_signal_14950, new_AGEMA_signal_14949, new_AGEMA_signal_14948, mcs1_mcs_mat1_3_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_12067, new_AGEMA_signal_12066, new_AGEMA_signal_12065, mcs1_mcs_mat1_3_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .c ({new_AGEMA_signal_13510, new_AGEMA_signal_13509, new_AGEMA_signal_13508, mcs1_mcs_mat1_3_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_10891, new_AGEMA_signal_10890, new_AGEMA_signal_10889, mcs1_mcs_mat1_3_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8875, new_AGEMA_signal_8874, new_AGEMA_signal_8873, mcs1_mcs_mat1_3_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_12067, new_AGEMA_signal_12066, new_AGEMA_signal_12065, mcs1_mcs_mat1_3_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4601], Fresh[4600], Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596]}), .c ({new_AGEMA_signal_12070, new_AGEMA_signal_12069, new_AGEMA_signal_12068, mcs1_mcs_mat1_3_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4607], Fresh[4606], Fresh[4605], Fresh[4604], Fresh[4603], Fresh[4602]}), .c ({new_AGEMA_signal_9709, new_AGEMA_signal_9708, new_AGEMA_signal_9707, mcs1_mcs_mat1_3_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610], Fresh[4609], Fresh[4608]}), .c ({new_AGEMA_signal_10891, new_AGEMA_signal_10890, new_AGEMA_signal_10889, mcs1_mcs_mat1_3_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_12073, new_AGEMA_signal_12072, new_AGEMA_signal_12071, mcs1_mcs_mat1_3_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_12082, new_AGEMA_signal_12081, new_AGEMA_signal_12080, mcs1_mcs_mat1_3_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_13513, new_AGEMA_signal_13512, new_AGEMA_signal_13511, mcs1_mcs_mat1_3_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_13516, new_AGEMA_signal_13515, new_AGEMA_signal_13514, mcs1_mcs_mat1_3_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_8878, new_AGEMA_signal_8877, new_AGEMA_signal_8876, mcs1_mcs_mat1_3_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_14953, new_AGEMA_signal_14952, new_AGEMA_signal_14951, mcs1_mcs_mat1_3_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_14956, new_AGEMA_signal_14955, new_AGEMA_signal_14954, mcs1_mcs_mat1_3_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_9712, new_AGEMA_signal_9711, new_AGEMA_signal_9710, mcs1_mcs_mat1_3_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_16144, new_AGEMA_signal_16143, new_AGEMA_signal_16142, mcs1_mcs_mat1_3_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8424, new_AGEMA_signal_8423, mcs1_mcs_mat1_3_mcs_out[50]}), .b ({new_AGEMA_signal_13516, new_AGEMA_signal_13515, new_AGEMA_signal_13514, mcs1_mcs_mat1_3_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_14956, new_AGEMA_signal_14955, new_AGEMA_signal_14954, mcs1_mcs_mat1_3_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_12076, new_AGEMA_signal_12075, new_AGEMA_signal_12074, mcs1_mcs_mat1_3_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .c ({new_AGEMA_signal_13516, new_AGEMA_signal_13515, new_AGEMA_signal_13514, mcs1_mcs_mat1_3_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_10894, new_AGEMA_signal_10893, new_AGEMA_signal_10892, mcs1_mcs_mat1_3_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_10897, new_AGEMA_signal_10896, new_AGEMA_signal_10895, mcs1_mcs_mat1_3_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_12076, new_AGEMA_signal_12075, new_AGEMA_signal_12074, mcs1_mcs_mat1_3_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_12079, new_AGEMA_signal_12078, new_AGEMA_signal_12077, mcs1_mcs_mat1_3_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_9712, new_AGEMA_signal_9711, new_AGEMA_signal_9710, mcs1_mcs_mat1_3_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_13519, new_AGEMA_signal_13518, new_AGEMA_signal_13517, mcs1_mcs_mat1_3_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614]}), .c ({new_AGEMA_signal_12082, new_AGEMA_signal_12081, new_AGEMA_signal_12080, mcs1_mcs_mat1_3_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620]}), .c ({new_AGEMA_signal_9712, new_AGEMA_signal_9711, new_AGEMA_signal_9710, mcs1_mcs_mat1_3_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4631], Fresh[4630], Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626]}), .c ({new_AGEMA_signal_10897, new_AGEMA_signal_10896, new_AGEMA_signal_10895, mcs1_mcs_mat1_3_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_14965, new_AGEMA_signal_14964, new_AGEMA_signal_14963, mcs1_mcs_mat1_3_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, new_AGEMA_signal_10316, mcs1_mcs_mat1_3_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_16147, new_AGEMA_signal_16146, new_AGEMA_signal_16145, mcs1_mcs_mat1_3_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_13528, new_AGEMA_signal_13527, new_AGEMA_signal_13526, mcs1_mcs_mat1_3_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_13522, new_AGEMA_signal_13521, new_AGEMA_signal_13520, mcs1_mcs_mat1_3_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_14959, new_AGEMA_signal_14958, new_AGEMA_signal_14957, mcs1_mcs_mat1_3_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_12088, new_AGEMA_signal_12087, new_AGEMA_signal_12086, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_9715, new_AGEMA_signal_9714, new_AGEMA_signal_9713, mcs1_mcs_mat1_3_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_13522, new_AGEMA_signal_13521, new_AGEMA_signal_13520, mcs1_mcs_mat1_3_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, new_AGEMA_signal_10316, mcs1_mcs_mat1_3_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_13525, new_AGEMA_signal_13524, new_AGEMA_signal_13523, mcs1_mcs_mat1_3_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_14962, new_AGEMA_signal_14961, new_AGEMA_signal_14960, mcs1_mcs_mat1_3_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_12085, new_AGEMA_signal_12084, new_AGEMA_signal_12083, mcs1_mcs_mat1_3_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_12088, new_AGEMA_signal_12087, new_AGEMA_signal_12086, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_13525, new_AGEMA_signal_13524, new_AGEMA_signal_13523, mcs1_mcs_mat1_3_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8880, new_AGEMA_signal_8879, mcs1_mcs_mat1_3_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_9715, new_AGEMA_signal_9714, new_AGEMA_signal_9713, mcs1_mcs_mat1_3_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_10318, new_AGEMA_signal_10317, new_AGEMA_signal_10316, mcs1_mcs_mat1_3_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_16150, new_AGEMA_signal_16149, new_AGEMA_signal_16148, mcs1_mcs_mat1_3_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .c ({new_AGEMA_signal_16999, new_AGEMA_signal_16998, new_AGEMA_signal_16997, mcs1_mcs_mat1_3_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_14965, new_AGEMA_signal_14964, new_AGEMA_signal_14963, mcs1_mcs_mat1_3_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_12088, new_AGEMA_signal_12087, new_AGEMA_signal_12086, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_16150, new_AGEMA_signal_16149, new_AGEMA_signal_16148, mcs1_mcs_mat1_3_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({new_AGEMA_signal_13528, new_AGEMA_signal_13527, new_AGEMA_signal_13526, mcs1_mcs_mat1_3_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_14965, new_AGEMA_signal_14964, new_AGEMA_signal_14963, mcs1_mcs_mat1_3_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({new_AGEMA_signal_12085, new_AGEMA_signal_12084, new_AGEMA_signal_12083, mcs1_mcs_mat1_3_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_13528, new_AGEMA_signal_13527, new_AGEMA_signal_13526, mcs1_mcs_mat1_3_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_8371, new_AGEMA_signal_8370, new_AGEMA_signal_8369, shiftr_out[112]}), .b ({new_AGEMA_signal_10900, new_AGEMA_signal_10899, new_AGEMA_signal_10898, mcs1_mcs_mat1_3_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_12085, new_AGEMA_signal_12084, new_AGEMA_signal_12083, mcs1_mcs_mat1_3_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10411, new_AGEMA_signal_10410, new_AGEMA_signal_10409, mcs1_mcs_mat1_3_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4637], Fresh[4636], Fresh[4635], Fresh[4634], Fresh[4633], Fresh[4632]}), .c ({new_AGEMA_signal_12088, new_AGEMA_signal_12087, new_AGEMA_signal_12086, mcs1_mcs_mat1_3_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8575, new_AGEMA_signal_8574, new_AGEMA_signal_8573, mcs1_mcs_mat1_3_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640], Fresh[4639], Fresh[4638]}), .c ({new_AGEMA_signal_9715, new_AGEMA_signal_9714, new_AGEMA_signal_9713, mcs1_mcs_mat1_3_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10212, new_AGEMA_signal_10211, mcs1_mcs_mat1_3_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644]}), .c ({new_AGEMA_signal_10900, new_AGEMA_signal_10899, new_AGEMA_signal_10898, mcs1_mcs_mat1_3_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_16153, new_AGEMA_signal_16152, new_AGEMA_signal_16151, mcs1_mcs_mat1_3_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .c ({new_AGEMA_signal_17002, new_AGEMA_signal_17001, new_AGEMA_signal_17000, mcs1_mcs_mat1_3_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_18394, new_AGEMA_signal_18393, new_AGEMA_signal_18392, mcs1_mcs_mat1_3_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .c ({new_AGEMA_signal_19039, new_AGEMA_signal_19038, new_AGEMA_signal_19037, mcs1_mcs_mat1_3_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_17710, new_AGEMA_signal_17709, new_AGEMA_signal_17708, mcs1_mcs_mat1_3_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .c ({new_AGEMA_signal_18391, new_AGEMA_signal_18390, new_AGEMA_signal_18389, mcs1_mcs_mat1_3_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_17005, new_AGEMA_signal_17004, new_AGEMA_signal_17003, mcs1_mcs_mat1_3_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_16153, new_AGEMA_signal_16152, new_AGEMA_signal_16151, mcs1_mcs_mat1_3_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_17710, new_AGEMA_signal_17709, new_AGEMA_signal_17708, mcs1_mcs_mat1_3_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_13531, new_AGEMA_signal_13530, new_AGEMA_signal_13529, mcs1_mcs_mat1_3_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_14968, new_AGEMA_signal_14967, new_AGEMA_signal_14966, mcs1_mcs_mat1_3_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_16153, new_AGEMA_signal_16152, new_AGEMA_signal_16151, mcs1_mcs_mat1_3_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_19042, new_AGEMA_signal_19041, new_AGEMA_signal_19040, mcs1_mcs_mat1_3_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_11389, new_AGEMA_signal_11388, new_AGEMA_signal_11387, shiftr_out[80]}), .c ({new_AGEMA_signal_19756, new_AGEMA_signal_19755, new_AGEMA_signal_19754, mcs1_mcs_mat1_3_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_13531, new_AGEMA_signal_13530, new_AGEMA_signal_13529, mcs1_mcs_mat1_3_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_18394, new_AGEMA_signal_18393, new_AGEMA_signal_18392, mcs1_mcs_mat1_3_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_19042, new_AGEMA_signal_19041, new_AGEMA_signal_19040, mcs1_mcs_mat1_3_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_17713, new_AGEMA_signal_17712, new_AGEMA_signal_17711, mcs1_mcs_mat1_3_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_17005, new_AGEMA_signal_17004, new_AGEMA_signal_17003, mcs1_mcs_mat1_3_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_18394, new_AGEMA_signal_18393, new_AGEMA_signal_18392, mcs1_mcs_mat1_3_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16615, new_AGEMA_signal_16614, new_AGEMA_signal_16613, mcs1_mcs_mat1_3_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650]}), .c ({new_AGEMA_signal_17713, new_AGEMA_signal_17712, new_AGEMA_signal_17711, mcs1_mcs_mat1_3_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12829, new_AGEMA_signal_12828, new_AGEMA_signal_12827, mcs1_mcs_mat1_3_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4661], Fresh[4660], Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656]}), .c ({new_AGEMA_signal_14968, new_AGEMA_signal_14967, new_AGEMA_signal_14966, mcs1_mcs_mat1_3_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15703, new_AGEMA_signal_15702, new_AGEMA_signal_15701, shiftr_out[83]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4667], Fresh[4666], Fresh[4665], Fresh[4664], Fresh[4663], Fresh[4662]}), .c ({new_AGEMA_signal_17005, new_AGEMA_signal_17004, new_AGEMA_signal_17003, mcs1_mcs_mat1_3_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_17008, new_AGEMA_signal_17007, new_AGEMA_signal_17006, mcs1_mcs_mat1_3_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_10906, new_AGEMA_signal_10905, new_AGEMA_signal_10904, mcs1_mcs_mat1_3_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_17716, new_AGEMA_signal_17715, new_AGEMA_signal_17714, mcs1_mcs_mat1_3_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_16156, new_AGEMA_signal_16155, new_AGEMA_signal_16154, mcs1_mcs_mat1_3_mcs_out[7]}), .b ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .c ({new_AGEMA_signal_17008, new_AGEMA_signal_17007, new_AGEMA_signal_17006, mcs1_mcs_mat1_3_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_14971, new_AGEMA_signal_14970, new_AGEMA_signal_14969, mcs1_mcs_mat1_3_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .c ({new_AGEMA_signal_16156, new_AGEMA_signal_16155, new_AGEMA_signal_16154, mcs1_mcs_mat1_3_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_13534, new_AGEMA_signal_13533, new_AGEMA_signal_13532, mcs1_mcs_mat1_3_mcs_out[6]}), .b ({new_AGEMA_signal_9721, new_AGEMA_signal_9720, new_AGEMA_signal_9719, mcs1_mcs_mat1_3_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_14971, new_AGEMA_signal_14970, new_AGEMA_signal_14969, mcs1_mcs_mat1_3_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_9718, new_AGEMA_signal_9717, new_AGEMA_signal_9716, mcs1_mcs_mat1_3_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_12091, new_AGEMA_signal_12090, new_AGEMA_signal_12089, mcs1_mcs_mat1_3_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_13534, new_AGEMA_signal_13533, new_AGEMA_signal_13532, mcs1_mcs_mat1_3_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10447, new_AGEMA_signal_10446, new_AGEMA_signal_10445, shiftr_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670], Fresh[4669], Fresh[4668]}), .c ({new_AGEMA_signal_12091, new_AGEMA_signal_12090, new_AGEMA_signal_12089, mcs1_mcs_mat1_3_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8611, new_AGEMA_signal_8610, new_AGEMA_signal_8609, shiftr_out[50]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674]}), .c ({new_AGEMA_signal_9721, new_AGEMA_signal_9720, new_AGEMA_signal_9719, mcs1_mcs_mat1_3_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10248, new_AGEMA_signal_10247, mcs1_mcs_mat1_3_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680]}), .c ({new_AGEMA_signal_10906, new_AGEMA_signal_10905, new_AGEMA_signal_10904, mcs1_mcs_mat1_3_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_10909, new_AGEMA_signal_10908, new_AGEMA_signal_10907, mcs1_mcs_mat1_3_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_12094, new_AGEMA_signal_12093, new_AGEMA_signal_12092, mcs1_mcs_mat1_3_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_13540, new_AGEMA_signal_13539, new_AGEMA_signal_13538, mcs1_mcs_mat1_3_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .b ({new_AGEMA_signal_10912, new_AGEMA_signal_10911, new_AGEMA_signal_10910, mcs1_mcs_mat1_3_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_12094, new_AGEMA_signal_12093, new_AGEMA_signal_12092, mcs1_mcs_mat1_3_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_13543, new_AGEMA_signal_13542, new_AGEMA_signal_13541, mcs1_mcs_mat1_3_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_9724, new_AGEMA_signal_9723, new_AGEMA_signal_9722, mcs1_mcs_mat1_3_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_14974, new_AGEMA_signal_14973, new_AGEMA_signal_14972, mcs1_mcs_mat1_3_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_13546, new_AGEMA_signal_13545, new_AGEMA_signal_13544, mcs1_mcs_mat1_3_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_12100, new_AGEMA_signal_12099, new_AGEMA_signal_12098, mcs1_mcs_mat1_3_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_14977, new_AGEMA_signal_14976, new_AGEMA_signal_14975, mcs1_mcs_mat1_3_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_12103, new_AGEMA_signal_12102, new_AGEMA_signal_12101, mcs1_mcs_mat1_3_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_8887, new_AGEMA_signal_8886, new_AGEMA_signal_8885, mcs1_mcs_mat1_3_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_13546, new_AGEMA_signal_13545, new_AGEMA_signal_13544, mcs1_mcs_mat1_3_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10464, new_AGEMA_signal_10463, shiftr_out[17]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4691], Fresh[4690], Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686]}), .c ({new_AGEMA_signal_12103, new_AGEMA_signal_12102, new_AGEMA_signal_12101, mcs1_mcs_mat1_3_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8628, new_AGEMA_signal_8627, shiftr_out[18]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4697], Fresh[4696], Fresh[4695], Fresh[4694], Fresh[4693], Fresh[4692]}), .c ({new_AGEMA_signal_9724, new_AGEMA_signal_9723, new_AGEMA_signal_9722, mcs1_mcs_mat1_3_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_3_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10267, new_AGEMA_signal_10266, new_AGEMA_signal_10265, mcs1_mcs_mat1_3_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700], Fresh[4699], Fresh[4698]}), .c ({new_AGEMA_signal_10912, new_AGEMA_signal_10911, new_AGEMA_signal_10910, mcs1_mcs_mat1_3_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U96 ( .a ({new_AGEMA_signal_17011, new_AGEMA_signal_17010, new_AGEMA_signal_17009, mcs1_mcs_mat1_4_n128}), .b ({new_AGEMA_signal_18397, new_AGEMA_signal_18396, new_AGEMA_signal_18395, mcs1_mcs_mat1_4_n127}), .c ({temp_next_s3[77], temp_next_s2[77], temp_next_s1[77], temp_next_s0[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U95 ( .a ({new_AGEMA_signal_15109, new_AGEMA_signal_15108, new_AGEMA_signal_15107, mcs1_mcs_mat1_4_mcs_out[41]}), .b ({new_AGEMA_signal_17773, new_AGEMA_signal_17772, new_AGEMA_signal_17771, mcs1_mcs_mat1_4_mcs_out[45]}), .c ({new_AGEMA_signal_18397, new_AGEMA_signal_18396, new_AGEMA_signal_18395, mcs1_mcs_mat1_4_n127}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U94 ( .a ({new_AGEMA_signal_10327, new_AGEMA_signal_10326, new_AGEMA_signal_10325, mcs1_mcs_mat1_4_mcs_out[33]}), .b ({new_AGEMA_signal_16231, new_AGEMA_signal_16230, new_AGEMA_signal_16229, mcs1_mcs_mat1_4_mcs_out[37]}), .c ({new_AGEMA_signal_17011, new_AGEMA_signal_17010, new_AGEMA_signal_17009, mcs1_mcs_mat1_4_n128}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U93 ( .a ({new_AGEMA_signal_17719, new_AGEMA_signal_17718, new_AGEMA_signal_17717, mcs1_mcs_mat1_4_n126}), .b ({new_AGEMA_signal_21241, new_AGEMA_signal_21240, new_AGEMA_signal_21239, mcs1_mcs_mat1_4_n125}), .c ({temp_next_s3[76], temp_next_s2[76], temp_next_s1[76], temp_next_s0[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U92 ( .a ({new_AGEMA_signal_13660, new_AGEMA_signal_13659, new_AGEMA_signal_13658, mcs1_mcs_mat1_4_mcs_out[40]}), .b ({new_AGEMA_signal_20620, new_AGEMA_signal_20619, new_AGEMA_signal_20618, mcs1_mcs_mat1_4_mcs_out[44]}), .c ({new_AGEMA_signal_21241, new_AGEMA_signal_21240, new_AGEMA_signal_21239, mcs1_mcs_mat1_4_n125}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U91 ( .a ({new_AGEMA_signal_17092, new_AGEMA_signal_17091, new_AGEMA_signal_17090, mcs1_mcs_mat1_4_mcs_out[32]}), .b ({new_AGEMA_signal_13666, new_AGEMA_signal_13665, new_AGEMA_signal_13664, mcs1_mcs_mat1_4_mcs_out[36]}), .c ({new_AGEMA_signal_17719, new_AGEMA_signal_17718, new_AGEMA_signal_17717, mcs1_mcs_mat1_4_n126}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U90 ( .a ({new_AGEMA_signal_14980, new_AGEMA_signal_14979, new_AGEMA_signal_14978, mcs1_mcs_mat1_4_n124}), .b ({new_AGEMA_signal_20569, new_AGEMA_signal_20568, new_AGEMA_signal_20567, mcs1_mcs_mat1_4_n123}), .c ({temp_next_s3[47], temp_next_s2[47], temp_next_s1[47], temp_next_s0[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U89 ( .a ({new_AGEMA_signal_13678, new_AGEMA_signal_13677, new_AGEMA_signal_13676, mcs1_mcs_mat1_4_mcs_out[27]}), .b ({new_AGEMA_signal_19813, new_AGEMA_signal_19812, new_AGEMA_signal_19811, mcs1_mcs_mat1_4_mcs_out[31]}), .c ({new_AGEMA_signal_20569, new_AGEMA_signal_20568, new_AGEMA_signal_20567, mcs1_mcs_mat1_4_n123}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U88 ( .a ({new_AGEMA_signal_13696, new_AGEMA_signal_13695, new_AGEMA_signal_13694, mcs1_mcs_mat1_4_mcs_out[19]}), .b ({new_AGEMA_signal_13687, new_AGEMA_signal_13686, new_AGEMA_signal_13685, mcs1_mcs_mat1_4_mcs_out[23]}), .c ({new_AGEMA_signal_14980, new_AGEMA_signal_14979, new_AGEMA_signal_14978, mcs1_mcs_mat1_4_n124}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U87 ( .a ({new_AGEMA_signal_16159, new_AGEMA_signal_16158, new_AGEMA_signal_16157, mcs1_mcs_mat1_4_n122}), .b ({new_AGEMA_signal_19759, new_AGEMA_signal_19758, new_AGEMA_signal_19757, mcs1_mcs_mat1_4_n121}), .c ({temp_next_s3[46], temp_next_s2[46], temp_next_s1[46], temp_next_s0[46]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U86 ( .a ({new_AGEMA_signal_15124, new_AGEMA_signal_15123, new_AGEMA_signal_15122, mcs1_mcs_mat1_4_mcs_out[26]}), .b ({new_AGEMA_signal_19096, new_AGEMA_signal_19095, new_AGEMA_signal_19094, mcs1_mcs_mat1_4_mcs_out[30]}), .c ({new_AGEMA_signal_19759, new_AGEMA_signal_19758, new_AGEMA_signal_19757, mcs1_mcs_mat1_4_n121}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U85 ( .a ({new_AGEMA_signal_15136, new_AGEMA_signal_15135, new_AGEMA_signal_15134, mcs1_mcs_mat1_4_mcs_out[18]}), .b ({new_AGEMA_signal_15130, new_AGEMA_signal_15129, new_AGEMA_signal_15128, mcs1_mcs_mat1_4_mcs_out[22]}), .c ({new_AGEMA_signal_16159, new_AGEMA_signal_16158, new_AGEMA_signal_16157, mcs1_mcs_mat1_4_n122}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U84 ( .a ({new_AGEMA_signal_17014, new_AGEMA_signal_17013, new_AGEMA_signal_17012, mcs1_mcs_mat1_4_n120}), .b ({new_AGEMA_signal_19048, new_AGEMA_signal_19047, new_AGEMA_signal_19046, mcs1_mcs_mat1_4_n119}), .c ({temp_next_s3[45], temp_next_s2[45], temp_next_s1[45], temp_next_s0[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U83 ( .a ({new_AGEMA_signal_16237, new_AGEMA_signal_16236, new_AGEMA_signal_16235, mcs1_mcs_mat1_4_mcs_out[25]}), .b ({new_AGEMA_signal_18448, new_AGEMA_signal_18447, new_AGEMA_signal_18446, mcs1_mcs_mat1_4_mcs_out[29]}), .c ({new_AGEMA_signal_19048, new_AGEMA_signal_19047, new_AGEMA_signal_19046, mcs1_mcs_mat1_4_n119}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U82 ( .a ({new_AGEMA_signal_16243, new_AGEMA_signal_16242, new_AGEMA_signal_16241, mcs1_mcs_mat1_4_mcs_out[17]}), .b ({new_AGEMA_signal_16240, new_AGEMA_signal_16239, new_AGEMA_signal_16238, mcs1_mcs_mat1_4_mcs_out[21]}), .c ({new_AGEMA_signal_17014, new_AGEMA_signal_17013, new_AGEMA_signal_17012, mcs1_mcs_mat1_4_n120}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U81 ( .a ({new_AGEMA_signal_14983, new_AGEMA_signal_14982, new_AGEMA_signal_14981, mcs1_mcs_mat1_4_n118}), .b ({new_AGEMA_signal_20575, new_AGEMA_signal_20574, new_AGEMA_signal_20573, mcs1_mcs_mat1_4_n117}), .c ({temp_next_s3[44], temp_next_s2[44], temp_next_s1[44], temp_next_s0[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U80 ( .a ({new_AGEMA_signal_13684, new_AGEMA_signal_13683, new_AGEMA_signal_13682, mcs1_mcs_mat1_4_mcs_out[24]}), .b ({new_AGEMA_signal_19816, new_AGEMA_signal_19815, new_AGEMA_signal_19814, mcs1_mcs_mat1_4_mcs_out[28]}), .c ({new_AGEMA_signal_20575, new_AGEMA_signal_20574, new_AGEMA_signal_20573, mcs1_mcs_mat1_4_n117}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U79 ( .a ({new_AGEMA_signal_13702, new_AGEMA_signal_13701, new_AGEMA_signal_13700, mcs1_mcs_mat1_4_mcs_out[16]}), .b ({new_AGEMA_signal_13693, new_AGEMA_signal_13692, new_AGEMA_signal_13691, mcs1_mcs_mat1_4_mcs_out[20]}), .c ({new_AGEMA_signal_14983, new_AGEMA_signal_14982, new_AGEMA_signal_14981, mcs1_mcs_mat1_4_n118}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U78 ( .a ({new_AGEMA_signal_20578, new_AGEMA_signal_20577, new_AGEMA_signal_20576, mcs1_mcs_mat1_4_n116}), .b ({new_AGEMA_signal_17017, new_AGEMA_signal_17016, new_AGEMA_signal_17015, mcs1_mcs_mat1_4_n115}), .c ({temp_next_s3[15], temp_next_s2[15], temp_next_s1[15], temp_next_s0[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U77 ( .a ({new_AGEMA_signal_13717, new_AGEMA_signal_13716, new_AGEMA_signal_13715, mcs1_mcs_mat1_4_mcs_out[3]}), .b ({new_AGEMA_signal_16252, new_AGEMA_signal_16251, new_AGEMA_signal_16250, mcs1_mcs_mat1_4_mcs_out[7]}), .c ({new_AGEMA_signal_17017, new_AGEMA_signal_17016, new_AGEMA_signal_17015, mcs1_mcs_mat1_4_n115}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U76 ( .a ({new_AGEMA_signal_11011, new_AGEMA_signal_11010, new_AGEMA_signal_11009, mcs1_mcs_mat1_4_mcs_out[11]}), .b ({new_AGEMA_signal_19819, new_AGEMA_signal_19818, new_AGEMA_signal_19817, mcs1_mcs_mat1_4_mcs_out[15]}), .c ({new_AGEMA_signal_20578, new_AGEMA_signal_20577, new_AGEMA_signal_20576, mcs1_mcs_mat1_4_n116}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U75 ( .a ({new_AGEMA_signal_17023, new_AGEMA_signal_17022, new_AGEMA_signal_17021, mcs1_mcs_mat1_4_n114}), .b ({new_AGEMA_signal_17020, new_AGEMA_signal_17019, new_AGEMA_signal_17018, mcs1_mcs_mat1_4_n113}), .c ({new_AGEMA_signal_17722, new_AGEMA_signal_17721, new_AGEMA_signal_17720, mcs_out[239]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U74 ( .a ({new_AGEMA_signal_16183, new_AGEMA_signal_16182, new_AGEMA_signal_16181, mcs1_mcs_mat1_4_mcs_out[123]}), .b ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_17020, new_AGEMA_signal_17019, new_AGEMA_signal_17018, mcs1_mcs_mat1_4_n113}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U73 ( .a ({new_AGEMA_signal_15022, new_AGEMA_signal_15021, new_AGEMA_signal_15020, mcs1_mcs_mat1_4_mcs_out[115]}), .b ({new_AGEMA_signal_16189, new_AGEMA_signal_16188, new_AGEMA_signal_16187, mcs1_mcs_mat1_4_mcs_out[119]}), .c ({new_AGEMA_signal_17023, new_AGEMA_signal_17022, new_AGEMA_signal_17021, mcs1_mcs_mat1_4_n114}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U72 ( .a ({new_AGEMA_signal_17026, new_AGEMA_signal_17025, new_AGEMA_signal_17024, mcs1_mcs_mat1_4_n112}), .b ({new_AGEMA_signal_17725, new_AGEMA_signal_17724, new_AGEMA_signal_17723, mcs1_mcs_mat1_4_n111}), .c ({new_AGEMA_signal_18400, new_AGEMA_signal_18399, new_AGEMA_signal_18398, mcs_out[238]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U71 ( .a ({new_AGEMA_signal_12106, new_AGEMA_signal_12105, new_AGEMA_signal_12104, mcs1_mcs_mat1_4_mcs_out[122]}), .b ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_17725, new_AGEMA_signal_17724, new_AGEMA_signal_17723, mcs1_mcs_mat1_4_n111}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U70 ( .a ({new_AGEMA_signal_13561, new_AGEMA_signal_13560, new_AGEMA_signal_13559, mcs1_mcs_mat1_4_mcs_out[114]}), .b ({new_AGEMA_signal_16192, new_AGEMA_signal_16191, new_AGEMA_signal_16190, mcs1_mcs_mat1_4_mcs_out[118]}), .c ({new_AGEMA_signal_17026, new_AGEMA_signal_17025, new_AGEMA_signal_17024, mcs1_mcs_mat1_4_n112}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U69 ( .a ({new_AGEMA_signal_19765, new_AGEMA_signal_19764, new_AGEMA_signal_19763, mcs1_mcs_mat1_4_n110}), .b ({new_AGEMA_signal_14986, new_AGEMA_signal_14985, new_AGEMA_signal_14984, mcs1_mcs_mat1_4_n109}), .c ({temp_next_s3[14], temp_next_s2[14], temp_next_s1[14], temp_next_s0[14]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U68 ( .a ({new_AGEMA_signal_13720, new_AGEMA_signal_13719, new_AGEMA_signal_13718, mcs1_mcs_mat1_4_mcs_out[2]}), .b ({new_AGEMA_signal_13714, new_AGEMA_signal_13713, new_AGEMA_signal_13712, mcs1_mcs_mat1_4_mcs_out[6]}), .c ({new_AGEMA_signal_14986, new_AGEMA_signal_14985, new_AGEMA_signal_14984, mcs1_mcs_mat1_4_n109}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U67 ( .a ({new_AGEMA_signal_15145, new_AGEMA_signal_15144, new_AGEMA_signal_15143, mcs1_mcs_mat1_4_mcs_out[10]}), .b ({new_AGEMA_signal_19102, new_AGEMA_signal_19101, new_AGEMA_signal_19100, mcs1_mcs_mat1_4_mcs_out[14]}), .c ({new_AGEMA_signal_19765, new_AGEMA_signal_19764, new_AGEMA_signal_19763, mcs1_mcs_mat1_4_n110}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U66 ( .a ({new_AGEMA_signal_16162, new_AGEMA_signal_16161, new_AGEMA_signal_16160, mcs1_mcs_mat1_4_n108}), .b ({new_AGEMA_signal_17728, new_AGEMA_signal_17727, new_AGEMA_signal_17726, mcs1_mcs_mat1_4_n107}), .c ({new_AGEMA_signal_18403, new_AGEMA_signal_18402, new_AGEMA_signal_18401, mcs_out[237]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U65 ( .a ({new_AGEMA_signal_16186, new_AGEMA_signal_16185, new_AGEMA_signal_16184, mcs1_mcs_mat1_4_mcs_out[121]}), .b ({new_AGEMA_signal_17059, new_AGEMA_signal_17058, new_AGEMA_signal_17057, mcs1_mcs_mat1_4_mcs_out[125]}), .c ({new_AGEMA_signal_17728, new_AGEMA_signal_17727, new_AGEMA_signal_17726, mcs1_mcs_mat1_4_n107}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U64 ( .a ({new_AGEMA_signal_12121, new_AGEMA_signal_12120, new_AGEMA_signal_12119, mcs1_mcs_mat1_4_mcs_out[113]}), .b ({new_AGEMA_signal_15019, new_AGEMA_signal_15018, new_AGEMA_signal_15017, mcs1_mcs_mat1_4_mcs_out[117]}), .c ({new_AGEMA_signal_16162, new_AGEMA_signal_16161, new_AGEMA_signal_16160, mcs1_mcs_mat1_4_n108}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U63 ( .a ({new_AGEMA_signal_17032, new_AGEMA_signal_17031, new_AGEMA_signal_17030, mcs1_mcs_mat1_4_n106}), .b ({new_AGEMA_signal_17029, new_AGEMA_signal_17028, new_AGEMA_signal_17027, mcs1_mcs_mat1_4_n105}), .c ({new_AGEMA_signal_17731, new_AGEMA_signal_17730, new_AGEMA_signal_17729, mcs_out[236]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U62 ( .a ({new_AGEMA_signal_15010, new_AGEMA_signal_15009, new_AGEMA_signal_15008, mcs1_mcs_mat1_4_mcs_out[120]}), .b ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_17029, new_AGEMA_signal_17028, new_AGEMA_signal_17027, mcs1_mcs_mat1_4_n105}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U61 ( .a ({new_AGEMA_signal_16195, new_AGEMA_signal_16194, new_AGEMA_signal_16193, mcs1_mcs_mat1_4_mcs_out[112]}), .b ({new_AGEMA_signal_13558, new_AGEMA_signal_13557, new_AGEMA_signal_13556, mcs1_mcs_mat1_4_mcs_out[116]}), .c ({new_AGEMA_signal_17032, new_AGEMA_signal_17031, new_AGEMA_signal_17030, mcs1_mcs_mat1_4_n106}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U60 ( .a ({new_AGEMA_signal_16165, new_AGEMA_signal_16164, new_AGEMA_signal_16163, mcs1_mcs_mat1_4_n104}), .b ({new_AGEMA_signal_20584, new_AGEMA_signal_20583, new_AGEMA_signal_20582, mcs1_mcs_mat1_4_n103}), .c ({new_AGEMA_signal_21253, new_AGEMA_signal_21252, new_AGEMA_signal_21251, mcs_out[207]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U59 ( .a ({new_AGEMA_signal_19789, new_AGEMA_signal_19788, new_AGEMA_signal_19787, mcs1_mcs_mat1_4_mcs_out[111]}), .b ({new_AGEMA_signal_16201, new_AGEMA_signal_16200, new_AGEMA_signal_16199, mcs1_mcs_mat1_4_mcs_out[99]}), .c ({new_AGEMA_signal_20584, new_AGEMA_signal_20583, new_AGEMA_signal_20582, mcs1_mcs_mat1_4_n103}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U58 ( .a ({new_AGEMA_signal_15043, new_AGEMA_signal_15042, new_AGEMA_signal_15041, mcs1_mcs_mat1_4_mcs_out[103]}), .b ({new_AGEMA_signal_15031, new_AGEMA_signal_15030, new_AGEMA_signal_15029, mcs1_mcs_mat1_4_mcs_out[107]}), .c ({new_AGEMA_signal_16165, new_AGEMA_signal_16164, new_AGEMA_signal_16163, mcs1_mcs_mat1_4_n104}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U57 ( .a ({new_AGEMA_signal_16168, new_AGEMA_signal_16167, new_AGEMA_signal_16166, mcs1_mcs_mat1_4_n102}), .b ({new_AGEMA_signal_20587, new_AGEMA_signal_20586, new_AGEMA_signal_20585, mcs1_mcs_mat1_4_n101}), .c ({new_AGEMA_signal_21256, new_AGEMA_signal_21255, new_AGEMA_signal_21254, mcs_out[206]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U56 ( .a ({new_AGEMA_signal_19792, new_AGEMA_signal_19791, new_AGEMA_signal_19790, mcs1_mcs_mat1_4_mcs_out[110]}), .b ({new_AGEMA_signal_13588, new_AGEMA_signal_13587, new_AGEMA_signal_13586, mcs1_mcs_mat1_4_mcs_out[98]}), .c ({new_AGEMA_signal_20587, new_AGEMA_signal_20586, new_AGEMA_signal_20585, mcs1_mcs_mat1_4_n101}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U55 ( .a ({new_AGEMA_signal_12136, new_AGEMA_signal_12135, new_AGEMA_signal_12134, mcs1_mcs_mat1_4_mcs_out[102]}), .b ({new_AGEMA_signal_15034, new_AGEMA_signal_15033, new_AGEMA_signal_15032, mcs1_mcs_mat1_4_mcs_out[106]}), .c ({new_AGEMA_signal_16168, new_AGEMA_signal_16167, new_AGEMA_signal_16166, mcs1_mcs_mat1_4_n102}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U54 ( .a ({new_AGEMA_signal_16171, new_AGEMA_signal_16170, new_AGEMA_signal_16169, mcs1_mcs_mat1_4_n100}), .b ({new_AGEMA_signal_20590, new_AGEMA_signal_20589, new_AGEMA_signal_20588, mcs1_mcs_mat1_4_n99}), .c ({new_AGEMA_signal_21259, new_AGEMA_signal_21258, new_AGEMA_signal_21257, mcs_out[205]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U53 ( .a ({new_AGEMA_signal_19795, new_AGEMA_signal_19794, new_AGEMA_signal_19793, mcs1_mcs_mat1_4_mcs_out[109]}), .b ({new_AGEMA_signal_10948, new_AGEMA_signal_10947, new_AGEMA_signal_10946, mcs1_mcs_mat1_4_mcs_out[97]}), .c ({new_AGEMA_signal_20590, new_AGEMA_signal_20589, new_AGEMA_signal_20588, mcs1_mcs_mat1_4_n99}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U52 ( .a ({new_AGEMA_signal_13582, new_AGEMA_signal_13581, new_AGEMA_signal_13580, mcs1_mcs_mat1_4_mcs_out[101]}), .b ({new_AGEMA_signal_15037, new_AGEMA_signal_15036, new_AGEMA_signal_15035, mcs1_mcs_mat1_4_mcs_out[105]}), .c ({new_AGEMA_signal_16171, new_AGEMA_signal_16170, new_AGEMA_signal_16169, mcs1_mcs_mat1_4_n100}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U51 ( .a ({new_AGEMA_signal_17035, new_AGEMA_signal_17034, new_AGEMA_signal_17033, mcs1_mcs_mat1_4_n98}), .b ({new_AGEMA_signal_20593, new_AGEMA_signal_20592, new_AGEMA_signal_20591, mcs1_mcs_mat1_4_n97}), .c ({new_AGEMA_signal_21262, new_AGEMA_signal_21261, new_AGEMA_signal_21260, mcs_out[204]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U50 ( .a ({new_AGEMA_signal_19798, new_AGEMA_signal_19797, new_AGEMA_signal_19796, mcs1_mcs_mat1_4_mcs_out[108]}), .b ({new_AGEMA_signal_17749, new_AGEMA_signal_17748, new_AGEMA_signal_17747, mcs1_mcs_mat1_4_mcs_out[96]}), .c ({new_AGEMA_signal_20593, new_AGEMA_signal_20592, new_AGEMA_signal_20591, mcs1_mcs_mat1_4_n97}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U49 ( .a ({new_AGEMA_signal_15046, new_AGEMA_signal_15045, new_AGEMA_signal_15044, mcs1_mcs_mat1_4_mcs_out[100]}), .b ({new_AGEMA_signal_16198, new_AGEMA_signal_16197, new_AGEMA_signal_16196, mcs1_mcs_mat1_4_mcs_out[104]}), .c ({new_AGEMA_signal_17035, new_AGEMA_signal_17034, new_AGEMA_signal_17033, mcs1_mcs_mat1_4_n98}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U48 ( .a ({new_AGEMA_signal_14989, new_AGEMA_signal_14988, new_AGEMA_signal_14987, mcs1_mcs_mat1_4_n96}), .b ({new_AGEMA_signal_19768, new_AGEMA_signal_19767, new_AGEMA_signal_19766, mcs1_mcs_mat1_4_n95}), .c ({new_AGEMA_signal_20596, new_AGEMA_signal_20595, new_AGEMA_signal_20594, mcs_out[175]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U47 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_19072, new_AGEMA_signal_19071, new_AGEMA_signal_19070, mcs1_mcs_mat1_4_mcs_out[95]}), .c ({new_AGEMA_signal_19768, new_AGEMA_signal_19767, new_AGEMA_signal_19766, mcs1_mcs_mat1_4_n95}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U46 ( .a ({new_AGEMA_signal_13597, new_AGEMA_signal_13596, new_AGEMA_signal_13595, mcs1_mcs_mat1_4_mcs_out[83]}), .b ({new_AGEMA_signal_12151, new_AGEMA_signal_12150, new_AGEMA_signal_12149, mcs1_mcs_mat1_4_mcs_out[87]}), .c ({new_AGEMA_signal_14989, new_AGEMA_signal_14988, new_AGEMA_signal_14987, mcs1_mcs_mat1_4_n96}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U45 ( .a ({new_AGEMA_signal_14992, new_AGEMA_signal_14991, new_AGEMA_signal_14990, mcs1_mcs_mat1_4_n94}), .b ({new_AGEMA_signal_18406, new_AGEMA_signal_18405, new_AGEMA_signal_18404, mcs1_mcs_mat1_4_n93}), .c ({new_AGEMA_signal_19051, new_AGEMA_signal_19050, new_AGEMA_signal_19049, mcs_out[174]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U43 ( .a ({new_AGEMA_signal_13600, new_AGEMA_signal_13599, new_AGEMA_signal_13598, mcs1_mcs_mat1_4_mcs_out[82]}), .b ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_14992, new_AGEMA_signal_14991, new_AGEMA_signal_14990, mcs1_mcs_mat1_4_n94}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U42 ( .a ({new_AGEMA_signal_14995, new_AGEMA_signal_14994, new_AGEMA_signal_14993, mcs1_mcs_mat1_4_n92}), .b ({new_AGEMA_signal_18409, new_AGEMA_signal_18408, new_AGEMA_signal_18407, mcs1_mcs_mat1_4_n91}), .c ({new_AGEMA_signal_19054, new_AGEMA_signal_19053, new_AGEMA_signal_19052, mcs_out[173]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U41 ( .a ({new_AGEMA_signal_10957, new_AGEMA_signal_10956, new_AGEMA_signal_10955, mcs1_mcs_mat1_4_mcs_out[89]}), .b ({new_AGEMA_signal_17755, new_AGEMA_signal_17754, new_AGEMA_signal_17753, mcs1_mcs_mat1_4_mcs_out[93]}), .c ({new_AGEMA_signal_18409, new_AGEMA_signal_18408, new_AGEMA_signal_18407, mcs1_mcs_mat1_4_n91}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U40 ( .a ({new_AGEMA_signal_13603, new_AGEMA_signal_13602, new_AGEMA_signal_13601, mcs1_mcs_mat1_4_mcs_out[81]}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_14995, new_AGEMA_signal_14994, new_AGEMA_signal_14993, mcs1_mcs_mat1_4_n92}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U39 ( .a ({new_AGEMA_signal_16174, new_AGEMA_signal_16173, new_AGEMA_signal_16172, mcs1_mcs_mat1_4_n90}), .b ({new_AGEMA_signal_20599, new_AGEMA_signal_20598, new_AGEMA_signal_20597, mcs1_mcs_mat1_4_n89}), .c ({new_AGEMA_signal_21265, new_AGEMA_signal_21264, new_AGEMA_signal_21263, mcs_out[172]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U38 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_19801, new_AGEMA_signal_19800, new_AGEMA_signal_19799, mcs1_mcs_mat1_4_mcs_out[92]}), .c ({new_AGEMA_signal_20599, new_AGEMA_signal_20598, new_AGEMA_signal_20597, mcs1_mcs_mat1_4_n89}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U37 ( .a ({new_AGEMA_signal_15055, new_AGEMA_signal_15054, new_AGEMA_signal_15053, mcs1_mcs_mat1_4_mcs_out[80]}), .b ({new_AGEMA_signal_13594, new_AGEMA_signal_13593, new_AGEMA_signal_13592, mcs1_mcs_mat1_4_mcs_out[84]}), .c ({new_AGEMA_signal_16174, new_AGEMA_signal_16173, new_AGEMA_signal_16172, mcs1_mcs_mat1_4_n90}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U36 ( .a ({new_AGEMA_signal_19771, new_AGEMA_signal_19770, new_AGEMA_signal_19769, mcs1_mcs_mat1_4_n88}), .b ({new_AGEMA_signal_14998, new_AGEMA_signal_14997, new_AGEMA_signal_14996, mcs1_mcs_mat1_4_n87}), .c ({temp_next_s3[13], temp_next_s2[13], temp_next_s1[13], temp_next_s0[13]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U35 ( .a ({new_AGEMA_signal_11017, new_AGEMA_signal_11016, new_AGEMA_signal_11015, mcs1_mcs_mat1_4_mcs_out[5]}), .b ({new_AGEMA_signal_13708, new_AGEMA_signal_13707, new_AGEMA_signal_13706, mcs1_mcs_mat1_4_mcs_out[9]}), .c ({new_AGEMA_signal_14998, new_AGEMA_signal_14997, new_AGEMA_signal_14996, mcs1_mcs_mat1_4_n87}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U34 ( .a ({new_AGEMA_signal_19105, new_AGEMA_signal_19104, new_AGEMA_signal_19103, mcs1_mcs_mat1_4_mcs_out[13]}), .b ({new_AGEMA_signal_15154, new_AGEMA_signal_15153, new_AGEMA_signal_15152, mcs1_mcs_mat1_4_mcs_out[1]}), .c ({new_AGEMA_signal_19771, new_AGEMA_signal_19770, new_AGEMA_signal_19769, mcs1_mcs_mat1_4_n88}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U33 ( .a ({new_AGEMA_signal_17038, new_AGEMA_signal_17037, new_AGEMA_signal_17036, mcs1_mcs_mat1_4_n86}), .b ({new_AGEMA_signal_19774, new_AGEMA_signal_19773, new_AGEMA_signal_19772, mcs1_mcs_mat1_4_n85}), .c ({new_AGEMA_signal_20605, new_AGEMA_signal_20604, new_AGEMA_signal_20603, mcs_out[143]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U32 ( .a ({new_AGEMA_signal_12166, new_AGEMA_signal_12165, new_AGEMA_signal_12164, mcs1_mcs_mat1_4_mcs_out[75]}), .b ({new_AGEMA_signal_19078, new_AGEMA_signal_19077, new_AGEMA_signal_19076, mcs1_mcs_mat1_4_mcs_out[79]}), .c ({new_AGEMA_signal_19774, new_AGEMA_signal_19773, new_AGEMA_signal_19772, mcs1_mcs_mat1_4_n85}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U31 ( .a ({new_AGEMA_signal_16216, new_AGEMA_signal_16215, new_AGEMA_signal_16214, mcs1_mcs_mat1_4_mcs_out[67]}), .b ({new_AGEMA_signal_15070, new_AGEMA_signal_15069, new_AGEMA_signal_15068, mcs1_mcs_mat1_4_mcs_out[71]}), .c ({new_AGEMA_signal_17038, new_AGEMA_signal_17037, new_AGEMA_signal_17036, mcs1_mcs_mat1_4_n86}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U30 ( .a ({new_AGEMA_signal_17044, new_AGEMA_signal_17043, new_AGEMA_signal_17042, mcs1_mcs_mat1_4_n84}), .b ({new_AGEMA_signal_17041, new_AGEMA_signal_17040, new_AGEMA_signal_17039, mcs1_mcs_mat1_4_n83}), .c ({new_AGEMA_signal_17734, new_AGEMA_signal_17733, new_AGEMA_signal_17732, mcs_out[142]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U29 ( .a ({new_AGEMA_signal_16204, new_AGEMA_signal_16203, new_AGEMA_signal_16202, mcs1_mcs_mat1_4_mcs_out[74]}), .b ({new_AGEMA_signal_15058, new_AGEMA_signal_15057, new_AGEMA_signal_15056, mcs1_mcs_mat1_4_mcs_out[78]}), .c ({new_AGEMA_signal_17041, new_AGEMA_signal_17040, new_AGEMA_signal_17039, mcs1_mcs_mat1_4_n83}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U28 ( .a ({new_AGEMA_signal_15079, new_AGEMA_signal_15078, new_AGEMA_signal_15077, mcs1_mcs_mat1_4_mcs_out[66]}), .b ({new_AGEMA_signal_16210, new_AGEMA_signal_16209, new_AGEMA_signal_16208, mcs1_mcs_mat1_4_mcs_out[70]}), .c ({new_AGEMA_signal_17044, new_AGEMA_signal_17043, new_AGEMA_signal_17042, mcs1_mcs_mat1_4_n84}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U27 ( .a ({new_AGEMA_signal_17047, new_AGEMA_signal_17046, new_AGEMA_signal_17045, mcs1_mcs_mat1_4_n82}), .b ({new_AGEMA_signal_18412, new_AGEMA_signal_18411, new_AGEMA_signal_18410, mcs1_mcs_mat1_4_n81}), .c ({new_AGEMA_signal_19057, new_AGEMA_signal_19056, new_AGEMA_signal_19055, mcs_out[141]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U26 ( .a ({new_AGEMA_signal_13612, new_AGEMA_signal_13611, new_AGEMA_signal_13610, mcs1_mcs_mat1_4_mcs_out[73]}), .b ({new_AGEMA_signal_17761, new_AGEMA_signal_17760, new_AGEMA_signal_17759, mcs1_mcs_mat1_4_mcs_out[77]}), .c ({new_AGEMA_signal_18412, new_AGEMA_signal_18411, new_AGEMA_signal_18410, mcs1_mcs_mat1_4_n81}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U25 ( .a ({new_AGEMA_signal_12184, new_AGEMA_signal_12183, new_AGEMA_signal_12182, mcs1_mcs_mat1_4_mcs_out[65]}), .b ({new_AGEMA_signal_16213, new_AGEMA_signal_16212, new_AGEMA_signal_16211, mcs1_mcs_mat1_4_mcs_out[69]}), .c ({new_AGEMA_signal_17047, new_AGEMA_signal_17046, new_AGEMA_signal_17045, mcs1_mcs_mat1_4_n82}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U24 ( .a ({new_AGEMA_signal_17737, new_AGEMA_signal_17736, new_AGEMA_signal_17735, mcs1_mcs_mat1_4_n80}), .b ({new_AGEMA_signal_20608, new_AGEMA_signal_20607, new_AGEMA_signal_20606, mcs1_mcs_mat1_4_n79}), .c ({new_AGEMA_signal_21268, new_AGEMA_signal_21267, new_AGEMA_signal_21266, mcs_out[140]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U23 ( .a ({new_AGEMA_signal_16207, new_AGEMA_signal_16206, new_AGEMA_signal_16205, mcs1_mcs_mat1_4_mcs_out[72]}), .b ({new_AGEMA_signal_19804, new_AGEMA_signal_19803, new_AGEMA_signal_19802, mcs1_mcs_mat1_4_mcs_out[76]}), .c ({new_AGEMA_signal_20608, new_AGEMA_signal_20607, new_AGEMA_signal_20606, mcs1_mcs_mat1_4_n79}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U22 ( .a ({new_AGEMA_signal_17080, new_AGEMA_signal_17079, new_AGEMA_signal_17078, mcs1_mcs_mat1_4_mcs_out[64]}), .b ({new_AGEMA_signal_15076, new_AGEMA_signal_15075, new_AGEMA_signal_15074, mcs1_mcs_mat1_4_mcs_out[68]}), .c ({new_AGEMA_signal_17737, new_AGEMA_signal_17736, new_AGEMA_signal_17735, mcs1_mcs_mat1_4_n80}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U21 ( .a ({new_AGEMA_signal_16177, new_AGEMA_signal_16176, new_AGEMA_signal_16175, mcs1_mcs_mat1_4_n78}), .b ({new_AGEMA_signal_19777, new_AGEMA_signal_19776, new_AGEMA_signal_19775, mcs1_mcs_mat1_4_n77}), .c ({temp_next_s3[111], temp_next_s2[111], temp_next_s1[111], temp_next_s0[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U20 ( .a ({new_AGEMA_signal_13630, new_AGEMA_signal_13629, new_AGEMA_signal_13628, mcs1_mcs_mat1_4_mcs_out[59]}), .b ({new_AGEMA_signal_19084, new_AGEMA_signal_19083, new_AGEMA_signal_19082, mcs1_mcs_mat1_4_mcs_out[63]}), .c ({new_AGEMA_signal_19777, new_AGEMA_signal_19776, new_AGEMA_signal_19775, mcs1_mcs_mat1_4_n77}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U19 ( .a ({new_AGEMA_signal_12214, new_AGEMA_signal_12213, new_AGEMA_signal_12212, mcs1_mcs_mat1_4_mcs_out[51]}), .b ({new_AGEMA_signal_15091, new_AGEMA_signal_15090, new_AGEMA_signal_15089, mcs1_mcs_mat1_4_mcs_out[55]}), .c ({new_AGEMA_signal_16177, new_AGEMA_signal_16176, new_AGEMA_signal_16175, mcs1_mcs_mat1_4_n78}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U18 ( .a ({new_AGEMA_signal_17050, new_AGEMA_signal_17049, new_AGEMA_signal_17048, mcs1_mcs_mat1_4_n76}), .b ({new_AGEMA_signal_19060, new_AGEMA_signal_19059, new_AGEMA_signal_19058, mcs1_mcs_mat1_4_n75}), .c ({temp_next_s3[110], temp_next_s2[110], temp_next_s1[110], temp_next_s0[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U17 ( .a ({new_AGEMA_signal_12190, new_AGEMA_signal_12189, new_AGEMA_signal_12188, mcs1_mcs_mat1_4_mcs_out[58]}), .b ({new_AGEMA_signal_18433, new_AGEMA_signal_18432, new_AGEMA_signal_18431, mcs1_mcs_mat1_4_mcs_out[62]}), .c ({new_AGEMA_signal_19060, new_AGEMA_signal_19059, new_AGEMA_signal_19058, mcs1_mcs_mat1_4_n75}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U16 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_16222, new_AGEMA_signal_16221, new_AGEMA_signal_16220, mcs1_mcs_mat1_4_mcs_out[54]}), .c ({new_AGEMA_signal_17050, new_AGEMA_signal_17049, new_AGEMA_signal_17048, mcs1_mcs_mat1_4_n76}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U15 ( .a ({new_AGEMA_signal_17053, new_AGEMA_signal_17052, new_AGEMA_signal_17051, mcs1_mcs_mat1_4_n74}), .b ({new_AGEMA_signal_19063, new_AGEMA_signal_19062, new_AGEMA_signal_19061, mcs1_mcs_mat1_4_n73}), .c ({temp_next_s3[109], temp_next_s2[109], temp_next_s1[109], temp_next_s0[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U14 ( .a ({new_AGEMA_signal_13633, new_AGEMA_signal_13632, new_AGEMA_signal_13631, mcs1_mcs_mat1_4_mcs_out[57]}), .b ({new_AGEMA_signal_18436, new_AGEMA_signal_18435, new_AGEMA_signal_18434, mcs1_mcs_mat1_4_mcs_out[61]}), .c ({new_AGEMA_signal_19063, new_AGEMA_signal_19062, new_AGEMA_signal_19061, mcs1_mcs_mat1_4_n73}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U13 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({new_AGEMA_signal_16225, new_AGEMA_signal_16224, new_AGEMA_signal_16223, mcs1_mcs_mat1_4_mcs_out[53]}), .c ({new_AGEMA_signal_17053, new_AGEMA_signal_17052, new_AGEMA_signal_17051, mcs1_mcs_mat1_4_n74}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U12 ( .a ({new_AGEMA_signal_16180, new_AGEMA_signal_16179, new_AGEMA_signal_16178, mcs1_mcs_mat1_4_n72}), .b ({new_AGEMA_signal_20614, new_AGEMA_signal_20613, new_AGEMA_signal_20612, mcs1_mcs_mat1_4_n71}), .c ({temp_next_s3[108], temp_next_s2[108], temp_next_s1[108], temp_next_s0[108]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U11 ( .a ({new_AGEMA_signal_15088, new_AGEMA_signal_15087, new_AGEMA_signal_15086, mcs1_mcs_mat1_4_mcs_out[56]}), .b ({new_AGEMA_signal_19807, new_AGEMA_signal_19806, new_AGEMA_signal_19805, mcs1_mcs_mat1_4_mcs_out[60]}), .c ({new_AGEMA_signal_20614, new_AGEMA_signal_20613, new_AGEMA_signal_20612, mcs1_mcs_mat1_4_n71}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U10 ( .a ({new_AGEMA_signal_13645, new_AGEMA_signal_13644, new_AGEMA_signal_13643, mcs1_mcs_mat1_4_mcs_out[48]}), .b ({new_AGEMA_signal_15097, new_AGEMA_signal_15096, new_AGEMA_signal_15095, mcs1_mcs_mat1_4_mcs_out[52]}), .c ({new_AGEMA_signal_16180, new_AGEMA_signal_16179, new_AGEMA_signal_16178, mcs1_mcs_mat1_4_n72}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U9 ( .a ({new_AGEMA_signal_17056, new_AGEMA_signal_17055, new_AGEMA_signal_17054, mcs1_mcs_mat1_4_n70}), .b ({new_AGEMA_signal_19786, new_AGEMA_signal_19785, new_AGEMA_signal_19784, mcs1_mcs_mat1_4_n69}), .c ({temp_next_s3[79], temp_next_s2[79], temp_next_s1[79], temp_next_s0[79]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U8 ( .a ({new_AGEMA_signal_15103, new_AGEMA_signal_15102, new_AGEMA_signal_15101, mcs1_mcs_mat1_4_mcs_out[43]}), .b ({new_AGEMA_signal_19090, new_AGEMA_signal_19089, new_AGEMA_signal_19088, mcs1_mcs_mat1_4_mcs_out[47]}), .c ({new_AGEMA_signal_19786, new_AGEMA_signal_19785, new_AGEMA_signal_19784, mcs1_mcs_mat1_4_n69}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U7 ( .a ({new_AGEMA_signal_15115, new_AGEMA_signal_15114, new_AGEMA_signal_15113, mcs1_mcs_mat1_4_mcs_out[35]}), .b ({new_AGEMA_signal_16228, new_AGEMA_signal_16227, new_AGEMA_signal_16226, mcs1_mcs_mat1_4_mcs_out[39]}), .c ({new_AGEMA_signal_17056, new_AGEMA_signal_17055, new_AGEMA_signal_17054, mcs1_mcs_mat1_4_n70}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U6 ( .a ({new_AGEMA_signal_15001, new_AGEMA_signal_15000, new_AGEMA_signal_14999, mcs1_mcs_mat1_4_n68}), .b ({new_AGEMA_signal_17740, new_AGEMA_signal_17739, new_AGEMA_signal_17738, mcs1_mcs_mat1_4_n67}), .c ({temp_next_s3[78], temp_next_s2[78], temp_next_s1[78], temp_next_s0[78]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U5 ( .a ({new_AGEMA_signal_15106, new_AGEMA_signal_15105, new_AGEMA_signal_15104, mcs1_mcs_mat1_4_mcs_out[42]}), .b ({new_AGEMA_signal_17086, new_AGEMA_signal_17085, new_AGEMA_signal_17084, mcs1_mcs_mat1_4_mcs_out[46]}), .c ({new_AGEMA_signal_17740, new_AGEMA_signal_17739, new_AGEMA_signal_17738, mcs1_mcs_mat1_4_n67}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U4 ( .a ({new_AGEMA_signal_13669, new_AGEMA_signal_13668, new_AGEMA_signal_13667, mcs1_mcs_mat1_4_mcs_out[34]}), .b ({new_AGEMA_signal_12226, new_AGEMA_signal_12225, new_AGEMA_signal_12224, mcs1_mcs_mat1_4_mcs_out[38]}), .c ({new_AGEMA_signal_15001, new_AGEMA_signal_15000, new_AGEMA_signal_14999, mcs1_mcs_mat1_4_n68}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U3 ( .a ({new_AGEMA_signal_21274, new_AGEMA_signal_21273, new_AGEMA_signal_21272, mcs1_mcs_mat1_4_n66}), .b ({new_AGEMA_signal_18418, new_AGEMA_signal_18417, new_AGEMA_signal_18416, mcs1_mcs_mat1_4_n65}), .c ({temp_next_s3[12], temp_next_s2[12], temp_next_s1[12], temp_next_s0[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U2 ( .a ({new_AGEMA_signal_17794, new_AGEMA_signal_17793, new_AGEMA_signal_17792, mcs1_mcs_mat1_4_mcs_out[4]}), .b ({new_AGEMA_signal_16249, new_AGEMA_signal_16248, new_AGEMA_signal_16247, mcs1_mcs_mat1_4_mcs_out[8]}), .c ({new_AGEMA_signal_18418, new_AGEMA_signal_18417, new_AGEMA_signal_18416, mcs1_mcs_mat1_4_n65}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_U1 ( .a ({new_AGEMA_signal_15157, new_AGEMA_signal_15156, new_AGEMA_signal_15155, mcs1_mcs_mat1_4_mcs_out[0]}), .b ({new_AGEMA_signal_20623, new_AGEMA_signal_20622, new_AGEMA_signal_20621, mcs1_mcs_mat1_4_mcs_out[12]}), .c ({new_AGEMA_signal_21274, new_AGEMA_signal_21273, new_AGEMA_signal_21272, mcs1_mcs_mat1_4_n66}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_15004, new_AGEMA_signal_15003, new_AGEMA_signal_15002, mcs1_mcs_mat1_4_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_16183, new_AGEMA_signal_16182, new_AGEMA_signal_16181, mcs1_mcs_mat1_4_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_13549, new_AGEMA_signal_13548, new_AGEMA_signal_13547, mcs1_mcs_mat1_4_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_8890, new_AGEMA_signal_8889, new_AGEMA_signal_8888, mcs1_mcs_mat1_4_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_15004, new_AGEMA_signal_15003, new_AGEMA_signal_15002, mcs1_mcs_mat1_4_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_9727, new_AGEMA_signal_9726, new_AGEMA_signal_9725, mcs1_mcs_mat1_4_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_10915, new_AGEMA_signal_10914, new_AGEMA_signal_10913, mcs1_mcs_mat1_4_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_12106, new_AGEMA_signal_12105, new_AGEMA_signal_12104, mcs1_mcs_mat1_4_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_9730, new_AGEMA_signal_9729, new_AGEMA_signal_9728, mcs1_mcs_mat1_4_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .c ({new_AGEMA_signal_10915, new_AGEMA_signal_10914, new_AGEMA_signal_10913, mcs1_mcs_mat1_4_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_15007, new_AGEMA_signal_15006, new_AGEMA_signal_15005, mcs1_mcs_mat1_4_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .c ({new_AGEMA_signal_16186, new_AGEMA_signal_16185, new_AGEMA_signal_16184, mcs1_mcs_mat1_4_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_13549, new_AGEMA_signal_13548, new_AGEMA_signal_13547, mcs1_mcs_mat1_4_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_15007, new_AGEMA_signal_15006, new_AGEMA_signal_15005, mcs1_mcs_mat1_4_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_12109, new_AGEMA_signal_12108, new_AGEMA_signal_12107, mcs1_mcs_mat1_4_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_10918, new_AGEMA_signal_10917, new_AGEMA_signal_10916, mcs1_mcs_mat1_4_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_13549, new_AGEMA_signal_13548, new_AGEMA_signal_13547, mcs1_mcs_mat1_4_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_13552, new_AGEMA_signal_13551, new_AGEMA_signal_13550, mcs1_mcs_mat1_4_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_15010, new_AGEMA_signal_15009, new_AGEMA_signal_15008, mcs1_mcs_mat1_4_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_12109, new_AGEMA_signal_12108, new_AGEMA_signal_12107, mcs1_mcs_mat1_4_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9730, new_AGEMA_signal_9729, new_AGEMA_signal_9728, mcs1_mcs_mat1_4_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_13552, new_AGEMA_signal_13551, new_AGEMA_signal_13550, mcs1_mcs_mat1_4_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704]}), .c ({new_AGEMA_signal_12109, new_AGEMA_signal_12108, new_AGEMA_signal_12107, mcs1_mcs_mat1_4_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710]}), .c ({new_AGEMA_signal_9730, new_AGEMA_signal_9729, new_AGEMA_signal_9728, mcs1_mcs_mat1_4_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4721], Fresh[4720], Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716]}), .c ({new_AGEMA_signal_10918, new_AGEMA_signal_10917, new_AGEMA_signal_10916, mcs1_mcs_mat1_4_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_15013, new_AGEMA_signal_15012, new_AGEMA_signal_15011, mcs1_mcs_mat1_4_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .c ({new_AGEMA_signal_16189, new_AGEMA_signal_16188, new_AGEMA_signal_16187, mcs1_mcs_mat1_4_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_13555, new_AGEMA_signal_13554, new_AGEMA_signal_13553, mcs1_mcs_mat1_4_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10927, new_AGEMA_signal_10926, new_AGEMA_signal_10925, mcs1_mcs_mat1_4_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_15013, new_AGEMA_signal_15012, new_AGEMA_signal_15011, mcs1_mcs_mat1_4_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_15016, new_AGEMA_signal_15015, new_AGEMA_signal_15014, mcs1_mcs_mat1_4_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_12115, new_AGEMA_signal_12114, new_AGEMA_signal_12113, mcs1_mcs_mat1_4_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_16192, new_AGEMA_signal_16191, new_AGEMA_signal_16190, mcs1_mcs_mat1_4_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_13555, new_AGEMA_signal_13554, new_AGEMA_signal_13553, mcs1_mcs_mat1_4_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .c ({new_AGEMA_signal_15016, new_AGEMA_signal_15015, new_AGEMA_signal_15014, mcs1_mcs_mat1_4_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_13555, new_AGEMA_signal_13554, new_AGEMA_signal_13553, mcs1_mcs_mat1_4_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_12112, new_AGEMA_signal_12111, new_AGEMA_signal_12110, mcs1_mcs_mat1_4_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_15019, new_AGEMA_signal_15018, new_AGEMA_signal_15017, mcs1_mcs_mat1_4_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_12118, new_AGEMA_signal_12117, new_AGEMA_signal_12116, mcs1_mcs_mat1_4_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_9733, new_AGEMA_signal_9732, new_AGEMA_signal_9731, mcs1_mcs_mat1_4_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_13555, new_AGEMA_signal_13554, new_AGEMA_signal_13553, mcs1_mcs_mat1_4_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_10924, new_AGEMA_signal_10923, new_AGEMA_signal_10922, mcs1_mcs_mat1_4_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_12115, new_AGEMA_signal_12114, new_AGEMA_signal_12113, mcs1_mcs_mat1_4_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_13558, new_AGEMA_signal_13557, new_AGEMA_signal_13556, mcs1_mcs_mat1_4_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_8893, new_AGEMA_signal_8892, new_AGEMA_signal_8891, mcs1_mcs_mat1_4_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_10927, new_AGEMA_signal_10926, new_AGEMA_signal_10925, mcs1_mcs_mat1_4_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_12115, new_AGEMA_signal_12114, new_AGEMA_signal_12113, mcs1_mcs_mat1_4_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_9733, new_AGEMA_signal_9732, new_AGEMA_signal_9731, mcs1_mcs_mat1_4_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_10924, new_AGEMA_signal_10923, new_AGEMA_signal_10922, mcs1_mcs_mat1_4_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4727], Fresh[4726], Fresh[4725], Fresh[4724], Fresh[4723], Fresh[4722]}), .c ({new_AGEMA_signal_12118, new_AGEMA_signal_12117, new_AGEMA_signal_12116, mcs1_mcs_mat1_4_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730], Fresh[4729], Fresh[4728]}), .c ({new_AGEMA_signal_9733, new_AGEMA_signal_9732, new_AGEMA_signal_9731, mcs1_mcs_mat1_4_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734]}), .c ({new_AGEMA_signal_10927, new_AGEMA_signal_10926, new_AGEMA_signal_10925, mcs1_mcs_mat1_4_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_13564, new_AGEMA_signal_13563, new_AGEMA_signal_13562, mcs1_mcs_mat1_4_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_9736, new_AGEMA_signal_9735, new_AGEMA_signal_9734, mcs1_mcs_mat1_4_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_15022, new_AGEMA_signal_15021, new_AGEMA_signal_15020, mcs1_mcs_mat1_4_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_10930, new_AGEMA_signal_10929, new_AGEMA_signal_10928, mcs1_mcs_mat1_4_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_10933, new_AGEMA_signal_10932, new_AGEMA_signal_10931, mcs1_mcs_mat1_4_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_12121, new_AGEMA_signal_12120, new_AGEMA_signal_12119, mcs1_mcs_mat1_4_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_13567, new_AGEMA_signal_13566, new_AGEMA_signal_13565, mcs1_mcs_mat1_4_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_15025, new_AGEMA_signal_15024, new_AGEMA_signal_15023, mcs1_mcs_mat1_4_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_16195, new_AGEMA_signal_16194, new_AGEMA_signal_16193, mcs1_mcs_mat1_4_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_13564, new_AGEMA_signal_13563, new_AGEMA_signal_13562, mcs1_mcs_mat1_4_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_15025, new_AGEMA_signal_15024, new_AGEMA_signal_15023, mcs1_mcs_mat1_4_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_8896, new_AGEMA_signal_8895, new_AGEMA_signal_8894, mcs1_mcs_mat1_4_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_12127, new_AGEMA_signal_12126, new_AGEMA_signal_12125, mcs1_mcs_mat1_4_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_13564, new_AGEMA_signal_13563, new_AGEMA_signal_13562, mcs1_mcs_mat1_4_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_9739, new_AGEMA_signal_9738, new_AGEMA_signal_9737, mcs1_mcs_mat1_4_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_12124, new_AGEMA_signal_12123, new_AGEMA_signal_12122, mcs1_mcs_mat1_4_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_13567, new_AGEMA_signal_13566, new_AGEMA_signal_13565, mcs1_mcs_mat1_4_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740]}), .c ({new_AGEMA_signal_12127, new_AGEMA_signal_12126, new_AGEMA_signal_12125, mcs1_mcs_mat1_4_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4751], Fresh[4750], Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746]}), .c ({new_AGEMA_signal_9739, new_AGEMA_signal_9738, new_AGEMA_signal_9737, mcs1_mcs_mat1_4_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4757], Fresh[4756], Fresh[4755], Fresh[4754], Fresh[4753], Fresh[4752]}), .c ({new_AGEMA_signal_10933, new_AGEMA_signal_10932, new_AGEMA_signal_10931, mcs1_mcs_mat1_4_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({new_AGEMA_signal_19066, new_AGEMA_signal_19065, new_AGEMA_signal_19064, mcs1_mcs_mat1_4_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_19789, new_AGEMA_signal_19788, new_AGEMA_signal_19787, mcs1_mcs_mat1_4_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({new_AGEMA_signal_19069, new_AGEMA_signal_19068, new_AGEMA_signal_19067, mcs1_mcs_mat1_4_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_19792, new_AGEMA_signal_19791, new_AGEMA_signal_19790, mcs1_mcs_mat1_4_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_17062, new_AGEMA_signal_17061, new_AGEMA_signal_17060, mcs1_mcs_mat1_4_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_19066, new_AGEMA_signal_19065, new_AGEMA_signal_19064, mcs1_mcs_mat1_4_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_19795, new_AGEMA_signal_19794, new_AGEMA_signal_19793, mcs1_mcs_mat1_4_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_15028, new_AGEMA_signal_15027, new_AGEMA_signal_15026, mcs1_mcs_mat1_4_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_18421, new_AGEMA_signal_18420, new_AGEMA_signal_18419, mcs1_mcs_mat1_4_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_19066, new_AGEMA_signal_19065, new_AGEMA_signal_19064, mcs1_mcs_mat1_4_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_17743, new_AGEMA_signal_17742, new_AGEMA_signal_17741, mcs1_mcs_mat1_4_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_19069, new_AGEMA_signal_19068, new_AGEMA_signal_19067, mcs1_mcs_mat1_4_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_19798, new_AGEMA_signal_19797, new_AGEMA_signal_19796, mcs1_mcs_mat1_4_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_18424, new_AGEMA_signal_18423, new_AGEMA_signal_18422, mcs1_mcs_mat1_4_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_19069, new_AGEMA_signal_19068, new_AGEMA_signal_19067, mcs1_mcs_mat1_4_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_17062, new_AGEMA_signal_17061, new_AGEMA_signal_17060, mcs1_mcs_mat1_4_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_17746, new_AGEMA_signal_17745, new_AGEMA_signal_17744, mcs1_mcs_mat1_4_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_18424, new_AGEMA_signal_18423, new_AGEMA_signal_18422, mcs1_mcs_mat1_4_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760], Fresh[4759], Fresh[4758]}), .c ({new_AGEMA_signal_17746, new_AGEMA_signal_17745, new_AGEMA_signal_17744, mcs1_mcs_mat1_4_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764]}), .c ({new_AGEMA_signal_15028, new_AGEMA_signal_15027, new_AGEMA_signal_15026, mcs1_mcs_mat1_4_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770]}), .c ({new_AGEMA_signal_17062, new_AGEMA_signal_17061, new_AGEMA_signal_17060, mcs1_mcs_mat1_4_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_13576, new_AGEMA_signal_13575, new_AGEMA_signal_13574, mcs1_mcs_mat1_4_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_13573, new_AGEMA_signal_13572, new_AGEMA_signal_13571, mcs1_mcs_mat1_4_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_15031, new_AGEMA_signal_15030, new_AGEMA_signal_15029, mcs1_mcs_mat1_4_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_13573, new_AGEMA_signal_13572, new_AGEMA_signal_13571, mcs1_mcs_mat1_4_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_10936, new_AGEMA_signal_10935, new_AGEMA_signal_10934, mcs1_mcs_mat1_4_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_15034, new_AGEMA_signal_15033, new_AGEMA_signal_15032, mcs1_mcs_mat1_4_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_9742, new_AGEMA_signal_9741, new_AGEMA_signal_9740, mcs1_mcs_mat1_4_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .c ({new_AGEMA_signal_10936, new_AGEMA_signal_10935, new_AGEMA_signal_10934, mcs1_mcs_mat1_4_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({new_AGEMA_signal_13573, new_AGEMA_signal_13572, new_AGEMA_signal_13571, mcs1_mcs_mat1_4_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_15037, new_AGEMA_signal_15036, new_AGEMA_signal_15035, mcs1_mcs_mat1_4_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_12133, new_AGEMA_signal_12132, new_AGEMA_signal_12131, mcs1_mcs_mat1_4_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_8899, new_AGEMA_signal_8898, new_AGEMA_signal_8897, mcs1_mcs_mat1_4_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_13573, new_AGEMA_signal_13572, new_AGEMA_signal_13571, mcs1_mcs_mat1_4_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_15040, new_AGEMA_signal_15039, new_AGEMA_signal_15038, mcs1_mcs_mat1_4_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_16198, new_AGEMA_signal_16197, new_AGEMA_signal_16196, mcs1_mcs_mat1_4_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_13576, new_AGEMA_signal_13575, new_AGEMA_signal_13574, mcs1_mcs_mat1_4_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_12133, new_AGEMA_signal_12132, new_AGEMA_signal_12131, mcs1_mcs_mat1_4_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_15040, new_AGEMA_signal_15039, new_AGEMA_signal_15038, mcs1_mcs_mat1_4_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_12130, new_AGEMA_signal_12129, new_AGEMA_signal_12128, mcs1_mcs_mat1_4_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .c ({new_AGEMA_signal_13576, new_AGEMA_signal_13575, new_AGEMA_signal_13574, mcs1_mcs_mat1_4_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_9742, new_AGEMA_signal_9741, new_AGEMA_signal_9740, mcs1_mcs_mat1_4_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_10939, new_AGEMA_signal_10938, new_AGEMA_signal_10937, mcs1_mcs_mat1_4_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_12130, new_AGEMA_signal_12129, new_AGEMA_signal_12128, mcs1_mcs_mat1_4_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4781], Fresh[4780], Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776]}), .c ({new_AGEMA_signal_12133, new_AGEMA_signal_12132, new_AGEMA_signal_12131, mcs1_mcs_mat1_4_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4787], Fresh[4786], Fresh[4785], Fresh[4784], Fresh[4783], Fresh[4782]}), .c ({new_AGEMA_signal_9742, new_AGEMA_signal_9741, new_AGEMA_signal_9740, mcs1_mcs_mat1_4_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790], Fresh[4789], Fresh[4788]}), .c ({new_AGEMA_signal_10939, new_AGEMA_signal_10938, new_AGEMA_signal_10937, mcs1_mcs_mat1_4_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_10942, new_AGEMA_signal_10941, new_AGEMA_signal_10940, mcs1_mcs_mat1_4_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_13579, new_AGEMA_signal_13578, new_AGEMA_signal_13577, mcs1_mcs_mat1_4_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_15043, new_AGEMA_signal_15042, new_AGEMA_signal_15041, mcs1_mcs_mat1_4_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_12145, new_AGEMA_signal_12144, new_AGEMA_signal_12143, mcs1_mcs_mat1_4_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_13579, new_AGEMA_signal_13578, new_AGEMA_signal_13577, mcs1_mcs_mat1_4_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_12139, new_AGEMA_signal_12138, new_AGEMA_signal_12137, mcs1_mcs_mat1_4_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_10945, new_AGEMA_signal_10944, new_AGEMA_signal_10943, mcs1_mcs_mat1_4_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_13582, new_AGEMA_signal_13581, new_AGEMA_signal_13580, mcs1_mcs_mat1_4_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_12142, new_AGEMA_signal_12141, new_AGEMA_signal_12140, mcs1_mcs_mat1_4_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_13585, new_AGEMA_signal_13584, new_AGEMA_signal_13583, mcs1_mcs_mat1_4_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_15046, new_AGEMA_signal_15045, new_AGEMA_signal_15044, mcs1_mcs_mat1_4_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_8902, new_AGEMA_signal_8901, new_AGEMA_signal_8900, mcs1_mcs_mat1_4_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_12145, new_AGEMA_signal_12144, new_AGEMA_signal_12143, mcs1_mcs_mat1_4_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_13585, new_AGEMA_signal_13584, new_AGEMA_signal_13583, mcs1_mcs_mat1_4_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_9745, new_AGEMA_signal_9744, new_AGEMA_signal_9743, mcs1_mcs_mat1_4_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .c ({new_AGEMA_signal_12142, new_AGEMA_signal_12141, new_AGEMA_signal_12140, mcs1_mcs_mat1_4_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794]}), .c ({new_AGEMA_signal_12145, new_AGEMA_signal_12144, new_AGEMA_signal_12143, mcs1_mcs_mat1_4_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800]}), .c ({new_AGEMA_signal_9745, new_AGEMA_signal_9744, new_AGEMA_signal_9743, mcs1_mcs_mat1_4_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4811], Fresh[4810], Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806]}), .c ({new_AGEMA_signal_10945, new_AGEMA_signal_10944, new_AGEMA_signal_10943, mcs1_mcs_mat1_4_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_17065, new_AGEMA_signal_17064, new_AGEMA_signal_17063, mcs1_mcs_mat1_4_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_10951, new_AGEMA_signal_10950, new_AGEMA_signal_10949, mcs1_mcs_mat1_4_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_17749, new_AGEMA_signal_17748, new_AGEMA_signal_17747, mcs1_mcs_mat1_4_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_16201, new_AGEMA_signal_16200, new_AGEMA_signal_16199, mcs1_mcs_mat1_4_mcs_out[99]}), .b ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .c ({new_AGEMA_signal_17065, new_AGEMA_signal_17064, new_AGEMA_signal_17063, mcs1_mcs_mat1_4_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_15049, new_AGEMA_signal_15048, new_AGEMA_signal_15047, mcs1_mcs_mat1_4_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .c ({new_AGEMA_signal_16201, new_AGEMA_signal_16200, new_AGEMA_signal_16199, mcs1_mcs_mat1_4_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_13588, new_AGEMA_signal_13587, new_AGEMA_signal_13586, mcs1_mcs_mat1_4_mcs_out[98]}), .b ({new_AGEMA_signal_9751, new_AGEMA_signal_9750, new_AGEMA_signal_9749, mcs1_mcs_mat1_4_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_15049, new_AGEMA_signal_15048, new_AGEMA_signal_15047, mcs1_mcs_mat1_4_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_9748, new_AGEMA_signal_9747, new_AGEMA_signal_9746, mcs1_mcs_mat1_4_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_12148, new_AGEMA_signal_12147, new_AGEMA_signal_12146, mcs1_mcs_mat1_4_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_13588, new_AGEMA_signal_13587, new_AGEMA_signal_13586, mcs1_mcs_mat1_4_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4817], Fresh[4816], Fresh[4815], Fresh[4814], Fresh[4813], Fresh[4812]}), .c ({new_AGEMA_signal_12148, new_AGEMA_signal_12147, new_AGEMA_signal_12146, mcs1_mcs_mat1_4_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820], Fresh[4819], Fresh[4818]}), .c ({new_AGEMA_signal_9751, new_AGEMA_signal_9750, new_AGEMA_signal_9749, mcs1_mcs_mat1_4_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824]}), .c ({new_AGEMA_signal_10951, new_AGEMA_signal_10950, new_AGEMA_signal_10949, mcs1_mcs_mat1_4_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_18427, new_AGEMA_signal_18426, new_AGEMA_signal_18425, mcs1_mcs_mat1_4_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_19072, new_AGEMA_signal_19071, new_AGEMA_signal_19070, mcs1_mcs_mat1_4_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_17071, new_AGEMA_signal_17070, new_AGEMA_signal_17069, mcs1_mcs_mat1_4_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_17074, new_AGEMA_signal_17073, new_AGEMA_signal_17072, mcs1_mcs_mat1_4_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_17755, new_AGEMA_signal_17754, new_AGEMA_signal_17753, mcs1_mcs_mat1_4_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_19075, new_AGEMA_signal_19074, new_AGEMA_signal_19073, mcs1_mcs_mat1_4_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_15052, new_AGEMA_signal_15051, new_AGEMA_signal_15050, mcs1_mcs_mat1_4_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_19801, new_AGEMA_signal_19800, new_AGEMA_signal_19799, mcs1_mcs_mat1_4_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_18427, new_AGEMA_signal_18426, new_AGEMA_signal_18425, mcs1_mcs_mat1_4_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .c ({new_AGEMA_signal_19075, new_AGEMA_signal_19074, new_AGEMA_signal_19073, mcs1_mcs_mat1_4_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_13591, new_AGEMA_signal_13590, new_AGEMA_signal_13589, mcs1_mcs_mat1_4_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_17758, new_AGEMA_signal_17757, new_AGEMA_signal_17756, mcs1_mcs_mat1_4_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_18427, new_AGEMA_signal_18426, new_AGEMA_signal_18425, mcs1_mcs_mat1_4_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830]}), .c ({new_AGEMA_signal_17758, new_AGEMA_signal_17757, new_AGEMA_signal_17756, mcs1_mcs_mat1_4_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4841], Fresh[4840], Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836]}), .c ({new_AGEMA_signal_15052, new_AGEMA_signal_15051, new_AGEMA_signal_15050, mcs1_mcs_mat1_4_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4847], Fresh[4846], Fresh[4845], Fresh[4844], Fresh[4843], Fresh[4842]}), .c ({new_AGEMA_signal_17074, new_AGEMA_signal_17073, new_AGEMA_signal_17072, mcs1_mcs_mat1_4_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_12160, new_AGEMA_signal_12159, new_AGEMA_signal_12158, mcs1_mcs_mat1_4_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_12163, new_AGEMA_signal_12162, new_AGEMA_signal_12161, mcs1_mcs_mat1_4_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_13597, new_AGEMA_signal_13596, new_AGEMA_signal_13595, mcs1_mcs_mat1_4_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_12154, new_AGEMA_signal_12153, new_AGEMA_signal_12152, mcs1_mcs_mat1_4_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_8908, new_AGEMA_signal_8907, new_AGEMA_signal_8906, mcs1_mcs_mat1_4_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_13600, new_AGEMA_signal_13599, new_AGEMA_signal_13598, mcs1_mcs_mat1_4_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_10960, new_AGEMA_signal_10959, new_AGEMA_signal_10958, mcs1_mcs_mat1_4_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_12154, new_AGEMA_signal_12153, new_AGEMA_signal_12152, mcs1_mcs_mat1_4_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_12157, new_AGEMA_signal_12156, new_AGEMA_signal_12155, mcs1_mcs_mat1_4_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_13603, new_AGEMA_signal_13602, new_AGEMA_signal_13601, mcs1_mcs_mat1_4_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_9754, new_AGEMA_signal_9753, new_AGEMA_signal_9752, mcs1_mcs_mat1_4_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_10960, new_AGEMA_signal_10959, new_AGEMA_signal_10958, mcs1_mcs_mat1_4_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_12157, new_AGEMA_signal_12156, new_AGEMA_signal_12155, mcs1_mcs_mat1_4_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_13606, new_AGEMA_signal_13605, new_AGEMA_signal_13604, mcs1_mcs_mat1_4_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .c ({new_AGEMA_signal_15055, new_AGEMA_signal_15054, new_AGEMA_signal_15053, mcs1_mcs_mat1_4_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_12160, new_AGEMA_signal_12159, new_AGEMA_signal_12158, mcs1_mcs_mat1_4_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_9754, new_AGEMA_signal_9753, new_AGEMA_signal_9752, mcs1_mcs_mat1_4_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_13606, new_AGEMA_signal_13605, new_AGEMA_signal_13604, mcs1_mcs_mat1_4_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850], Fresh[4849], Fresh[4848]}), .c ({new_AGEMA_signal_12163, new_AGEMA_signal_12162, new_AGEMA_signal_12161, mcs1_mcs_mat1_4_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854]}), .c ({new_AGEMA_signal_9754, new_AGEMA_signal_9753, new_AGEMA_signal_9752, mcs1_mcs_mat1_4_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860]}), .c ({new_AGEMA_signal_10960, new_AGEMA_signal_10959, new_AGEMA_signal_10958, mcs1_mcs_mat1_4_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_18430, new_AGEMA_signal_18429, new_AGEMA_signal_18428, mcs1_mcs_mat1_4_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_19078, new_AGEMA_signal_19077, new_AGEMA_signal_19076, mcs1_mcs_mat1_4_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_17077, new_AGEMA_signal_17076, new_AGEMA_signal_17075, mcs1_mcs_mat1_4_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_17761, new_AGEMA_signal_17760, new_AGEMA_signal_17759, mcs1_mcs_mat1_4_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_19081, new_AGEMA_signal_19080, new_AGEMA_signal_19079, mcs1_mcs_mat1_4_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_15061, new_AGEMA_signal_15060, new_AGEMA_signal_15059, mcs1_mcs_mat1_4_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_19804, new_AGEMA_signal_19803, new_AGEMA_signal_19802, mcs1_mcs_mat1_4_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_18430, new_AGEMA_signal_18429, new_AGEMA_signal_18428, mcs1_mcs_mat1_4_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .c ({new_AGEMA_signal_19081, new_AGEMA_signal_19080, new_AGEMA_signal_19079, mcs1_mcs_mat1_4_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_13609, new_AGEMA_signal_13608, new_AGEMA_signal_13607, mcs1_mcs_mat1_4_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_17764, new_AGEMA_signal_17763, new_AGEMA_signal_17762, mcs1_mcs_mat1_4_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_18430, new_AGEMA_signal_18429, new_AGEMA_signal_18428, mcs1_mcs_mat1_4_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4871], Fresh[4870], Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866]}), .c ({new_AGEMA_signal_17764, new_AGEMA_signal_17763, new_AGEMA_signal_17762, mcs1_mcs_mat1_4_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4877], Fresh[4876], Fresh[4875], Fresh[4874], Fresh[4873], Fresh[4872]}), .c ({new_AGEMA_signal_15061, new_AGEMA_signal_15060, new_AGEMA_signal_15059, mcs1_mcs_mat1_4_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880], Fresh[4879], Fresh[4878]}), .c ({new_AGEMA_signal_17077, new_AGEMA_signal_17076, new_AGEMA_signal_17075, mcs1_mcs_mat1_4_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_15064, new_AGEMA_signal_15063, new_AGEMA_signal_15062, mcs1_mcs_mat1_4_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_16204, new_AGEMA_signal_16203, new_AGEMA_signal_16202, mcs1_mcs_mat1_4_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_13615, new_AGEMA_signal_13614, new_AGEMA_signal_13613, mcs1_mcs_mat1_4_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_12169, new_AGEMA_signal_12168, new_AGEMA_signal_12167, mcs1_mcs_mat1_4_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_15064, new_AGEMA_signal_15063, new_AGEMA_signal_15062, mcs1_mcs_mat1_4_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({new_AGEMA_signal_10321, new_AGEMA_signal_10320, new_AGEMA_signal_10319, mcs1_mcs_mat1_4_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_12166, new_AGEMA_signal_12165, new_AGEMA_signal_12164, mcs1_mcs_mat1_4_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_12169, new_AGEMA_signal_12168, new_AGEMA_signal_12167, mcs1_mcs_mat1_4_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_10321, new_AGEMA_signal_10320, new_AGEMA_signal_10319, mcs1_mcs_mat1_4_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_13612, new_AGEMA_signal_13611, new_AGEMA_signal_13610, mcs1_mcs_mat1_4_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_9757, new_AGEMA_signal_9756, new_AGEMA_signal_9755, mcs1_mcs_mat1_4_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_9760, new_AGEMA_signal_9759, new_AGEMA_signal_9758, mcs1_mcs_mat1_4_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_10321, new_AGEMA_signal_10320, new_AGEMA_signal_10319, mcs1_mcs_mat1_4_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_10963, new_AGEMA_signal_10962, new_AGEMA_signal_10961, mcs1_mcs_mat1_4_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .c ({new_AGEMA_signal_12169, new_AGEMA_signal_12168, new_AGEMA_signal_12167, mcs1_mcs_mat1_4_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_15067, new_AGEMA_signal_15066, new_AGEMA_signal_15065, mcs1_mcs_mat1_4_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_9757, new_AGEMA_signal_9756, new_AGEMA_signal_9755, mcs1_mcs_mat1_4_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_16207, new_AGEMA_signal_16206, new_AGEMA_signal_16205, mcs1_mcs_mat1_4_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_13615, new_AGEMA_signal_13614, new_AGEMA_signal_13613, mcs1_mcs_mat1_4_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_10963, new_AGEMA_signal_10962, new_AGEMA_signal_10961, mcs1_mcs_mat1_4_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_15067, new_AGEMA_signal_15066, new_AGEMA_signal_15065, mcs1_mcs_mat1_4_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .b ({new_AGEMA_signal_12172, new_AGEMA_signal_12171, new_AGEMA_signal_12170, mcs1_mcs_mat1_4_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_13615, new_AGEMA_signal_13614, new_AGEMA_signal_13613, mcs1_mcs_mat1_4_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884]}), .c ({new_AGEMA_signal_12172, new_AGEMA_signal_12171, new_AGEMA_signal_12170, mcs1_mcs_mat1_4_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890]}), .c ({new_AGEMA_signal_9760, new_AGEMA_signal_9759, new_AGEMA_signal_9758, mcs1_mcs_mat1_4_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4901], Fresh[4900], Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896]}), .c ({new_AGEMA_signal_10963, new_AGEMA_signal_10962, new_AGEMA_signal_10961, mcs1_mcs_mat1_4_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_13618, new_AGEMA_signal_13617, new_AGEMA_signal_13616, mcs1_mcs_mat1_4_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_10966, new_AGEMA_signal_10965, new_AGEMA_signal_10964, mcs1_mcs_mat1_4_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_15070, new_AGEMA_signal_15069, new_AGEMA_signal_15068, mcs1_mcs_mat1_4_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_12178, new_AGEMA_signal_12177, new_AGEMA_signal_12176, mcs1_mcs_mat1_4_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_15073, new_AGEMA_signal_15072, new_AGEMA_signal_15071, mcs1_mcs_mat1_4_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_16210, new_AGEMA_signal_16209, new_AGEMA_signal_16208, mcs1_mcs_mat1_4_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_13618, new_AGEMA_signal_13617, new_AGEMA_signal_13616, mcs1_mcs_mat1_4_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_15073, new_AGEMA_signal_15072, new_AGEMA_signal_15071, mcs1_mcs_mat1_4_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_16213, new_AGEMA_signal_16212, new_AGEMA_signal_16211, mcs1_mcs_mat1_4_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_10966, new_AGEMA_signal_10965, new_AGEMA_signal_10964, mcs1_mcs_mat1_4_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_13621, new_AGEMA_signal_13620, new_AGEMA_signal_13619, mcs1_mcs_mat1_4_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_15073, new_AGEMA_signal_15072, new_AGEMA_signal_15071, mcs1_mcs_mat1_4_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({new_AGEMA_signal_9763, new_AGEMA_signal_9762, new_AGEMA_signal_9761, mcs1_mcs_mat1_4_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_10966, new_AGEMA_signal_10965, new_AGEMA_signal_10964, mcs1_mcs_mat1_4_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_12175, new_AGEMA_signal_12174, new_AGEMA_signal_12173, mcs1_mcs_mat1_4_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .c ({new_AGEMA_signal_13618, new_AGEMA_signal_13617, new_AGEMA_signal_13616, mcs1_mcs_mat1_4_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_10969, new_AGEMA_signal_10968, new_AGEMA_signal_10967, mcs1_mcs_mat1_4_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8914, new_AGEMA_signal_8913, new_AGEMA_signal_8912, mcs1_mcs_mat1_4_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_12175, new_AGEMA_signal_12174, new_AGEMA_signal_12173, mcs1_mcs_mat1_4_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_13621, new_AGEMA_signal_13620, new_AGEMA_signal_13619, mcs1_mcs_mat1_4_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_12178, new_AGEMA_signal_12177, new_AGEMA_signal_12176, mcs1_mcs_mat1_4_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_15076, new_AGEMA_signal_15075, new_AGEMA_signal_15074, mcs1_mcs_mat1_4_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_10969, new_AGEMA_signal_10968, new_AGEMA_signal_10967, mcs1_mcs_mat1_4_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_12178, new_AGEMA_signal_12177, new_AGEMA_signal_12176, mcs1_mcs_mat1_4_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({new_AGEMA_signal_12181, new_AGEMA_signal_12180, new_AGEMA_signal_12179, mcs1_mcs_mat1_4_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_13621, new_AGEMA_signal_13620, new_AGEMA_signal_13619, mcs1_mcs_mat1_4_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4907], Fresh[4906], Fresh[4905], Fresh[4904], Fresh[4903], Fresh[4902]}), .c ({new_AGEMA_signal_12181, new_AGEMA_signal_12180, new_AGEMA_signal_12179, mcs1_mcs_mat1_4_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910], Fresh[4909], Fresh[4908]}), .c ({new_AGEMA_signal_9763, new_AGEMA_signal_9762, new_AGEMA_signal_9761, mcs1_mcs_mat1_4_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914]}), .c ({new_AGEMA_signal_10969, new_AGEMA_signal_10968, new_AGEMA_signal_10967, mcs1_mcs_mat1_4_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_15082, new_AGEMA_signal_15081, new_AGEMA_signal_15080, mcs1_mcs_mat1_4_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .c ({new_AGEMA_signal_16216, new_AGEMA_signal_16215, new_AGEMA_signal_16214, mcs1_mcs_mat1_4_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({new_AGEMA_signal_13624, new_AGEMA_signal_13623, new_AGEMA_signal_13622, mcs1_mcs_mat1_4_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_15079, new_AGEMA_signal_15078, new_AGEMA_signal_15077, mcs1_mcs_mat1_4_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_16219, new_AGEMA_signal_16218, new_AGEMA_signal_16217, mcs1_mcs_mat1_4_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_10972, new_AGEMA_signal_10971, new_AGEMA_signal_10970, mcs1_mcs_mat1_4_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_17080, new_AGEMA_signal_17079, new_AGEMA_signal_17078, mcs1_mcs_mat1_4_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_15082, new_AGEMA_signal_15081, new_AGEMA_signal_15080, mcs1_mcs_mat1_4_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .c ({new_AGEMA_signal_16219, new_AGEMA_signal_16218, new_AGEMA_signal_16217, mcs1_mcs_mat1_4_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_9766, new_AGEMA_signal_9765, new_AGEMA_signal_9764, mcs1_mcs_mat1_4_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_13624, new_AGEMA_signal_13623, new_AGEMA_signal_13622, mcs1_mcs_mat1_4_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_15082, new_AGEMA_signal_15081, new_AGEMA_signal_15080, mcs1_mcs_mat1_4_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_8917, new_AGEMA_signal_8916, new_AGEMA_signal_8915, mcs1_mcs_mat1_4_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_12187, new_AGEMA_signal_12186, new_AGEMA_signal_12185, mcs1_mcs_mat1_4_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_13624, new_AGEMA_signal_13623, new_AGEMA_signal_13622, mcs1_mcs_mat1_4_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920]}), .c ({new_AGEMA_signal_12187, new_AGEMA_signal_12186, new_AGEMA_signal_12185, mcs1_mcs_mat1_4_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4931], Fresh[4930], Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926]}), .c ({new_AGEMA_signal_9766, new_AGEMA_signal_9765, new_AGEMA_signal_9764, mcs1_mcs_mat1_4_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4937], Fresh[4936], Fresh[4935], Fresh[4934], Fresh[4933], Fresh[4932]}), .c ({new_AGEMA_signal_10972, new_AGEMA_signal_10971, new_AGEMA_signal_10970, mcs1_mcs_mat1_4_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_18439, new_AGEMA_signal_18438, new_AGEMA_signal_18437, mcs1_mcs_mat1_4_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_17083, new_AGEMA_signal_17082, new_AGEMA_signal_17081, mcs1_mcs_mat1_4_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_19084, new_AGEMA_signal_19083, new_AGEMA_signal_19082, mcs1_mcs_mat1_4_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_15085, new_AGEMA_signal_15084, new_AGEMA_signal_15083, mcs1_mcs_mat1_4_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_17767, new_AGEMA_signal_17766, new_AGEMA_signal_17765, mcs1_mcs_mat1_4_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_18433, new_AGEMA_signal_18432, new_AGEMA_signal_18431, mcs1_mcs_mat1_4_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({new_AGEMA_signal_17770, new_AGEMA_signal_17769, new_AGEMA_signal_17768, mcs1_mcs_mat1_4_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_18436, new_AGEMA_signal_18435, new_AGEMA_signal_18434, mcs1_mcs_mat1_4_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940], Fresh[4939], Fresh[4938]}), .c ({new_AGEMA_signal_17770, new_AGEMA_signal_17769, new_AGEMA_signal_17768, mcs1_mcs_mat1_4_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944]}), .c ({new_AGEMA_signal_15085, new_AGEMA_signal_15084, new_AGEMA_signal_15083, mcs1_mcs_mat1_4_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950]}), .c ({new_AGEMA_signal_17083, new_AGEMA_signal_17082, new_AGEMA_signal_17081, mcs1_mcs_mat1_4_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_9772, new_AGEMA_signal_9771, new_AGEMA_signal_9770, mcs1_mcs_mat1_4_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_10975, new_AGEMA_signal_10974, new_AGEMA_signal_10973, mcs1_mcs_mat1_4_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_12190, new_AGEMA_signal_12189, new_AGEMA_signal_12188, mcs1_mcs_mat1_4_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_9775, new_AGEMA_signal_9774, new_AGEMA_signal_9773, mcs1_mcs_mat1_4_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_12193, new_AGEMA_signal_12192, new_AGEMA_signal_12191, mcs1_mcs_mat1_4_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_13633, new_AGEMA_signal_13632, new_AGEMA_signal_13631, mcs1_mcs_mat1_4_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_13636, new_AGEMA_signal_13635, new_AGEMA_signal_13634, mcs1_mcs_mat1_4_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_12196, new_AGEMA_signal_12195, new_AGEMA_signal_12194, mcs1_mcs_mat1_4_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_15088, new_AGEMA_signal_15087, new_AGEMA_signal_15086, mcs1_mcs_mat1_4_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_12199, new_AGEMA_signal_12198, new_AGEMA_signal_12197, mcs1_mcs_mat1_4_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_13636, new_AGEMA_signal_13635, new_AGEMA_signal_13634, mcs1_mcs_mat1_4_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4961], Fresh[4960], Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956]}), .c ({new_AGEMA_signal_12199, new_AGEMA_signal_12198, new_AGEMA_signal_12197, mcs1_mcs_mat1_4_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4967], Fresh[4966], Fresh[4965], Fresh[4964], Fresh[4963], Fresh[4962]}), .c ({new_AGEMA_signal_9775, new_AGEMA_signal_9774, new_AGEMA_signal_9773, mcs1_mcs_mat1_4_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970], Fresh[4969], Fresh[4968]}), .c ({new_AGEMA_signal_10975, new_AGEMA_signal_10974, new_AGEMA_signal_10973, mcs1_mcs_mat1_4_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_12205, new_AGEMA_signal_12204, new_AGEMA_signal_12203, mcs1_mcs_mat1_4_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_13639, new_AGEMA_signal_13638, new_AGEMA_signal_13637, mcs1_mcs_mat1_4_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_15091, new_AGEMA_signal_15090, new_AGEMA_signal_15089, mcs1_mcs_mat1_4_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_15094, new_AGEMA_signal_15093, new_AGEMA_signal_15092, mcs1_mcs_mat1_4_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_12202, new_AGEMA_signal_12201, new_AGEMA_signal_12200, mcs1_mcs_mat1_4_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_16222, new_AGEMA_signal_16221, new_AGEMA_signal_16220, mcs1_mcs_mat1_4_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_10978, new_AGEMA_signal_10977, new_AGEMA_signal_10976, mcs1_mcs_mat1_4_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_12202, new_AGEMA_signal_12201, new_AGEMA_signal_12200, mcs1_mcs_mat1_4_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({new_AGEMA_signal_15094, new_AGEMA_signal_15093, new_AGEMA_signal_15092, mcs1_mcs_mat1_4_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_16225, new_AGEMA_signal_16224, new_AGEMA_signal_16223, mcs1_mcs_mat1_4_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_8923, new_AGEMA_signal_8922, new_AGEMA_signal_8921, mcs1_mcs_mat1_4_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_13639, new_AGEMA_signal_13638, new_AGEMA_signal_13637, mcs1_mcs_mat1_4_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_15094, new_AGEMA_signal_15093, new_AGEMA_signal_15092, mcs1_mcs_mat1_4_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_9778, new_AGEMA_signal_9777, new_AGEMA_signal_9776, mcs1_mcs_mat1_4_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_12211, new_AGEMA_signal_12210, new_AGEMA_signal_12209, mcs1_mcs_mat1_4_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_13639, new_AGEMA_signal_13638, new_AGEMA_signal_13637, mcs1_mcs_mat1_4_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_12208, new_AGEMA_signal_12207, new_AGEMA_signal_12206, mcs1_mcs_mat1_4_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_13642, new_AGEMA_signal_13641, new_AGEMA_signal_13640, mcs1_mcs_mat1_4_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_15097, new_AGEMA_signal_15096, new_AGEMA_signal_15095, mcs1_mcs_mat1_4_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_12205, new_AGEMA_signal_12204, new_AGEMA_signal_12203, mcs1_mcs_mat1_4_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_9778, new_AGEMA_signal_9777, new_AGEMA_signal_9776, mcs1_mcs_mat1_4_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_13642, new_AGEMA_signal_13641, new_AGEMA_signal_13640, mcs1_mcs_mat1_4_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_10978, new_AGEMA_signal_10977, new_AGEMA_signal_10976, mcs1_mcs_mat1_4_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_12205, new_AGEMA_signal_12204, new_AGEMA_signal_12203, mcs1_mcs_mat1_4_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974]}), .c ({new_AGEMA_signal_12211, new_AGEMA_signal_12210, new_AGEMA_signal_12209, mcs1_mcs_mat1_4_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980]}), .c ({new_AGEMA_signal_9778, new_AGEMA_signal_9777, new_AGEMA_signal_9776, mcs1_mcs_mat1_4_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4991], Fresh[4990], Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986]}), .c ({new_AGEMA_signal_10978, new_AGEMA_signal_10977, new_AGEMA_signal_10976, mcs1_mcs_mat1_4_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_17089, new_AGEMA_signal_17088, new_AGEMA_signal_17087, mcs1_mcs_mat1_4_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_17773, new_AGEMA_signal_17772, new_AGEMA_signal_17771, mcs1_mcs_mat1_4_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_19810, new_AGEMA_signal_19809, new_AGEMA_signal_19808, mcs1_mcs_mat1_4_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_15100, new_AGEMA_signal_15099, new_AGEMA_signal_15098, mcs1_mcs_mat1_4_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_20620, new_AGEMA_signal_20619, new_AGEMA_signal_20618, mcs1_mcs_mat1_4_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_19090, new_AGEMA_signal_19089, new_AGEMA_signal_19088, mcs1_mcs_mat1_4_mcs_out[47]}), .b ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .c ({new_AGEMA_signal_19810, new_AGEMA_signal_19809, new_AGEMA_signal_19808, mcs1_mcs_mat1_4_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_18442, new_AGEMA_signal_18441, new_AGEMA_signal_18440, mcs1_mcs_mat1_4_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .c ({new_AGEMA_signal_19090, new_AGEMA_signal_19089, new_AGEMA_signal_19088, mcs1_mcs_mat1_4_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_13648, new_AGEMA_signal_13647, new_AGEMA_signal_13646, mcs1_mcs_mat1_4_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_17776, new_AGEMA_signal_17775, new_AGEMA_signal_17774, mcs1_mcs_mat1_4_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_18442, new_AGEMA_signal_18441, new_AGEMA_signal_18440, mcs1_mcs_mat1_4_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[4997], Fresh[4996], Fresh[4995], Fresh[4994], Fresh[4993], Fresh[4992]}), .c ({new_AGEMA_signal_17776, new_AGEMA_signal_17775, new_AGEMA_signal_17774, mcs1_mcs_mat1_4_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000], Fresh[4999], Fresh[4998]}), .c ({new_AGEMA_signal_15100, new_AGEMA_signal_15099, new_AGEMA_signal_15098, mcs1_mcs_mat1_4_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004]}), .c ({new_AGEMA_signal_17089, new_AGEMA_signal_17088, new_AGEMA_signal_17087, mcs1_mcs_mat1_4_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_13651, new_AGEMA_signal_13650, new_AGEMA_signal_13649, mcs1_mcs_mat1_4_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_10981, new_AGEMA_signal_10980, new_AGEMA_signal_10979, mcs1_mcs_mat1_4_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_15103, new_AGEMA_signal_15102, new_AGEMA_signal_15101, mcs1_mcs_mat1_4_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_12217, new_AGEMA_signal_12216, new_AGEMA_signal_12215, mcs1_mcs_mat1_4_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9781, new_AGEMA_signal_9780, new_AGEMA_signal_9779, mcs1_mcs_mat1_4_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_13651, new_AGEMA_signal_13650, new_AGEMA_signal_13649, mcs1_mcs_mat1_4_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_13654, new_AGEMA_signal_13653, new_AGEMA_signal_13652, mcs1_mcs_mat1_4_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_12223, new_AGEMA_signal_12222, new_AGEMA_signal_12221, mcs1_mcs_mat1_4_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_15106, new_AGEMA_signal_15105, new_AGEMA_signal_15104, mcs1_mcs_mat1_4_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_13657, new_AGEMA_signal_13656, new_AGEMA_signal_13655, mcs1_mcs_mat1_4_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_8926, new_AGEMA_signal_8925, new_AGEMA_signal_8924, mcs1_mcs_mat1_4_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_15109, new_AGEMA_signal_15108, new_AGEMA_signal_15107, mcs1_mcs_mat1_4_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_12217, new_AGEMA_signal_12216, new_AGEMA_signal_12215, mcs1_mcs_mat1_4_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_10984, new_AGEMA_signal_10983, new_AGEMA_signal_10982, mcs1_mcs_mat1_4_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_13657, new_AGEMA_signal_13656, new_AGEMA_signal_13655, mcs1_mcs_mat1_4_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_12220, new_AGEMA_signal_12219, new_AGEMA_signal_12218, mcs1_mcs_mat1_4_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_10984, new_AGEMA_signal_10983, new_AGEMA_signal_10982, mcs1_mcs_mat1_4_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_13660, new_AGEMA_signal_13659, new_AGEMA_signal_13658, mcs1_mcs_mat1_4_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010]}), .c ({new_AGEMA_signal_12223, new_AGEMA_signal_12222, new_AGEMA_signal_12221, mcs1_mcs_mat1_4_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5021], Fresh[5020], Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016]}), .c ({new_AGEMA_signal_9781, new_AGEMA_signal_9780, new_AGEMA_signal_9779, mcs1_mcs_mat1_4_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5027], Fresh[5026], Fresh[5025], Fresh[5024], Fresh[5023], Fresh[5022]}), .c ({new_AGEMA_signal_10984, new_AGEMA_signal_10983, new_AGEMA_signal_10982, mcs1_mcs_mat1_4_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_15112, new_AGEMA_signal_15111, new_AGEMA_signal_15110, mcs1_mcs_mat1_4_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_8929, new_AGEMA_signal_8928, new_AGEMA_signal_8927, mcs1_mcs_mat1_4_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_16228, new_AGEMA_signal_16227, new_AGEMA_signal_16226, mcs1_mcs_mat1_4_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_10990, new_AGEMA_signal_10989, new_AGEMA_signal_10988, mcs1_mcs_mat1_4_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_10987, new_AGEMA_signal_10986, new_AGEMA_signal_10985, mcs1_mcs_mat1_4_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_12226, new_AGEMA_signal_12225, new_AGEMA_signal_12224, mcs1_mcs_mat1_4_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({new_AGEMA_signal_15112, new_AGEMA_signal_15111, new_AGEMA_signal_15110, mcs1_mcs_mat1_4_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_16231, new_AGEMA_signal_16230, new_AGEMA_signal_16229, mcs1_mcs_mat1_4_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_12229, new_AGEMA_signal_12228, new_AGEMA_signal_12227, mcs1_mcs_mat1_4_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_13663, new_AGEMA_signal_13662, new_AGEMA_signal_13661, mcs1_mcs_mat1_4_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_15112, new_AGEMA_signal_15111, new_AGEMA_signal_15110, mcs1_mcs_mat1_4_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_12232, new_AGEMA_signal_12231, new_AGEMA_signal_12230, mcs1_mcs_mat1_4_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_10993, new_AGEMA_signal_10992, new_AGEMA_signal_10991, mcs1_mcs_mat1_4_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_13663, new_AGEMA_signal_13662, new_AGEMA_signal_13661, mcs1_mcs_mat1_4_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_12232, new_AGEMA_signal_12231, new_AGEMA_signal_12230, mcs1_mcs_mat1_4_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_10990, new_AGEMA_signal_10989, new_AGEMA_signal_10988, mcs1_mcs_mat1_4_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_13666, new_AGEMA_signal_13665, new_AGEMA_signal_13664, mcs1_mcs_mat1_4_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .b ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, new_AGEMA_signal_10322, mcs1_mcs_mat1_4_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_10990, new_AGEMA_signal_10989, new_AGEMA_signal_10988, mcs1_mcs_mat1_4_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({new_AGEMA_signal_9784, new_AGEMA_signal_9783, new_AGEMA_signal_9782, mcs1_mcs_mat1_4_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_10324, new_AGEMA_signal_10323, new_AGEMA_signal_10322, mcs1_mcs_mat1_4_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030], Fresh[5029], Fresh[5028]}), .c ({new_AGEMA_signal_12232, new_AGEMA_signal_12231, new_AGEMA_signal_12230, mcs1_mcs_mat1_4_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034]}), .c ({new_AGEMA_signal_9784, new_AGEMA_signal_9783, new_AGEMA_signal_9782, mcs1_mcs_mat1_4_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040]}), .c ({new_AGEMA_signal_10993, new_AGEMA_signal_10992, new_AGEMA_signal_10991, mcs1_mcs_mat1_4_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_12235, new_AGEMA_signal_12234, new_AGEMA_signal_12233, mcs1_mcs_mat1_4_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_10996, new_AGEMA_signal_10995, new_AGEMA_signal_10994, mcs1_mcs_mat1_4_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_13669, new_AGEMA_signal_13668, new_AGEMA_signal_13667, mcs1_mcs_mat1_4_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_9787, new_AGEMA_signal_9786, new_AGEMA_signal_9785, mcs1_mcs_mat1_4_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_10327, new_AGEMA_signal_10326, new_AGEMA_signal_10325, mcs1_mcs_mat1_4_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_16234, new_AGEMA_signal_16233, new_AGEMA_signal_16232, mcs1_mcs_mat1_4_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_12238, new_AGEMA_signal_12237, new_AGEMA_signal_12236, mcs1_mcs_mat1_4_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_17092, new_AGEMA_signal_17091, new_AGEMA_signal_17090, mcs1_mcs_mat1_4_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5051], Fresh[5050], Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046]}), .c ({new_AGEMA_signal_12238, new_AGEMA_signal_12237, new_AGEMA_signal_12236, mcs1_mcs_mat1_4_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5057], Fresh[5056], Fresh[5055], Fresh[5054], Fresh[5053], Fresh[5052]}), .c ({new_AGEMA_signal_9787, new_AGEMA_signal_9786, new_AGEMA_signal_9785, mcs1_mcs_mat1_4_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060], Fresh[5059], Fresh[5058]}), .c ({new_AGEMA_signal_10996, new_AGEMA_signal_10995, new_AGEMA_signal_10994, mcs1_mcs_mat1_4_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_19093, new_AGEMA_signal_19092, new_AGEMA_signal_19091, mcs1_mcs_mat1_4_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_18445, new_AGEMA_signal_18444, new_AGEMA_signal_18443, mcs1_mcs_mat1_4_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_19813, new_AGEMA_signal_19812, new_AGEMA_signal_19811, mcs1_mcs_mat1_4_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_15121, new_AGEMA_signal_15120, new_AGEMA_signal_15119, mcs1_mcs_mat1_4_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_18448, new_AGEMA_signal_18447, new_AGEMA_signal_18446, mcs1_mcs_mat1_4_mcs_out[29]}), .c ({new_AGEMA_signal_19093, new_AGEMA_signal_19092, new_AGEMA_signal_19091, mcs1_mcs_mat1_4_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_15118, new_AGEMA_signal_15117, new_AGEMA_signal_15116, mcs1_mcs_mat1_4_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_18445, new_AGEMA_signal_18444, new_AGEMA_signal_18443, mcs1_mcs_mat1_4_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_19096, new_AGEMA_signal_19095, new_AGEMA_signal_19094, mcs1_mcs_mat1_4_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_17785, new_AGEMA_signal_17784, new_AGEMA_signal_17783, mcs1_mcs_mat1_4_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .c ({new_AGEMA_signal_18445, new_AGEMA_signal_18444, new_AGEMA_signal_18443, mcs1_mcs_mat1_4_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_19099, new_AGEMA_signal_19098, new_AGEMA_signal_19097, mcs1_mcs_mat1_4_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_17779, new_AGEMA_signal_17778, new_AGEMA_signal_17777, mcs1_mcs_mat1_4_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_19816, new_AGEMA_signal_19815, new_AGEMA_signal_19814, mcs1_mcs_mat1_4_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_18451, new_AGEMA_signal_18450, new_AGEMA_signal_18449, mcs1_mcs_mat1_4_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_17782, new_AGEMA_signal_17781, new_AGEMA_signal_17780, mcs1_mcs_mat1_4_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_19099, new_AGEMA_signal_19098, new_AGEMA_signal_19097, mcs1_mcs_mat1_4_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_17095, new_AGEMA_signal_17094, new_AGEMA_signal_17093, mcs1_mcs_mat1_4_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_17782, new_AGEMA_signal_17781, new_AGEMA_signal_17780, mcs1_mcs_mat1_4_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_17785, new_AGEMA_signal_17784, new_AGEMA_signal_17783, mcs1_mcs_mat1_4_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_15121, new_AGEMA_signal_15120, new_AGEMA_signal_15119, mcs1_mcs_mat1_4_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_18451, new_AGEMA_signal_18450, new_AGEMA_signal_18449, mcs1_mcs_mat1_4_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064]}), .c ({new_AGEMA_signal_17785, new_AGEMA_signal_17784, new_AGEMA_signal_17783, mcs1_mcs_mat1_4_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070]}), .c ({new_AGEMA_signal_15121, new_AGEMA_signal_15120, new_AGEMA_signal_15119, mcs1_mcs_mat1_4_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5081], Fresh[5080], Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076]}), .c ({new_AGEMA_signal_17095, new_AGEMA_signal_17094, new_AGEMA_signal_17093, mcs1_mcs_mat1_4_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_12241, new_AGEMA_signal_12240, new_AGEMA_signal_12239, mcs1_mcs_mat1_4_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_13678, new_AGEMA_signal_13677, new_AGEMA_signal_13676, mcs1_mcs_mat1_4_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_10999, new_AGEMA_signal_10998, new_AGEMA_signal_10997, mcs1_mcs_mat1_4_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_9790, new_AGEMA_signal_9789, new_AGEMA_signal_9788, mcs1_mcs_mat1_4_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_12241, new_AGEMA_signal_12240, new_AGEMA_signal_12239, mcs1_mcs_mat1_4_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_13681, new_AGEMA_signal_13680, new_AGEMA_signal_13679, mcs1_mcs_mat1_4_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_15124, new_AGEMA_signal_15123, new_AGEMA_signal_15122, mcs1_mcs_mat1_4_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_12247, new_AGEMA_signal_12246, new_AGEMA_signal_12245, mcs1_mcs_mat1_4_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_9790, new_AGEMA_signal_9789, new_AGEMA_signal_9788, mcs1_mcs_mat1_4_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_13681, new_AGEMA_signal_13680, new_AGEMA_signal_13679, mcs1_mcs_mat1_4_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_15127, new_AGEMA_signal_15126, new_AGEMA_signal_15125, mcs1_mcs_mat1_4_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .c ({new_AGEMA_signal_16237, new_AGEMA_signal_16236, new_AGEMA_signal_16235, mcs1_mcs_mat1_4_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_12247, new_AGEMA_signal_12246, new_AGEMA_signal_12245, mcs1_mcs_mat1_4_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_13684, new_AGEMA_signal_13683, new_AGEMA_signal_13682, mcs1_mcs_mat1_4_mcs_out[24]}), .c ({new_AGEMA_signal_15127, new_AGEMA_signal_15126, new_AGEMA_signal_15125, mcs1_mcs_mat1_4_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_12244, new_AGEMA_signal_12243, new_AGEMA_signal_12242, mcs1_mcs_mat1_4_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .c ({new_AGEMA_signal_13684, new_AGEMA_signal_13683, new_AGEMA_signal_13682, mcs1_mcs_mat1_4_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_10999, new_AGEMA_signal_10998, new_AGEMA_signal_10997, mcs1_mcs_mat1_4_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_8935, new_AGEMA_signal_8934, new_AGEMA_signal_8933, mcs1_mcs_mat1_4_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_12244, new_AGEMA_signal_12243, new_AGEMA_signal_12242, mcs1_mcs_mat1_4_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5087], Fresh[5086], Fresh[5085], Fresh[5084], Fresh[5083], Fresh[5082]}), .c ({new_AGEMA_signal_12247, new_AGEMA_signal_12246, new_AGEMA_signal_12245, mcs1_mcs_mat1_4_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090], Fresh[5089], Fresh[5088]}), .c ({new_AGEMA_signal_9790, new_AGEMA_signal_9789, new_AGEMA_signal_9788, mcs1_mcs_mat1_4_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094]}), .c ({new_AGEMA_signal_10999, new_AGEMA_signal_10998, new_AGEMA_signal_10997, mcs1_mcs_mat1_4_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_12250, new_AGEMA_signal_12249, new_AGEMA_signal_12248, mcs1_mcs_mat1_4_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .c ({new_AGEMA_signal_13687, new_AGEMA_signal_13686, new_AGEMA_signal_13685, mcs1_mcs_mat1_4_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_11002, new_AGEMA_signal_11001, new_AGEMA_signal_11000, mcs1_mcs_mat1_4_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_9793, new_AGEMA_signal_9792, new_AGEMA_signal_9791, mcs1_mcs_mat1_4_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_12250, new_AGEMA_signal_12249, new_AGEMA_signal_12248, mcs1_mcs_mat1_4_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_13690, new_AGEMA_signal_13689, new_AGEMA_signal_13688, mcs1_mcs_mat1_4_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .c ({new_AGEMA_signal_15130, new_AGEMA_signal_15129, new_AGEMA_signal_15128, mcs1_mcs_mat1_4_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_12256, new_AGEMA_signal_12255, new_AGEMA_signal_12254, mcs1_mcs_mat1_4_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_9793, new_AGEMA_signal_9792, new_AGEMA_signal_9791, mcs1_mcs_mat1_4_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_13690, new_AGEMA_signal_13689, new_AGEMA_signal_13688, mcs1_mcs_mat1_4_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_15133, new_AGEMA_signal_15132, new_AGEMA_signal_15131, mcs1_mcs_mat1_4_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_8404, new_AGEMA_signal_8403, new_AGEMA_signal_8402, mcs1_mcs_mat1_4_mcs_out[86]}), .c ({new_AGEMA_signal_16240, new_AGEMA_signal_16239, new_AGEMA_signal_16238, mcs1_mcs_mat1_4_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_12256, new_AGEMA_signal_12255, new_AGEMA_signal_12254, mcs1_mcs_mat1_4_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_13693, new_AGEMA_signal_13692, new_AGEMA_signal_13691, mcs1_mcs_mat1_4_mcs_out[20]}), .c ({new_AGEMA_signal_15133, new_AGEMA_signal_15132, new_AGEMA_signal_15131, mcs1_mcs_mat1_4_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_12253, new_AGEMA_signal_12252, new_AGEMA_signal_12251, mcs1_mcs_mat1_4_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .c ({new_AGEMA_signal_13693, new_AGEMA_signal_13692, new_AGEMA_signal_13691, mcs1_mcs_mat1_4_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_11002, new_AGEMA_signal_11001, new_AGEMA_signal_11000, mcs1_mcs_mat1_4_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_8938, new_AGEMA_signal_8937, new_AGEMA_signal_8936, mcs1_mcs_mat1_4_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_12253, new_AGEMA_signal_12252, new_AGEMA_signal_12251, mcs1_mcs_mat1_4_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100]}), .c ({new_AGEMA_signal_12256, new_AGEMA_signal_12255, new_AGEMA_signal_12254, mcs1_mcs_mat1_4_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5111], Fresh[5110], Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106]}), .c ({new_AGEMA_signal_9793, new_AGEMA_signal_9792, new_AGEMA_signal_9791, mcs1_mcs_mat1_4_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5117], Fresh[5116], Fresh[5115], Fresh[5114], Fresh[5113], Fresh[5112]}), .c ({new_AGEMA_signal_11002, new_AGEMA_signal_11001, new_AGEMA_signal_11000, mcs1_mcs_mat1_4_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_12259, new_AGEMA_signal_12258, new_AGEMA_signal_12257, mcs1_mcs_mat1_4_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_12268, new_AGEMA_signal_12267, new_AGEMA_signal_12266, mcs1_mcs_mat1_4_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_13696, new_AGEMA_signal_13695, new_AGEMA_signal_13694, mcs1_mcs_mat1_4_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_13699, new_AGEMA_signal_13698, new_AGEMA_signal_13697, mcs1_mcs_mat1_4_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_8941, new_AGEMA_signal_8940, new_AGEMA_signal_8939, mcs1_mcs_mat1_4_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_15136, new_AGEMA_signal_15135, new_AGEMA_signal_15134, mcs1_mcs_mat1_4_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_15139, new_AGEMA_signal_15138, new_AGEMA_signal_15137, mcs1_mcs_mat1_4_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_9796, new_AGEMA_signal_9795, new_AGEMA_signal_9794, mcs1_mcs_mat1_4_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_16243, new_AGEMA_signal_16242, new_AGEMA_signal_16241, mcs1_mcs_mat1_4_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_8422, new_AGEMA_signal_8421, new_AGEMA_signal_8420, mcs1_mcs_mat1_4_mcs_out[50]}), .b ({new_AGEMA_signal_13699, new_AGEMA_signal_13698, new_AGEMA_signal_13697, mcs1_mcs_mat1_4_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_15139, new_AGEMA_signal_15138, new_AGEMA_signal_15137, mcs1_mcs_mat1_4_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_12262, new_AGEMA_signal_12261, new_AGEMA_signal_12260, mcs1_mcs_mat1_4_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .c ({new_AGEMA_signal_13699, new_AGEMA_signal_13698, new_AGEMA_signal_13697, mcs1_mcs_mat1_4_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_11005, new_AGEMA_signal_11004, new_AGEMA_signal_11003, mcs1_mcs_mat1_4_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_11008, new_AGEMA_signal_11007, new_AGEMA_signal_11006, mcs1_mcs_mat1_4_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_12262, new_AGEMA_signal_12261, new_AGEMA_signal_12260, mcs1_mcs_mat1_4_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_12265, new_AGEMA_signal_12264, new_AGEMA_signal_12263, mcs1_mcs_mat1_4_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_9796, new_AGEMA_signal_9795, new_AGEMA_signal_9794, mcs1_mcs_mat1_4_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_13702, new_AGEMA_signal_13701, new_AGEMA_signal_13700, mcs1_mcs_mat1_4_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120], Fresh[5119], Fresh[5118]}), .c ({new_AGEMA_signal_12268, new_AGEMA_signal_12267, new_AGEMA_signal_12266, mcs1_mcs_mat1_4_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124]}), .c ({new_AGEMA_signal_9796, new_AGEMA_signal_9795, new_AGEMA_signal_9794, mcs1_mcs_mat1_4_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130]}), .c ({new_AGEMA_signal_11008, new_AGEMA_signal_11007, new_AGEMA_signal_11006, mcs1_mcs_mat1_4_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_19108, new_AGEMA_signal_19107, new_AGEMA_signal_19106, mcs1_mcs_mat1_4_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_16246, new_AGEMA_signal_16245, new_AGEMA_signal_16244, mcs1_mcs_mat1_4_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_19819, new_AGEMA_signal_19818, new_AGEMA_signal_19817, mcs1_mcs_mat1_4_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_18460, new_AGEMA_signal_18459, new_AGEMA_signal_18458, mcs1_mcs_mat1_4_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_18454, new_AGEMA_signal_18453, new_AGEMA_signal_18452, mcs1_mcs_mat1_4_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_19102, new_AGEMA_signal_19101, new_AGEMA_signal_19100, mcs1_mcs_mat1_4_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_17791, new_AGEMA_signal_17790, new_AGEMA_signal_17789, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_15142, new_AGEMA_signal_15141, new_AGEMA_signal_15140, mcs1_mcs_mat1_4_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_18454, new_AGEMA_signal_18453, new_AGEMA_signal_18452, mcs1_mcs_mat1_4_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_16246, new_AGEMA_signal_16245, new_AGEMA_signal_16244, mcs1_mcs_mat1_4_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_18457, new_AGEMA_signal_18456, new_AGEMA_signal_18455, mcs1_mcs_mat1_4_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_19105, new_AGEMA_signal_19104, new_AGEMA_signal_19103, mcs1_mcs_mat1_4_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_17788, new_AGEMA_signal_17787, new_AGEMA_signal_17786, mcs1_mcs_mat1_4_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_17791, new_AGEMA_signal_17790, new_AGEMA_signal_17789, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_18457, new_AGEMA_signal_18456, new_AGEMA_signal_18455, mcs1_mcs_mat1_4_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_13705, new_AGEMA_signal_13704, new_AGEMA_signal_13703, mcs1_mcs_mat1_4_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_15142, new_AGEMA_signal_15141, new_AGEMA_signal_15140, mcs1_mcs_mat1_4_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_16246, new_AGEMA_signal_16245, new_AGEMA_signal_16244, mcs1_mcs_mat1_4_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_19822, new_AGEMA_signal_19821, new_AGEMA_signal_19820, mcs1_mcs_mat1_4_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .c ({new_AGEMA_signal_20623, new_AGEMA_signal_20622, new_AGEMA_signal_20621, mcs1_mcs_mat1_4_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_19108, new_AGEMA_signal_19107, new_AGEMA_signal_19106, mcs1_mcs_mat1_4_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_17791, new_AGEMA_signal_17790, new_AGEMA_signal_17789, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_19822, new_AGEMA_signal_19821, new_AGEMA_signal_19820, mcs1_mcs_mat1_4_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({new_AGEMA_signal_18460, new_AGEMA_signal_18459, new_AGEMA_signal_18458, mcs1_mcs_mat1_4_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_19108, new_AGEMA_signal_19107, new_AGEMA_signal_19106, mcs1_mcs_mat1_4_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({new_AGEMA_signal_17788, new_AGEMA_signal_17787, new_AGEMA_signal_17786, mcs1_mcs_mat1_4_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_18460, new_AGEMA_signal_18459, new_AGEMA_signal_18458, mcs1_mcs_mat1_4_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_11380, new_AGEMA_signal_11379, new_AGEMA_signal_11378, shiftr_out[108]}), .b ({new_AGEMA_signal_17098, new_AGEMA_signal_17097, new_AGEMA_signal_17096, mcs1_mcs_mat1_4_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_17788, new_AGEMA_signal_17787, new_AGEMA_signal_17786, mcs1_mcs_mat1_4_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16606, new_AGEMA_signal_16605, new_AGEMA_signal_16604, mcs1_mcs_mat1_4_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5141], Fresh[5140], Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136]}), .c ({new_AGEMA_signal_17791, new_AGEMA_signal_17790, new_AGEMA_signal_17789, mcs1_mcs_mat1_4_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12820, new_AGEMA_signal_12819, new_AGEMA_signal_12818, mcs1_mcs_mat1_4_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5147], Fresh[5146], Fresh[5145], Fresh[5144], Fresh[5143], Fresh[5142]}), .c ({new_AGEMA_signal_15142, new_AGEMA_signal_15141, new_AGEMA_signal_15140, mcs1_mcs_mat1_4_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15694, new_AGEMA_signal_15693, new_AGEMA_signal_15692, mcs1_mcs_mat1_4_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150], Fresh[5149], Fresh[5148]}), .c ({new_AGEMA_signal_17098, new_AGEMA_signal_17097, new_AGEMA_signal_17096, mcs1_mcs_mat1_4_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, new_AGEMA_signal_10328, mcs1_mcs_mat1_4_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .c ({new_AGEMA_signal_11011, new_AGEMA_signal_11010, new_AGEMA_signal_11009, mcs1_mcs_mat1_4_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_13711, new_AGEMA_signal_13710, new_AGEMA_signal_13709, mcs1_mcs_mat1_4_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .c ({new_AGEMA_signal_15145, new_AGEMA_signal_15144, new_AGEMA_signal_15143, mcs1_mcs_mat1_4_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_12271, new_AGEMA_signal_12270, new_AGEMA_signal_12269, mcs1_mcs_mat1_4_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .c ({new_AGEMA_signal_13708, new_AGEMA_signal_13707, new_AGEMA_signal_13706, mcs1_mcs_mat1_4_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_11014, new_AGEMA_signal_11013, new_AGEMA_signal_11012, mcs1_mcs_mat1_4_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, new_AGEMA_signal_10328, mcs1_mcs_mat1_4_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_12271, new_AGEMA_signal_12270, new_AGEMA_signal_12269, mcs1_mcs_mat1_4_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_8944, new_AGEMA_signal_8943, new_AGEMA_signal_8942, mcs1_mcs_mat1_4_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_9799, new_AGEMA_signal_9798, new_AGEMA_signal_9797, mcs1_mcs_mat1_4_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_10330, new_AGEMA_signal_10329, new_AGEMA_signal_10328, mcs1_mcs_mat1_4_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_15148, new_AGEMA_signal_15147, new_AGEMA_signal_15146, mcs1_mcs_mat1_4_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_8386, new_AGEMA_signal_8385, new_AGEMA_signal_8384, shiftr_out[76]}), .c ({new_AGEMA_signal_16249, new_AGEMA_signal_16248, new_AGEMA_signal_16247, mcs1_mcs_mat1_4_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_8944, new_AGEMA_signal_8943, new_AGEMA_signal_8942, mcs1_mcs_mat1_4_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_13711, new_AGEMA_signal_13710, new_AGEMA_signal_13709, mcs1_mcs_mat1_4_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_15148, new_AGEMA_signal_15147, new_AGEMA_signal_15146, mcs1_mcs_mat1_4_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_12274, new_AGEMA_signal_12273, new_AGEMA_signal_12272, mcs1_mcs_mat1_4_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_11014, new_AGEMA_signal_11013, new_AGEMA_signal_11012, mcs1_mcs_mat1_4_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_13711, new_AGEMA_signal_13710, new_AGEMA_signal_13709, mcs1_mcs_mat1_4_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10425, new_AGEMA_signal_10424, mcs1_mcs_mat1_4_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154]}), .c ({new_AGEMA_signal_12274, new_AGEMA_signal_12273, new_AGEMA_signal_12272, mcs1_mcs_mat1_4_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8590, new_AGEMA_signal_8589, new_AGEMA_signal_8588, mcs1_mcs_mat1_4_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160]}), .c ({new_AGEMA_signal_9799, new_AGEMA_signal_9798, new_AGEMA_signal_9797, mcs1_mcs_mat1_4_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10228, new_AGEMA_signal_10227, new_AGEMA_signal_10226, shiftr_out[79]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5171], Fresh[5170], Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166]}), .c ({new_AGEMA_signal_11014, new_AGEMA_signal_11013, new_AGEMA_signal_11012, mcs1_mcs_mat1_4_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_17101, new_AGEMA_signal_17100, new_AGEMA_signal_17099, mcs1_mcs_mat1_4_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_11020, new_AGEMA_signal_11019, new_AGEMA_signal_11018, mcs1_mcs_mat1_4_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_17794, new_AGEMA_signal_17793, new_AGEMA_signal_17792, mcs1_mcs_mat1_4_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_16252, new_AGEMA_signal_16251, new_AGEMA_signal_16250, mcs1_mcs_mat1_4_mcs_out[7]}), .b ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .c ({new_AGEMA_signal_17101, new_AGEMA_signal_17100, new_AGEMA_signal_17099, mcs1_mcs_mat1_4_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_15151, new_AGEMA_signal_15150, new_AGEMA_signal_15149, mcs1_mcs_mat1_4_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .c ({new_AGEMA_signal_16252, new_AGEMA_signal_16251, new_AGEMA_signal_16250, mcs1_mcs_mat1_4_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_13714, new_AGEMA_signal_13713, new_AGEMA_signal_13712, mcs1_mcs_mat1_4_mcs_out[6]}), .b ({new_AGEMA_signal_9805, new_AGEMA_signal_9804, new_AGEMA_signal_9803, mcs1_mcs_mat1_4_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_15151, new_AGEMA_signal_15150, new_AGEMA_signal_15149, mcs1_mcs_mat1_4_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_9802, new_AGEMA_signal_9801, new_AGEMA_signal_9800, mcs1_mcs_mat1_4_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_12277, new_AGEMA_signal_12276, new_AGEMA_signal_12275, mcs1_mcs_mat1_4_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_13714, new_AGEMA_signal_13713, new_AGEMA_signal_13712, mcs1_mcs_mat1_4_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10444, new_AGEMA_signal_10443, new_AGEMA_signal_10442, shiftr_out[45]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5177], Fresh[5176], Fresh[5175], Fresh[5174], Fresh[5173], Fresh[5172]}), .c ({new_AGEMA_signal_12277, new_AGEMA_signal_12276, new_AGEMA_signal_12275, mcs1_mcs_mat1_4_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8608, new_AGEMA_signal_8607, new_AGEMA_signal_8606, shiftr_out[46]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180], Fresh[5179], Fresh[5178]}), .c ({new_AGEMA_signal_9805, new_AGEMA_signal_9804, new_AGEMA_signal_9803, mcs1_mcs_mat1_4_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10246, new_AGEMA_signal_10245, new_AGEMA_signal_10244, mcs1_mcs_mat1_4_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184]}), .c ({new_AGEMA_signal_11020, new_AGEMA_signal_11019, new_AGEMA_signal_11018, mcs1_mcs_mat1_4_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_11023, new_AGEMA_signal_11022, new_AGEMA_signal_11021, mcs1_mcs_mat1_4_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_12280, new_AGEMA_signal_12279, new_AGEMA_signal_12278, mcs1_mcs_mat1_4_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_13720, new_AGEMA_signal_13719, new_AGEMA_signal_13718, mcs1_mcs_mat1_4_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .b ({new_AGEMA_signal_11026, new_AGEMA_signal_11025, new_AGEMA_signal_11024, mcs1_mcs_mat1_4_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_12280, new_AGEMA_signal_12279, new_AGEMA_signal_12278, mcs1_mcs_mat1_4_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_13723, new_AGEMA_signal_13722, new_AGEMA_signal_13721, mcs1_mcs_mat1_4_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_9808, new_AGEMA_signal_9807, new_AGEMA_signal_9806, mcs1_mcs_mat1_4_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_15154, new_AGEMA_signal_15153, new_AGEMA_signal_15152, mcs1_mcs_mat1_4_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_13726, new_AGEMA_signal_13725, new_AGEMA_signal_13724, mcs1_mcs_mat1_4_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_12286, new_AGEMA_signal_12285, new_AGEMA_signal_12284, mcs1_mcs_mat1_4_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_15157, new_AGEMA_signal_15156, new_AGEMA_signal_15155, mcs1_mcs_mat1_4_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_12289, new_AGEMA_signal_12288, new_AGEMA_signal_12287, mcs1_mcs_mat1_4_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_8950, new_AGEMA_signal_8949, new_AGEMA_signal_8948, mcs1_mcs_mat1_4_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_13726, new_AGEMA_signal_13725, new_AGEMA_signal_13724, mcs1_mcs_mat1_4_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10462, new_AGEMA_signal_10461, new_AGEMA_signal_10460, shiftr_out[13]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190]}), .c ({new_AGEMA_signal_12289, new_AGEMA_signal_12288, new_AGEMA_signal_12287, mcs1_mcs_mat1_4_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8626, new_AGEMA_signal_8625, new_AGEMA_signal_8624, shiftr_out[14]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5201], Fresh[5200], Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196]}), .c ({new_AGEMA_signal_9808, new_AGEMA_signal_9807, new_AGEMA_signal_9806, mcs1_mcs_mat1_4_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_4_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10264, new_AGEMA_signal_10263, new_AGEMA_signal_10262, mcs1_mcs_mat1_4_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5207], Fresh[5206], Fresh[5205], Fresh[5204], Fresh[5203], Fresh[5202]}), .c ({new_AGEMA_signal_11026, new_AGEMA_signal_11025, new_AGEMA_signal_11024, mcs1_mcs_mat1_4_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U96 ( .a ({new_AGEMA_signal_17104, new_AGEMA_signal_17103, new_AGEMA_signal_17102, mcs1_mcs_mat1_5_n128}), .b ({new_AGEMA_signal_16255, new_AGEMA_signal_16254, new_AGEMA_signal_16253, mcs1_mcs_mat1_5_n127}), .c ({temp_next_s3[73], temp_next_s2[73], temp_next_s1[73], temp_next_s0[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U95 ( .a ({new_AGEMA_signal_15286, new_AGEMA_signal_15285, new_AGEMA_signal_15284, mcs1_mcs_mat1_5_mcs_out[41]}), .b ({new_AGEMA_signal_12397, new_AGEMA_signal_12396, new_AGEMA_signal_12395, mcs1_mcs_mat1_5_mcs_out[45]}), .c ({new_AGEMA_signal_16255, new_AGEMA_signal_16254, new_AGEMA_signal_16253, mcs1_mcs_mat1_5_n127}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U94 ( .a ({new_AGEMA_signal_16354, new_AGEMA_signal_16353, new_AGEMA_signal_16352, mcs1_mcs_mat1_5_mcs_out[33]}), .b ({new_AGEMA_signal_16351, new_AGEMA_signal_16350, new_AGEMA_signal_16349, mcs1_mcs_mat1_5_mcs_out[37]}), .c ({new_AGEMA_signal_17104, new_AGEMA_signal_17103, new_AGEMA_signal_17102, mcs1_mcs_mat1_5_n128}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U93 ( .a ({new_AGEMA_signal_21277, new_AGEMA_signal_21276, new_AGEMA_signal_21275, mcs1_mcs_mat1_5_n126}), .b ({new_AGEMA_signal_17800, new_AGEMA_signal_17799, new_AGEMA_signal_17798, mcs1_mcs_mat1_5_n125}), .c ({temp_next_s3[72], temp_next_s2[72], temp_next_s1[72], temp_next_s0[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U92 ( .a ({new_AGEMA_signal_13840, new_AGEMA_signal_13839, new_AGEMA_signal_13838, mcs1_mcs_mat1_5_mcs_out[40]}), .b ({new_AGEMA_signal_17164, new_AGEMA_signal_17163, new_AGEMA_signal_17162, mcs1_mcs_mat1_5_mcs_out[44]}), .c ({new_AGEMA_signal_17800, new_AGEMA_signal_17799, new_AGEMA_signal_17798, mcs1_mcs_mat1_5_n125}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U91 ( .a ({new_AGEMA_signal_20665, new_AGEMA_signal_20664, new_AGEMA_signal_20663, mcs1_mcs_mat1_5_mcs_out[32]}), .b ({new_AGEMA_signal_13846, new_AGEMA_signal_13845, new_AGEMA_signal_13844, mcs1_mcs_mat1_5_mcs_out[36]}), .c ({new_AGEMA_signal_21277, new_AGEMA_signal_21276, new_AGEMA_signal_21275, mcs1_mcs_mat1_5_n126}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U90 ( .a ({new_AGEMA_signal_19111, new_AGEMA_signal_19110, new_AGEMA_signal_19109, mcs1_mcs_mat1_5_n124}), .b ({new_AGEMA_signal_17107, new_AGEMA_signal_17106, new_AGEMA_signal_17105, mcs1_mcs_mat1_5_n123}), .c ({temp_next_s3[43], temp_next_s2[43], temp_next_s1[43], temp_next_s0[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U89 ( .a ({new_AGEMA_signal_13861, new_AGEMA_signal_13860, new_AGEMA_signal_13859, mcs1_mcs_mat1_5_mcs_out[27]}), .b ({new_AGEMA_signal_16357, new_AGEMA_signal_16356, new_AGEMA_signal_16355, mcs1_mcs_mat1_5_mcs_out[31]}), .c ({new_AGEMA_signal_17107, new_AGEMA_signal_17106, new_AGEMA_signal_17105, mcs1_mcs_mat1_5_n123}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U88 ( .a ({new_AGEMA_signal_18514, new_AGEMA_signal_18513, new_AGEMA_signal_18512, mcs1_mcs_mat1_5_mcs_out[19]}), .b ({new_AGEMA_signal_13870, new_AGEMA_signal_13869, new_AGEMA_signal_13868, mcs1_mcs_mat1_5_mcs_out[23]}), .c ({new_AGEMA_signal_19111, new_AGEMA_signal_19110, new_AGEMA_signal_19109, mcs1_mcs_mat1_5_n124}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U87 ( .a ({new_AGEMA_signal_19828, new_AGEMA_signal_19827, new_AGEMA_signal_19826, mcs1_mcs_mat1_5_n122}), .b ({new_AGEMA_signal_16258, new_AGEMA_signal_16257, new_AGEMA_signal_16256, mcs1_mcs_mat1_5_n121}), .c ({temp_next_s3[42], temp_next_s2[42], temp_next_s1[42], temp_next_s0[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U86 ( .a ({new_AGEMA_signal_15304, new_AGEMA_signal_15303, new_AGEMA_signal_15302, mcs1_mcs_mat1_5_mcs_out[26]}), .b ({new_AGEMA_signal_15298, new_AGEMA_signal_15297, new_AGEMA_signal_15296, mcs1_mcs_mat1_5_mcs_out[30]}), .c ({new_AGEMA_signal_16258, new_AGEMA_signal_16257, new_AGEMA_signal_16256, mcs1_mcs_mat1_5_n121}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U85 ( .a ({new_AGEMA_signal_19174, new_AGEMA_signal_19173, new_AGEMA_signal_19172, mcs1_mcs_mat1_5_mcs_out[18]}), .b ({new_AGEMA_signal_15310, new_AGEMA_signal_15309, new_AGEMA_signal_15308, mcs1_mcs_mat1_5_mcs_out[22]}), .c ({new_AGEMA_signal_19828, new_AGEMA_signal_19827, new_AGEMA_signal_19826, mcs1_mcs_mat1_5_n122}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U84 ( .a ({new_AGEMA_signal_20629, new_AGEMA_signal_20628, new_AGEMA_signal_20627, mcs1_mcs_mat1_5_n120}), .b ({new_AGEMA_signal_17110, new_AGEMA_signal_17109, new_AGEMA_signal_17108, mcs1_mcs_mat1_5_n119}), .c ({temp_next_s3[41], temp_next_s2[41], temp_next_s1[41], temp_next_s0[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U83 ( .a ({new_AGEMA_signal_16363, new_AGEMA_signal_16362, new_AGEMA_signal_16361, mcs1_mcs_mat1_5_mcs_out[25]}), .b ({new_AGEMA_signal_13855, new_AGEMA_signal_13854, new_AGEMA_signal_13853, mcs1_mcs_mat1_5_mcs_out[29]}), .c ({new_AGEMA_signal_17110, new_AGEMA_signal_17109, new_AGEMA_signal_17108, mcs1_mcs_mat1_5_n119}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U82 ( .a ({new_AGEMA_signal_19894, new_AGEMA_signal_19893, new_AGEMA_signal_19892, mcs1_mcs_mat1_5_mcs_out[17]}), .b ({new_AGEMA_signal_16366, new_AGEMA_signal_16365, new_AGEMA_signal_16364, mcs1_mcs_mat1_5_mcs_out[21]}), .c ({new_AGEMA_signal_20629, new_AGEMA_signal_20628, new_AGEMA_signal_20627, mcs1_mcs_mat1_5_n120}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U81 ( .a ({new_AGEMA_signal_19114, new_AGEMA_signal_19113, new_AGEMA_signal_19112, mcs1_mcs_mat1_5_n118}), .b ({new_AGEMA_signal_17113, new_AGEMA_signal_17112, new_AGEMA_signal_17111, mcs1_mcs_mat1_5_n117}), .c ({temp_next_s3[40], temp_next_s2[40], temp_next_s1[40], temp_next_s0[40]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U80 ( .a ({new_AGEMA_signal_13867, new_AGEMA_signal_13866, new_AGEMA_signal_13865, mcs1_mcs_mat1_5_mcs_out[24]}), .b ({new_AGEMA_signal_16360, new_AGEMA_signal_16359, new_AGEMA_signal_16358, mcs1_mcs_mat1_5_mcs_out[28]}), .c ({new_AGEMA_signal_17113, new_AGEMA_signal_17112, new_AGEMA_signal_17111, mcs1_mcs_mat1_5_n117}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U79 ( .a ({new_AGEMA_signal_18520, new_AGEMA_signal_18519, new_AGEMA_signal_18518, mcs1_mcs_mat1_5_mcs_out[16]}), .b ({new_AGEMA_signal_13876, new_AGEMA_signal_13875, new_AGEMA_signal_13874, mcs1_mcs_mat1_5_mcs_out[20]}), .c ({new_AGEMA_signal_19114, new_AGEMA_signal_19113, new_AGEMA_signal_19112, mcs1_mcs_mat1_5_n118}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U78 ( .a ({new_AGEMA_signal_17116, new_AGEMA_signal_17115, new_AGEMA_signal_17114, mcs1_mcs_mat1_5_n116}), .b ({new_AGEMA_signal_19117, new_AGEMA_signal_19116, new_AGEMA_signal_19115, mcs1_mcs_mat1_5_n115}), .c ({temp_next_s3[11], temp_next_s2[11], temp_next_s1[11], temp_next_s0[11]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U77 ( .a ({new_AGEMA_signal_18523, new_AGEMA_signal_18522, new_AGEMA_signal_18521, mcs1_mcs_mat1_5_mcs_out[3]}), .b ({new_AGEMA_signal_16378, new_AGEMA_signal_16377, new_AGEMA_signal_16376, mcs1_mcs_mat1_5_mcs_out[7]}), .c ({new_AGEMA_signal_19117, new_AGEMA_signal_19116, new_AGEMA_signal_19115, mcs1_mcs_mat1_5_n115}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U76 ( .a ({new_AGEMA_signal_11131, new_AGEMA_signal_11130, new_AGEMA_signal_11129, mcs1_mcs_mat1_5_mcs_out[11]}), .b ({new_AGEMA_signal_16369, new_AGEMA_signal_16368, new_AGEMA_signal_16367, mcs1_mcs_mat1_5_mcs_out[15]}), .c ({new_AGEMA_signal_17116, new_AGEMA_signal_17115, new_AGEMA_signal_17114, mcs1_mcs_mat1_5_n116}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U75 ( .a ({new_AGEMA_signal_19837, new_AGEMA_signal_19836, new_AGEMA_signal_19835, mcs1_mcs_mat1_5_n114}), .b ({new_AGEMA_signal_17119, new_AGEMA_signal_17118, new_AGEMA_signal_17117, mcs1_mcs_mat1_5_n113}), .c ({new_AGEMA_signal_20632, new_AGEMA_signal_20631, new_AGEMA_signal_20630, mcs_out[235]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U74 ( .a ({new_AGEMA_signal_16291, new_AGEMA_signal_16290, new_AGEMA_signal_16289, mcs1_mcs_mat1_5_mcs_out[123]}), .b ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_17119, new_AGEMA_signal_17118, new_AGEMA_signal_17117, mcs1_mcs_mat1_5_n113}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U73 ( .a ({new_AGEMA_signal_19153, new_AGEMA_signal_19152, new_AGEMA_signal_19151, mcs1_mcs_mat1_5_mcs_out[115]}), .b ({new_AGEMA_signal_16297, new_AGEMA_signal_16296, new_AGEMA_signal_16295, mcs1_mcs_mat1_5_mcs_out[119]}), .c ({new_AGEMA_signal_19837, new_AGEMA_signal_19836, new_AGEMA_signal_19835, mcs1_mcs_mat1_5_n114}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U72 ( .a ({new_AGEMA_signal_19120, new_AGEMA_signal_19119, new_AGEMA_signal_19118, mcs1_mcs_mat1_5_n112}), .b ({new_AGEMA_signal_13729, new_AGEMA_signal_13728, new_AGEMA_signal_13727, mcs1_mcs_mat1_5_n111}), .c ({new_AGEMA_signal_19840, new_AGEMA_signal_19839, new_AGEMA_signal_19838, mcs_out[234]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U71 ( .a ({new_AGEMA_signal_12292, new_AGEMA_signal_12291, new_AGEMA_signal_12290, mcs1_mcs_mat1_5_mcs_out[122]}), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_13729, new_AGEMA_signal_13728, new_AGEMA_signal_13727, mcs1_mcs_mat1_5_n111}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U70 ( .a ({new_AGEMA_signal_18478, new_AGEMA_signal_18477, new_AGEMA_signal_18476, mcs1_mcs_mat1_5_mcs_out[114]}), .b ({new_AGEMA_signal_16300, new_AGEMA_signal_16299, new_AGEMA_signal_16298, mcs1_mcs_mat1_5_mcs_out[118]}), .c ({new_AGEMA_signal_19120, new_AGEMA_signal_19119, new_AGEMA_signal_19118, mcs1_mcs_mat1_5_n112}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U69 ( .a ({new_AGEMA_signal_16261, new_AGEMA_signal_16260, new_AGEMA_signal_16259, mcs1_mcs_mat1_5_n110}), .b ({new_AGEMA_signal_19123, new_AGEMA_signal_19122, new_AGEMA_signal_19121, mcs1_mcs_mat1_5_n109}), .c ({temp_next_s3[10], temp_next_s2[10], temp_next_s1[10], temp_next_s0[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U68 ( .a ({new_AGEMA_signal_18526, new_AGEMA_signal_18525, new_AGEMA_signal_18524, mcs1_mcs_mat1_5_mcs_out[2]}), .b ({new_AGEMA_signal_13897, new_AGEMA_signal_13896, new_AGEMA_signal_13895, mcs1_mcs_mat1_5_mcs_out[6]}), .c ({new_AGEMA_signal_19123, new_AGEMA_signal_19122, new_AGEMA_signal_19121, mcs1_mcs_mat1_5_n109}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U67 ( .a ({new_AGEMA_signal_15328, new_AGEMA_signal_15327, new_AGEMA_signal_15326, mcs1_mcs_mat1_5_mcs_out[10]}), .b ({new_AGEMA_signal_15319, new_AGEMA_signal_15318, new_AGEMA_signal_15317, mcs1_mcs_mat1_5_mcs_out[14]}), .c ({new_AGEMA_signal_16261, new_AGEMA_signal_16260, new_AGEMA_signal_16259, mcs1_mcs_mat1_5_n110}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U66 ( .a ({new_AGEMA_signal_18463, new_AGEMA_signal_18462, new_AGEMA_signal_18461, mcs1_mcs_mat1_5_n108}), .b ({new_AGEMA_signal_17122, new_AGEMA_signal_17121, new_AGEMA_signal_17120, mcs1_mcs_mat1_5_n107}), .c ({new_AGEMA_signal_19126, new_AGEMA_signal_19125, new_AGEMA_signal_19124, mcs_out[233]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U65 ( .a ({new_AGEMA_signal_16294, new_AGEMA_signal_16293, new_AGEMA_signal_16292, mcs1_mcs_mat1_5_mcs_out[121]}), .b ({new_AGEMA_signal_11029, new_AGEMA_signal_11028, new_AGEMA_signal_11027, mcs1_mcs_mat1_5_mcs_out[125]}), .c ({new_AGEMA_signal_17122, new_AGEMA_signal_17121, new_AGEMA_signal_17120, mcs1_mcs_mat1_5_n107}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U64 ( .a ({new_AGEMA_signal_17812, new_AGEMA_signal_17811, new_AGEMA_signal_17810, mcs1_mcs_mat1_5_mcs_out[113]}), .b ({new_AGEMA_signal_15187, new_AGEMA_signal_15186, new_AGEMA_signal_15185, mcs1_mcs_mat1_5_mcs_out[117]}), .c ({new_AGEMA_signal_18463, new_AGEMA_signal_18462, new_AGEMA_signal_18461, mcs1_mcs_mat1_5_n108}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U63 ( .a ({new_AGEMA_signal_20635, new_AGEMA_signal_20634, new_AGEMA_signal_20633, mcs1_mcs_mat1_5_n106}), .b ({new_AGEMA_signal_16264, new_AGEMA_signal_16263, new_AGEMA_signal_16262, mcs1_mcs_mat1_5_n105}), .c ({new_AGEMA_signal_21283, new_AGEMA_signal_21282, new_AGEMA_signal_21281, mcs_out[232]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U62 ( .a ({new_AGEMA_signal_15178, new_AGEMA_signal_15177, new_AGEMA_signal_15176, mcs1_mcs_mat1_5_mcs_out[120]}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_16264, new_AGEMA_signal_16263, new_AGEMA_signal_16262, mcs1_mcs_mat1_5_n105}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U61 ( .a ({new_AGEMA_signal_19879, new_AGEMA_signal_19878, new_AGEMA_signal_19877, mcs1_mcs_mat1_5_mcs_out[112]}), .b ({new_AGEMA_signal_13747, new_AGEMA_signal_13746, new_AGEMA_signal_13745, mcs1_mcs_mat1_5_mcs_out[116]}), .c ({new_AGEMA_signal_20635, new_AGEMA_signal_20634, new_AGEMA_signal_20633, mcs1_mcs_mat1_5_n106}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U60 ( .a ({new_AGEMA_signal_16267, new_AGEMA_signal_16266, new_AGEMA_signal_16265, mcs1_mcs_mat1_5_n104}), .b ({new_AGEMA_signal_20638, new_AGEMA_signal_20637, new_AGEMA_signal_20636, mcs1_mcs_mat1_5_n103}), .c ({new_AGEMA_signal_21286, new_AGEMA_signal_21285, new_AGEMA_signal_21284, mcs_out[203]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U59 ( .a ({new_AGEMA_signal_16303, new_AGEMA_signal_16302, new_AGEMA_signal_16301, mcs1_mcs_mat1_5_mcs_out[111]}), .b ({new_AGEMA_signal_19882, new_AGEMA_signal_19881, new_AGEMA_signal_19880, mcs1_mcs_mat1_5_mcs_out[99]}), .c ({new_AGEMA_signal_20638, new_AGEMA_signal_20637, new_AGEMA_signal_20636, mcs1_mcs_mat1_5_n103}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U58 ( .a ({new_AGEMA_signal_15214, new_AGEMA_signal_15213, new_AGEMA_signal_15212, mcs1_mcs_mat1_5_mcs_out[103]}), .b ({new_AGEMA_signal_15202, new_AGEMA_signal_15201, new_AGEMA_signal_15200, mcs1_mcs_mat1_5_mcs_out[107]}), .c ({new_AGEMA_signal_16267, new_AGEMA_signal_16266, new_AGEMA_signal_16265, mcs1_mcs_mat1_5_n104}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U57 ( .a ({new_AGEMA_signal_16270, new_AGEMA_signal_16269, new_AGEMA_signal_16268, mcs1_mcs_mat1_5_n102}), .b ({new_AGEMA_signal_19129, new_AGEMA_signal_19128, new_AGEMA_signal_19127, mcs1_mcs_mat1_5_n101}), .c ({new_AGEMA_signal_19846, new_AGEMA_signal_19845, new_AGEMA_signal_19844, mcs_out[202]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U56 ( .a ({new_AGEMA_signal_16306, new_AGEMA_signal_16305, new_AGEMA_signal_16304, mcs1_mcs_mat1_5_mcs_out[110]}), .b ({new_AGEMA_signal_18487, new_AGEMA_signal_18486, new_AGEMA_signal_18485, mcs1_mcs_mat1_5_mcs_out[98]}), .c ({new_AGEMA_signal_19129, new_AGEMA_signal_19128, new_AGEMA_signal_19127, mcs1_mcs_mat1_5_n101}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U55 ( .a ({new_AGEMA_signal_12319, new_AGEMA_signal_12318, new_AGEMA_signal_12317, mcs1_mcs_mat1_5_mcs_out[102]}), .b ({new_AGEMA_signal_15205, new_AGEMA_signal_15204, new_AGEMA_signal_15203, mcs1_mcs_mat1_5_mcs_out[106]}), .c ({new_AGEMA_signal_16270, new_AGEMA_signal_16269, new_AGEMA_signal_16268, mcs1_mcs_mat1_5_n102}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U54 ( .a ({new_AGEMA_signal_16273, new_AGEMA_signal_16272, new_AGEMA_signal_16271, mcs1_mcs_mat1_5_n100}), .b ({new_AGEMA_signal_17803, new_AGEMA_signal_17802, new_AGEMA_signal_17801, mcs1_mcs_mat1_5_n99}), .c ({new_AGEMA_signal_18466, new_AGEMA_signal_18465, new_AGEMA_signal_18464, mcs_out[201]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U53 ( .a ({new_AGEMA_signal_16309, new_AGEMA_signal_16308, new_AGEMA_signal_16307, mcs1_mcs_mat1_5_mcs_out[109]}), .b ({new_AGEMA_signal_17152, new_AGEMA_signal_17151, new_AGEMA_signal_17150, mcs1_mcs_mat1_5_mcs_out[97]}), .c ({new_AGEMA_signal_17803, new_AGEMA_signal_17802, new_AGEMA_signal_17801, mcs1_mcs_mat1_5_n99}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U52 ( .a ({new_AGEMA_signal_13768, new_AGEMA_signal_13767, new_AGEMA_signal_13766, mcs1_mcs_mat1_5_mcs_out[101]}), .b ({new_AGEMA_signal_15208, new_AGEMA_signal_15207, new_AGEMA_signal_15206, mcs1_mcs_mat1_5_mcs_out[105]}), .c ({new_AGEMA_signal_16273, new_AGEMA_signal_16272, new_AGEMA_signal_16271, mcs1_mcs_mat1_5_n100}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U51 ( .a ({new_AGEMA_signal_17125, new_AGEMA_signal_17124, new_AGEMA_signal_17123, mcs1_mcs_mat1_5_n98}), .b ({new_AGEMA_signal_21697, new_AGEMA_signal_21696, new_AGEMA_signal_21695, mcs1_mcs_mat1_5_n97}), .c ({new_AGEMA_signal_21838, new_AGEMA_signal_21837, new_AGEMA_signal_21836, mcs_out[200]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U50 ( .a ({new_AGEMA_signal_16312, new_AGEMA_signal_16311, new_AGEMA_signal_16310, mcs1_mcs_mat1_5_mcs_out[108]}), .b ({new_AGEMA_signal_21295, new_AGEMA_signal_21294, new_AGEMA_signal_21293, mcs1_mcs_mat1_5_mcs_out[96]}), .c ({new_AGEMA_signal_21697, new_AGEMA_signal_21696, new_AGEMA_signal_21695, mcs1_mcs_mat1_5_n97}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U49 ( .a ({new_AGEMA_signal_15217, new_AGEMA_signal_15216, new_AGEMA_signal_15215, mcs1_mcs_mat1_5_mcs_out[100]}), .b ({new_AGEMA_signal_16315, new_AGEMA_signal_16314, new_AGEMA_signal_16313, mcs1_mcs_mat1_5_mcs_out[104]}), .c ({new_AGEMA_signal_17125, new_AGEMA_signal_17124, new_AGEMA_signal_17123, mcs1_mcs_mat1_5_n98}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U48 ( .a ({new_AGEMA_signal_19132, new_AGEMA_signal_19131, new_AGEMA_signal_19130, mcs1_mcs_mat1_5_n96}), .b ({new_AGEMA_signal_16276, new_AGEMA_signal_16275, new_AGEMA_signal_16274, mcs1_mcs_mat1_5_n95}), .c ({new_AGEMA_signal_19849, new_AGEMA_signal_19848, new_AGEMA_signal_19847, mcs_out[171]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U47 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_15226, new_AGEMA_signal_15225, new_AGEMA_signal_15224, mcs1_mcs_mat1_5_mcs_out[95]}), .c ({new_AGEMA_signal_16276, new_AGEMA_signal_16275, new_AGEMA_signal_16274, mcs1_mcs_mat1_5_n95}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U46 ( .a ({new_AGEMA_signal_18490, new_AGEMA_signal_18489, new_AGEMA_signal_18488, mcs1_mcs_mat1_5_mcs_out[83]}), .b ({new_AGEMA_signal_12340, new_AGEMA_signal_12339, new_AGEMA_signal_12338, mcs1_mcs_mat1_5_mcs_out[87]}), .c ({new_AGEMA_signal_19132, new_AGEMA_signal_19131, new_AGEMA_signal_19130, mcs1_mcs_mat1_5_n96}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U45 ( .a ({new_AGEMA_signal_19135, new_AGEMA_signal_19134, new_AGEMA_signal_19133, mcs1_mcs_mat1_5_n94}), .b ({new_AGEMA_signal_13732, new_AGEMA_signal_13731, new_AGEMA_signal_13730, mcs1_mcs_mat1_5_n93}), .c ({new_AGEMA_signal_19852, new_AGEMA_signal_19851, new_AGEMA_signal_19850, mcs_out[170]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U43 ( .a ({new_AGEMA_signal_18493, new_AGEMA_signal_18492, new_AGEMA_signal_18491, mcs1_mcs_mat1_5_mcs_out[82]}), .b ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_19135, new_AGEMA_signal_19134, new_AGEMA_signal_19133, mcs1_mcs_mat1_5_n94}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U42 ( .a ({new_AGEMA_signal_19138, new_AGEMA_signal_19137, new_AGEMA_signal_19136, mcs1_mcs_mat1_5_n92}), .b ({new_AGEMA_signal_13735, new_AGEMA_signal_13734, new_AGEMA_signal_13733, mcs1_mcs_mat1_5_n91}), .c ({new_AGEMA_signal_19855, new_AGEMA_signal_19854, new_AGEMA_signal_19853, mcs_out[169]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U41 ( .a ({new_AGEMA_signal_11074, new_AGEMA_signal_11073, new_AGEMA_signal_11072, mcs1_mcs_mat1_5_mcs_out[89]}), .b ({new_AGEMA_signal_12334, new_AGEMA_signal_12333, new_AGEMA_signal_12332, mcs1_mcs_mat1_5_mcs_out[93]}), .c ({new_AGEMA_signal_13735, new_AGEMA_signal_13734, new_AGEMA_signal_13733, mcs1_mcs_mat1_5_n91}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U40 ( .a ({new_AGEMA_signal_18496, new_AGEMA_signal_18495, new_AGEMA_signal_18494, mcs1_mcs_mat1_5_mcs_out[81]}), .b ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_19138, new_AGEMA_signal_19137, new_AGEMA_signal_19136, mcs1_mcs_mat1_5_n92}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U39 ( .a ({new_AGEMA_signal_19858, new_AGEMA_signal_19857, new_AGEMA_signal_19856, mcs1_mcs_mat1_5_n90}), .b ({new_AGEMA_signal_17128, new_AGEMA_signal_17127, new_AGEMA_signal_17126, mcs1_mcs_mat1_5_n89}), .c ({new_AGEMA_signal_20641, new_AGEMA_signal_20640, new_AGEMA_signal_20639, mcs_out[168]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U38 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_16318, new_AGEMA_signal_16317, new_AGEMA_signal_16316, mcs1_mcs_mat1_5_mcs_out[92]}), .c ({new_AGEMA_signal_17128, new_AGEMA_signal_17127, new_AGEMA_signal_17126, mcs1_mcs_mat1_5_n89}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U37 ( .a ({new_AGEMA_signal_19162, new_AGEMA_signal_19161, new_AGEMA_signal_19160, mcs1_mcs_mat1_5_mcs_out[80]}), .b ({new_AGEMA_signal_13780, new_AGEMA_signal_13779, new_AGEMA_signal_13778, mcs1_mcs_mat1_5_mcs_out[84]}), .c ({new_AGEMA_signal_19858, new_AGEMA_signal_19857, new_AGEMA_signal_19856, mcs1_mcs_mat1_5_n90}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U36 ( .a ({new_AGEMA_signal_19861, new_AGEMA_signal_19860, new_AGEMA_signal_19859, mcs1_mcs_mat1_5_n88}), .b ({new_AGEMA_signal_15160, new_AGEMA_signal_15159, new_AGEMA_signal_15158, mcs1_mcs_mat1_5_n87}), .c ({temp_next_s3[9], temp_next_s2[9], temp_next_s1[9], temp_next_s0[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U35 ( .a ({new_AGEMA_signal_11137, new_AGEMA_signal_11136, new_AGEMA_signal_11135, mcs1_mcs_mat1_5_mcs_out[5]}), .b ({new_AGEMA_signal_13891, new_AGEMA_signal_13890, new_AGEMA_signal_13889, mcs1_mcs_mat1_5_mcs_out[9]}), .c ({new_AGEMA_signal_15160, new_AGEMA_signal_15159, new_AGEMA_signal_15158, mcs1_mcs_mat1_5_n87}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U34 ( .a ({new_AGEMA_signal_15322, new_AGEMA_signal_15321, new_AGEMA_signal_15320, mcs1_mcs_mat1_5_mcs_out[13]}), .b ({new_AGEMA_signal_19180, new_AGEMA_signal_19179, new_AGEMA_signal_19178, mcs1_mcs_mat1_5_mcs_out[1]}), .c ({new_AGEMA_signal_19861, new_AGEMA_signal_19860, new_AGEMA_signal_19859, mcs1_mcs_mat1_5_n88}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U33 ( .a ({new_AGEMA_signal_20647, new_AGEMA_signal_20646, new_AGEMA_signal_20645, mcs1_mcs_mat1_5_n86}), .b ({new_AGEMA_signal_16279, new_AGEMA_signal_16278, new_AGEMA_signal_16277, mcs1_mcs_mat1_5_n85}), .c ({new_AGEMA_signal_21289, new_AGEMA_signal_21288, new_AGEMA_signal_21287, mcs_out[139]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U32 ( .a ({new_AGEMA_signal_12349, new_AGEMA_signal_12348, new_AGEMA_signal_12347, mcs1_mcs_mat1_5_mcs_out[75]}), .b ({new_AGEMA_signal_15235, new_AGEMA_signal_15234, new_AGEMA_signal_15233, mcs1_mcs_mat1_5_mcs_out[79]}), .c ({new_AGEMA_signal_16279, new_AGEMA_signal_16278, new_AGEMA_signal_16277, mcs1_mcs_mat1_5_n85}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U31 ( .a ({new_AGEMA_signal_19885, new_AGEMA_signal_19884, new_AGEMA_signal_19883, mcs1_mcs_mat1_5_mcs_out[67]}), .b ({new_AGEMA_signal_15247, new_AGEMA_signal_15246, new_AGEMA_signal_15245, mcs1_mcs_mat1_5_mcs_out[71]}), .c ({new_AGEMA_signal_20647, new_AGEMA_signal_20646, new_AGEMA_signal_20645, mcs1_mcs_mat1_5_n86}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U30 ( .a ({new_AGEMA_signal_19864, new_AGEMA_signal_19863, new_AGEMA_signal_19862, mcs1_mcs_mat1_5_n84}), .b ({new_AGEMA_signal_17131, new_AGEMA_signal_17130, new_AGEMA_signal_17129, mcs1_mcs_mat1_5_n83}), .c ({new_AGEMA_signal_20650, new_AGEMA_signal_20649, new_AGEMA_signal_20648, mcs_out[138]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U29 ( .a ({new_AGEMA_signal_16324, new_AGEMA_signal_16323, new_AGEMA_signal_16322, mcs1_mcs_mat1_5_mcs_out[74]}), .b ({new_AGEMA_signal_9832, new_AGEMA_signal_9831, new_AGEMA_signal_9830, mcs1_mcs_mat1_5_mcs_out[78]}), .c ({new_AGEMA_signal_17131, new_AGEMA_signal_17130, new_AGEMA_signal_17129, mcs1_mcs_mat1_5_n83}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U28 ( .a ({new_AGEMA_signal_19165, new_AGEMA_signal_19164, new_AGEMA_signal_19163, mcs1_mcs_mat1_5_mcs_out[66]}), .b ({new_AGEMA_signal_16330, new_AGEMA_signal_16329, new_AGEMA_signal_16328, mcs1_mcs_mat1_5_mcs_out[70]}), .c ({new_AGEMA_signal_19864, new_AGEMA_signal_19863, new_AGEMA_signal_19862, mcs1_mcs_mat1_5_n84}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U27 ( .a ({new_AGEMA_signal_18469, new_AGEMA_signal_18468, new_AGEMA_signal_18467, mcs1_mcs_mat1_5_n82}), .b ({new_AGEMA_signal_15163, new_AGEMA_signal_15162, new_AGEMA_signal_15161, mcs1_mcs_mat1_5_n81}), .c ({new_AGEMA_signal_19141, new_AGEMA_signal_19140, new_AGEMA_signal_19139, mcs_out[137]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U26 ( .a ({new_AGEMA_signal_13789, new_AGEMA_signal_13788, new_AGEMA_signal_13787, mcs1_mcs_mat1_5_mcs_out[73]}), .b ({new_AGEMA_signal_12343, new_AGEMA_signal_12342, new_AGEMA_signal_12341, mcs1_mcs_mat1_5_mcs_out[77]}), .c ({new_AGEMA_signal_15163, new_AGEMA_signal_15162, new_AGEMA_signal_15161, mcs1_mcs_mat1_5_n81}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U25 ( .a ({new_AGEMA_signal_17836, new_AGEMA_signal_17835, new_AGEMA_signal_17834, mcs1_mcs_mat1_5_mcs_out[65]}), .b ({new_AGEMA_signal_16333, new_AGEMA_signal_16332, new_AGEMA_signal_16331, mcs1_mcs_mat1_5_mcs_out[69]}), .c ({new_AGEMA_signal_18469, new_AGEMA_signal_18468, new_AGEMA_signal_18467, mcs1_mcs_mat1_5_n82}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U24 ( .a ({new_AGEMA_signal_21292, new_AGEMA_signal_21291, new_AGEMA_signal_21290, mcs1_mcs_mat1_5_n80}), .b ({new_AGEMA_signal_17134, new_AGEMA_signal_17133, new_AGEMA_signal_17132, mcs1_mcs_mat1_5_n79}), .c ({new_AGEMA_signal_21700, new_AGEMA_signal_21699, new_AGEMA_signal_21698, mcs_out[136]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U23 ( .a ({new_AGEMA_signal_16327, new_AGEMA_signal_16326, new_AGEMA_signal_16325, mcs1_mcs_mat1_5_mcs_out[72]}), .b ({new_AGEMA_signal_16321, new_AGEMA_signal_16320, new_AGEMA_signal_16319, mcs1_mcs_mat1_5_mcs_out[76]}), .c ({new_AGEMA_signal_17134, new_AGEMA_signal_17133, new_AGEMA_signal_17132, mcs1_mcs_mat1_5_n79}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U22 ( .a ({new_AGEMA_signal_20662, new_AGEMA_signal_20661, new_AGEMA_signal_20660, mcs1_mcs_mat1_5_mcs_out[64]}), .b ({new_AGEMA_signal_15253, new_AGEMA_signal_15252, new_AGEMA_signal_15251, mcs1_mcs_mat1_5_mcs_out[68]}), .c ({new_AGEMA_signal_21292, new_AGEMA_signal_21291, new_AGEMA_signal_21290, mcs1_mcs_mat1_5_n80}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U21 ( .a ({new_AGEMA_signal_18472, new_AGEMA_signal_18471, new_AGEMA_signal_18470, mcs1_mcs_mat1_5_n78}), .b ({new_AGEMA_signal_16282, new_AGEMA_signal_16281, new_AGEMA_signal_16280, mcs1_mcs_mat1_5_n77}), .c ({temp_next_s3[107], temp_next_s2[107], temp_next_s1[107], temp_next_s0[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U20 ( .a ({new_AGEMA_signal_13813, new_AGEMA_signal_13812, new_AGEMA_signal_13811, mcs1_mcs_mat1_5_mcs_out[59]}), .b ({new_AGEMA_signal_15259, new_AGEMA_signal_15258, new_AGEMA_signal_15257, mcs1_mcs_mat1_5_mcs_out[63]}), .c ({new_AGEMA_signal_16282, new_AGEMA_signal_16281, new_AGEMA_signal_16280, mcs1_mcs_mat1_5_n77}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U19 ( .a ({new_AGEMA_signal_17842, new_AGEMA_signal_17841, new_AGEMA_signal_17840, mcs1_mcs_mat1_5_mcs_out[51]}), .b ({new_AGEMA_signal_15268, new_AGEMA_signal_15267, new_AGEMA_signal_15266, mcs1_mcs_mat1_5_mcs_out[55]}), .c ({new_AGEMA_signal_18472, new_AGEMA_signal_18471, new_AGEMA_signal_18470, mcs1_mcs_mat1_5_n78}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U18 ( .a ({new_AGEMA_signal_17137, new_AGEMA_signal_17136, new_AGEMA_signal_17135, mcs1_mcs_mat1_5_n76}), .b ({new_AGEMA_signal_15166, new_AGEMA_signal_15165, new_AGEMA_signal_15164, mcs1_mcs_mat1_5_n75}), .c ({temp_next_s3[106], temp_next_s2[106], temp_next_s1[106], temp_next_s0[106]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U17 ( .a ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, new_AGEMA_signal_12371, mcs1_mcs_mat1_5_mcs_out[58]}), .b ({new_AGEMA_signal_13804, new_AGEMA_signal_13803, new_AGEMA_signal_13802, mcs1_mcs_mat1_5_mcs_out[62]}), .c ({new_AGEMA_signal_15166, new_AGEMA_signal_15165, new_AGEMA_signal_15164, mcs1_mcs_mat1_5_n75}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U16 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_16339, new_AGEMA_signal_16338, new_AGEMA_signal_16337, mcs1_mcs_mat1_5_mcs_out[54]}), .c ({new_AGEMA_signal_17137, new_AGEMA_signal_17136, new_AGEMA_signal_17135, mcs1_mcs_mat1_5_n76}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U15 ( .a ({new_AGEMA_signal_17140, new_AGEMA_signal_17139, new_AGEMA_signal_17138, mcs1_mcs_mat1_5_n74}), .b ({new_AGEMA_signal_15169, new_AGEMA_signal_15168, new_AGEMA_signal_15167, mcs1_mcs_mat1_5_n73}), .c ({temp_next_s3[105], temp_next_s2[105], temp_next_s1[105], temp_next_s0[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U14 ( .a ({new_AGEMA_signal_13816, new_AGEMA_signal_13815, new_AGEMA_signal_13814, mcs1_mcs_mat1_5_mcs_out[57]}), .b ({new_AGEMA_signal_13807, new_AGEMA_signal_13806, new_AGEMA_signal_13805, mcs1_mcs_mat1_5_mcs_out[61]}), .c ({new_AGEMA_signal_15169, new_AGEMA_signal_15168, new_AGEMA_signal_15167, mcs1_mcs_mat1_5_n73}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U13 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({new_AGEMA_signal_16342, new_AGEMA_signal_16341, new_AGEMA_signal_16340, mcs1_mcs_mat1_5_mcs_out[53]}), .c ({new_AGEMA_signal_17140, new_AGEMA_signal_17139, new_AGEMA_signal_17138, mcs1_mcs_mat1_5_n74}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U12 ( .a ({new_AGEMA_signal_19147, new_AGEMA_signal_19146, new_AGEMA_signal_19145, mcs1_mcs_mat1_5_n72}), .b ({new_AGEMA_signal_17143, new_AGEMA_signal_17142, new_AGEMA_signal_17141, mcs1_mcs_mat1_5_n71}), .c ({temp_next_s3[104], temp_next_s2[104], temp_next_s1[104], temp_next_s0[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U11 ( .a ({new_AGEMA_signal_15265, new_AGEMA_signal_15264, new_AGEMA_signal_15263, mcs1_mcs_mat1_5_mcs_out[56]}), .b ({new_AGEMA_signal_16336, new_AGEMA_signal_16335, new_AGEMA_signal_16334, mcs1_mcs_mat1_5_mcs_out[60]}), .c ({new_AGEMA_signal_17143, new_AGEMA_signal_17142, new_AGEMA_signal_17141, mcs1_mcs_mat1_5_n71}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U10 ( .a ({new_AGEMA_signal_18505, new_AGEMA_signal_18504, new_AGEMA_signal_18503, mcs1_mcs_mat1_5_mcs_out[48]}), .b ({new_AGEMA_signal_15274, new_AGEMA_signal_15273, new_AGEMA_signal_15272, mcs1_mcs_mat1_5_mcs_out[52]}), .c ({new_AGEMA_signal_19147, new_AGEMA_signal_19146, new_AGEMA_signal_19145, mcs1_mcs_mat1_5_n72}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U9 ( .a ({new_AGEMA_signal_19870, new_AGEMA_signal_19869, new_AGEMA_signal_19868, mcs1_mcs_mat1_5_n70}), .b ({new_AGEMA_signal_16285, new_AGEMA_signal_16284, new_AGEMA_signal_16283, mcs1_mcs_mat1_5_n69}), .c ({temp_next_s3[75], temp_next_s2[75], temp_next_s1[75], temp_next_s0[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U8 ( .a ({new_AGEMA_signal_15280, new_AGEMA_signal_15279, new_AGEMA_signal_15278, mcs1_mcs_mat1_5_mcs_out[43]}), .b ({new_AGEMA_signal_15277, new_AGEMA_signal_15276, new_AGEMA_signal_15275, mcs1_mcs_mat1_5_mcs_out[47]}), .c ({new_AGEMA_signal_16285, new_AGEMA_signal_16284, new_AGEMA_signal_16283, mcs1_mcs_mat1_5_n69}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U7 ( .a ({new_AGEMA_signal_19171, new_AGEMA_signal_19170, new_AGEMA_signal_19169, mcs1_mcs_mat1_5_mcs_out[35]}), .b ({new_AGEMA_signal_16348, new_AGEMA_signal_16347, new_AGEMA_signal_16346, mcs1_mcs_mat1_5_mcs_out[39]}), .c ({new_AGEMA_signal_19870, new_AGEMA_signal_19869, new_AGEMA_signal_19868, mcs1_mcs_mat1_5_n70}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U6 ( .a ({new_AGEMA_signal_19150, new_AGEMA_signal_19149, new_AGEMA_signal_19148, mcs1_mcs_mat1_5_n68}), .b ({new_AGEMA_signal_16288, new_AGEMA_signal_16287, new_AGEMA_signal_16286, mcs1_mcs_mat1_5_n67}), .c ({temp_next_s3[74], temp_next_s2[74], temp_next_s1[74], temp_next_s0[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U5 ( .a ({new_AGEMA_signal_15283, new_AGEMA_signal_15282, new_AGEMA_signal_15281, mcs1_mcs_mat1_5_mcs_out[42]}), .b ({new_AGEMA_signal_11098, new_AGEMA_signal_11097, new_AGEMA_signal_11096, mcs1_mcs_mat1_5_mcs_out[46]}), .c ({new_AGEMA_signal_16288, new_AGEMA_signal_16287, new_AGEMA_signal_16286, mcs1_mcs_mat1_5_n67}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U4 ( .a ({new_AGEMA_signal_18508, new_AGEMA_signal_18507, new_AGEMA_signal_18506, mcs1_mcs_mat1_5_mcs_out[34]}), .b ({new_AGEMA_signal_12412, new_AGEMA_signal_12411, new_AGEMA_signal_12410, mcs1_mcs_mat1_5_mcs_out[38]}), .c ({new_AGEMA_signal_19150, new_AGEMA_signal_19149, new_AGEMA_signal_19148, mcs1_mcs_mat1_5_n68}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U3 ( .a ({new_AGEMA_signal_19876, new_AGEMA_signal_19875, new_AGEMA_signal_19874, mcs1_mcs_mat1_5_n66}), .b ({new_AGEMA_signal_18475, new_AGEMA_signal_18474, new_AGEMA_signal_18473, mcs1_mcs_mat1_5_n65}), .c ({temp_next_s3[8], temp_next_s2[8], temp_next_s1[8], temp_next_s0[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U2 ( .a ({new_AGEMA_signal_17863, new_AGEMA_signal_17862, new_AGEMA_signal_17861, mcs1_mcs_mat1_5_mcs_out[4]}), .b ({new_AGEMA_signal_16375, new_AGEMA_signal_16374, new_AGEMA_signal_16373, mcs1_mcs_mat1_5_mcs_out[8]}), .c ({new_AGEMA_signal_18475, new_AGEMA_signal_18474, new_AGEMA_signal_18473, mcs1_mcs_mat1_5_n65}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_U1 ( .a ({new_AGEMA_signal_19183, new_AGEMA_signal_19182, new_AGEMA_signal_19181, mcs1_mcs_mat1_5_mcs_out[0]}), .b ({new_AGEMA_signal_17176, new_AGEMA_signal_17175, new_AGEMA_signal_17174, mcs1_mcs_mat1_5_mcs_out[12]}), .c ({new_AGEMA_signal_19876, new_AGEMA_signal_19875, new_AGEMA_signal_19874, mcs1_mcs_mat1_5_n66}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_15172, new_AGEMA_signal_15171, new_AGEMA_signal_15170, mcs1_mcs_mat1_5_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_16291, new_AGEMA_signal_16290, new_AGEMA_signal_16289, mcs1_mcs_mat1_5_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_13738, new_AGEMA_signal_13737, new_AGEMA_signal_13736, mcs1_mcs_mat1_5_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_8953, new_AGEMA_signal_8952, new_AGEMA_signal_8951, mcs1_mcs_mat1_5_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_15172, new_AGEMA_signal_15171, new_AGEMA_signal_15170, mcs1_mcs_mat1_5_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_9811, new_AGEMA_signal_9810, new_AGEMA_signal_9809, mcs1_mcs_mat1_5_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_11032, new_AGEMA_signal_11031, new_AGEMA_signal_11030, mcs1_mcs_mat1_5_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_12292, new_AGEMA_signal_12291, new_AGEMA_signal_12290, mcs1_mcs_mat1_5_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_9814, new_AGEMA_signal_9813, new_AGEMA_signal_9812, mcs1_mcs_mat1_5_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .c ({new_AGEMA_signal_11032, new_AGEMA_signal_11031, new_AGEMA_signal_11030, mcs1_mcs_mat1_5_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_15175, new_AGEMA_signal_15174, new_AGEMA_signal_15173, mcs1_mcs_mat1_5_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .c ({new_AGEMA_signal_16294, new_AGEMA_signal_16293, new_AGEMA_signal_16292, mcs1_mcs_mat1_5_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_13738, new_AGEMA_signal_13737, new_AGEMA_signal_13736, mcs1_mcs_mat1_5_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_15175, new_AGEMA_signal_15174, new_AGEMA_signal_15173, mcs1_mcs_mat1_5_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_12295, new_AGEMA_signal_12294, new_AGEMA_signal_12293, mcs1_mcs_mat1_5_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_11035, new_AGEMA_signal_11034, new_AGEMA_signal_11033, mcs1_mcs_mat1_5_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_13738, new_AGEMA_signal_13737, new_AGEMA_signal_13736, mcs1_mcs_mat1_5_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_13741, new_AGEMA_signal_13740, new_AGEMA_signal_13739, mcs1_mcs_mat1_5_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_15178, new_AGEMA_signal_15177, new_AGEMA_signal_15176, mcs1_mcs_mat1_5_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_12295, new_AGEMA_signal_12294, new_AGEMA_signal_12293, mcs1_mcs_mat1_5_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9814, new_AGEMA_signal_9813, new_AGEMA_signal_9812, mcs1_mcs_mat1_5_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_13741, new_AGEMA_signal_13740, new_AGEMA_signal_13739, mcs1_mcs_mat1_5_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5213], Fresh[5212], Fresh[5211], Fresh[5210], Fresh[5209], Fresh[5208]}), .c ({new_AGEMA_signal_12295, new_AGEMA_signal_12294, new_AGEMA_signal_12293, mcs1_mcs_mat1_5_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5219], Fresh[5218], Fresh[5217], Fresh[5216], Fresh[5215], Fresh[5214]}), .c ({new_AGEMA_signal_9814, new_AGEMA_signal_9813, new_AGEMA_signal_9812, mcs1_mcs_mat1_5_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5225], Fresh[5224], Fresh[5223], Fresh[5222], Fresh[5221], Fresh[5220]}), .c ({new_AGEMA_signal_11035, new_AGEMA_signal_11034, new_AGEMA_signal_11033, mcs1_mcs_mat1_5_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_15181, new_AGEMA_signal_15180, new_AGEMA_signal_15179, mcs1_mcs_mat1_5_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .c ({new_AGEMA_signal_16297, new_AGEMA_signal_16296, new_AGEMA_signal_16295, mcs1_mcs_mat1_5_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_13744, new_AGEMA_signal_13743, new_AGEMA_signal_13742, mcs1_mcs_mat1_5_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_11044, new_AGEMA_signal_11043, new_AGEMA_signal_11042, mcs1_mcs_mat1_5_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_15181, new_AGEMA_signal_15180, new_AGEMA_signal_15179, mcs1_mcs_mat1_5_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_15184, new_AGEMA_signal_15183, new_AGEMA_signal_15182, mcs1_mcs_mat1_5_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_12301, new_AGEMA_signal_12300, new_AGEMA_signal_12299, mcs1_mcs_mat1_5_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_16300, new_AGEMA_signal_16299, new_AGEMA_signal_16298, mcs1_mcs_mat1_5_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_13744, new_AGEMA_signal_13743, new_AGEMA_signal_13742, mcs1_mcs_mat1_5_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .c ({new_AGEMA_signal_15184, new_AGEMA_signal_15183, new_AGEMA_signal_15182, mcs1_mcs_mat1_5_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_13744, new_AGEMA_signal_13743, new_AGEMA_signal_13742, mcs1_mcs_mat1_5_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_12298, new_AGEMA_signal_12297, new_AGEMA_signal_12296, mcs1_mcs_mat1_5_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_15187, new_AGEMA_signal_15186, new_AGEMA_signal_15185, mcs1_mcs_mat1_5_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_12304, new_AGEMA_signal_12303, new_AGEMA_signal_12302, mcs1_mcs_mat1_5_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_9817, new_AGEMA_signal_9816, new_AGEMA_signal_9815, mcs1_mcs_mat1_5_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_13744, new_AGEMA_signal_13743, new_AGEMA_signal_13742, mcs1_mcs_mat1_5_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_11041, new_AGEMA_signal_11040, new_AGEMA_signal_11039, mcs1_mcs_mat1_5_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_12301, new_AGEMA_signal_12300, new_AGEMA_signal_12299, mcs1_mcs_mat1_5_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_13747, new_AGEMA_signal_13746, new_AGEMA_signal_13745, mcs1_mcs_mat1_5_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_8956, new_AGEMA_signal_8955, new_AGEMA_signal_8954, mcs1_mcs_mat1_5_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_11044, new_AGEMA_signal_11043, new_AGEMA_signal_11042, mcs1_mcs_mat1_5_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_12301, new_AGEMA_signal_12300, new_AGEMA_signal_12299, mcs1_mcs_mat1_5_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_9817, new_AGEMA_signal_9816, new_AGEMA_signal_9815, mcs1_mcs_mat1_5_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_11041, new_AGEMA_signal_11040, new_AGEMA_signal_11039, mcs1_mcs_mat1_5_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5231], Fresh[5230], Fresh[5229], Fresh[5228], Fresh[5227], Fresh[5226]}), .c ({new_AGEMA_signal_12304, new_AGEMA_signal_12303, new_AGEMA_signal_12302, mcs1_mcs_mat1_5_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5237], Fresh[5236], Fresh[5235], Fresh[5234], Fresh[5233], Fresh[5232]}), .c ({new_AGEMA_signal_9817, new_AGEMA_signal_9816, new_AGEMA_signal_9815, mcs1_mcs_mat1_5_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5243], Fresh[5242], Fresh[5241], Fresh[5240], Fresh[5239], Fresh[5238]}), .c ({new_AGEMA_signal_11044, new_AGEMA_signal_11043, new_AGEMA_signal_11042, mcs1_mcs_mat1_5_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_18481, new_AGEMA_signal_18480, new_AGEMA_signal_18479, mcs1_mcs_mat1_5_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_15190, new_AGEMA_signal_15189, new_AGEMA_signal_15188, mcs1_mcs_mat1_5_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_19153, new_AGEMA_signal_19152, new_AGEMA_signal_19151, mcs1_mcs_mat1_5_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_17146, new_AGEMA_signal_17145, new_AGEMA_signal_17144, mcs1_mcs_mat1_5_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_17149, new_AGEMA_signal_17148, new_AGEMA_signal_17147, mcs1_mcs_mat1_5_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_17812, new_AGEMA_signal_17811, new_AGEMA_signal_17810, mcs1_mcs_mat1_5_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_18484, new_AGEMA_signal_18483, new_AGEMA_signal_18482, mcs1_mcs_mat1_5_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_19156, new_AGEMA_signal_19155, new_AGEMA_signal_19154, mcs1_mcs_mat1_5_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_19879, new_AGEMA_signal_19878, new_AGEMA_signal_19877, mcs1_mcs_mat1_5_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_18481, new_AGEMA_signal_18480, new_AGEMA_signal_18479, mcs1_mcs_mat1_5_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_19156, new_AGEMA_signal_19155, new_AGEMA_signal_19154, mcs1_mcs_mat1_5_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_13750, new_AGEMA_signal_13749, new_AGEMA_signal_13748, mcs1_mcs_mat1_5_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_17818, new_AGEMA_signal_17817, new_AGEMA_signal_17816, mcs1_mcs_mat1_5_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_18481, new_AGEMA_signal_18480, new_AGEMA_signal_18479, mcs1_mcs_mat1_5_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_15193, new_AGEMA_signal_15192, new_AGEMA_signal_15191, mcs1_mcs_mat1_5_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_17815, new_AGEMA_signal_17814, new_AGEMA_signal_17813, mcs1_mcs_mat1_5_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_18484, new_AGEMA_signal_18483, new_AGEMA_signal_18482, mcs1_mcs_mat1_5_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5249], Fresh[5248], Fresh[5247], Fresh[5246], Fresh[5245], Fresh[5244]}), .c ({new_AGEMA_signal_17818, new_AGEMA_signal_17817, new_AGEMA_signal_17816, mcs1_mcs_mat1_5_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5255], Fresh[5254], Fresh[5253], Fresh[5252], Fresh[5251], Fresh[5250]}), .c ({new_AGEMA_signal_15193, new_AGEMA_signal_15192, new_AGEMA_signal_15191, mcs1_mcs_mat1_5_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5261], Fresh[5260], Fresh[5259], Fresh[5258], Fresh[5257], Fresh[5256]}), .c ({new_AGEMA_signal_17149, new_AGEMA_signal_17148, new_AGEMA_signal_17147, mcs1_mcs_mat1_5_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({new_AGEMA_signal_15196, new_AGEMA_signal_15195, new_AGEMA_signal_15194, mcs1_mcs_mat1_5_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_16303, new_AGEMA_signal_16302, new_AGEMA_signal_16301, mcs1_mcs_mat1_5_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({new_AGEMA_signal_15199, new_AGEMA_signal_15198, new_AGEMA_signal_15197, mcs1_mcs_mat1_5_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_16306, new_AGEMA_signal_16305, new_AGEMA_signal_16304, mcs1_mcs_mat1_5_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_11047, new_AGEMA_signal_11046, new_AGEMA_signal_11045, mcs1_mcs_mat1_5_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_15196, new_AGEMA_signal_15195, new_AGEMA_signal_15194, mcs1_mcs_mat1_5_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_16309, new_AGEMA_signal_16308, new_AGEMA_signal_16307, mcs1_mcs_mat1_5_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_9820, new_AGEMA_signal_9819, new_AGEMA_signal_9818, mcs1_mcs_mat1_5_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_13753, new_AGEMA_signal_13752, new_AGEMA_signal_13751, mcs1_mcs_mat1_5_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_15196, new_AGEMA_signal_15195, new_AGEMA_signal_15194, mcs1_mcs_mat1_5_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_12307, new_AGEMA_signal_12306, new_AGEMA_signal_12305, mcs1_mcs_mat1_5_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_15199, new_AGEMA_signal_15198, new_AGEMA_signal_15197, mcs1_mcs_mat1_5_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_16312, new_AGEMA_signal_16311, new_AGEMA_signal_16310, mcs1_mcs_mat1_5_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_13756, new_AGEMA_signal_13755, new_AGEMA_signal_13754, mcs1_mcs_mat1_5_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_15199, new_AGEMA_signal_15198, new_AGEMA_signal_15197, mcs1_mcs_mat1_5_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_11047, new_AGEMA_signal_11046, new_AGEMA_signal_11045, mcs1_mcs_mat1_5_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_12310, new_AGEMA_signal_12309, new_AGEMA_signal_12308, mcs1_mcs_mat1_5_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_13756, new_AGEMA_signal_13755, new_AGEMA_signal_13754, mcs1_mcs_mat1_5_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5267], Fresh[5266], Fresh[5265], Fresh[5264], Fresh[5263], Fresh[5262]}), .c ({new_AGEMA_signal_12310, new_AGEMA_signal_12309, new_AGEMA_signal_12308, mcs1_mcs_mat1_5_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5273], Fresh[5272], Fresh[5271], Fresh[5270], Fresh[5269], Fresh[5268]}), .c ({new_AGEMA_signal_9820, new_AGEMA_signal_9819, new_AGEMA_signal_9818, mcs1_mcs_mat1_5_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5279], Fresh[5278], Fresh[5277], Fresh[5276], Fresh[5275], Fresh[5274]}), .c ({new_AGEMA_signal_11047, new_AGEMA_signal_11046, new_AGEMA_signal_11045, mcs1_mcs_mat1_5_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_13762, new_AGEMA_signal_13761, new_AGEMA_signal_13760, mcs1_mcs_mat1_5_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_13759, new_AGEMA_signal_13758, new_AGEMA_signal_13757, mcs1_mcs_mat1_5_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_15202, new_AGEMA_signal_15201, new_AGEMA_signal_15200, mcs1_mcs_mat1_5_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_13759, new_AGEMA_signal_13758, new_AGEMA_signal_13757, mcs1_mcs_mat1_5_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_11050, new_AGEMA_signal_11049, new_AGEMA_signal_11048, mcs1_mcs_mat1_5_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_15205, new_AGEMA_signal_15204, new_AGEMA_signal_15203, mcs1_mcs_mat1_5_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_9823, new_AGEMA_signal_9822, new_AGEMA_signal_9821, mcs1_mcs_mat1_5_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .c ({new_AGEMA_signal_11050, new_AGEMA_signal_11049, new_AGEMA_signal_11048, mcs1_mcs_mat1_5_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({new_AGEMA_signal_13759, new_AGEMA_signal_13758, new_AGEMA_signal_13757, mcs1_mcs_mat1_5_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_15208, new_AGEMA_signal_15207, new_AGEMA_signal_15206, mcs1_mcs_mat1_5_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_12316, new_AGEMA_signal_12315, new_AGEMA_signal_12314, mcs1_mcs_mat1_5_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_8962, new_AGEMA_signal_8961, new_AGEMA_signal_8960, mcs1_mcs_mat1_5_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_13759, new_AGEMA_signal_13758, new_AGEMA_signal_13757, mcs1_mcs_mat1_5_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_15211, new_AGEMA_signal_15210, new_AGEMA_signal_15209, mcs1_mcs_mat1_5_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_16315, new_AGEMA_signal_16314, new_AGEMA_signal_16313, mcs1_mcs_mat1_5_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_13762, new_AGEMA_signal_13761, new_AGEMA_signal_13760, mcs1_mcs_mat1_5_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_12316, new_AGEMA_signal_12315, new_AGEMA_signal_12314, mcs1_mcs_mat1_5_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_15211, new_AGEMA_signal_15210, new_AGEMA_signal_15209, mcs1_mcs_mat1_5_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_12313, new_AGEMA_signal_12312, new_AGEMA_signal_12311, mcs1_mcs_mat1_5_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .c ({new_AGEMA_signal_13762, new_AGEMA_signal_13761, new_AGEMA_signal_13760, mcs1_mcs_mat1_5_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_9823, new_AGEMA_signal_9822, new_AGEMA_signal_9821, mcs1_mcs_mat1_5_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_11053, new_AGEMA_signal_11052, new_AGEMA_signal_11051, mcs1_mcs_mat1_5_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_12313, new_AGEMA_signal_12312, new_AGEMA_signal_12311, mcs1_mcs_mat1_5_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5285], Fresh[5284], Fresh[5283], Fresh[5282], Fresh[5281], Fresh[5280]}), .c ({new_AGEMA_signal_12316, new_AGEMA_signal_12315, new_AGEMA_signal_12314, mcs1_mcs_mat1_5_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5291], Fresh[5290], Fresh[5289], Fresh[5288], Fresh[5287], Fresh[5286]}), .c ({new_AGEMA_signal_9823, new_AGEMA_signal_9822, new_AGEMA_signal_9821, mcs1_mcs_mat1_5_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5297], Fresh[5296], Fresh[5295], Fresh[5294], Fresh[5293], Fresh[5292]}), .c ({new_AGEMA_signal_11053, new_AGEMA_signal_11052, new_AGEMA_signal_11051, mcs1_mcs_mat1_5_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_11056, new_AGEMA_signal_11055, new_AGEMA_signal_11054, mcs1_mcs_mat1_5_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_13765, new_AGEMA_signal_13764, new_AGEMA_signal_13763, mcs1_mcs_mat1_5_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_15214, new_AGEMA_signal_15213, new_AGEMA_signal_15212, mcs1_mcs_mat1_5_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_12328, new_AGEMA_signal_12327, new_AGEMA_signal_12326, mcs1_mcs_mat1_5_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_13765, new_AGEMA_signal_13764, new_AGEMA_signal_13763, mcs1_mcs_mat1_5_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_12322, new_AGEMA_signal_12321, new_AGEMA_signal_12320, mcs1_mcs_mat1_5_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_11059, new_AGEMA_signal_11058, new_AGEMA_signal_11057, mcs1_mcs_mat1_5_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_13768, new_AGEMA_signal_13767, new_AGEMA_signal_13766, mcs1_mcs_mat1_5_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_12325, new_AGEMA_signal_12324, new_AGEMA_signal_12323, mcs1_mcs_mat1_5_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_13771, new_AGEMA_signal_13770, new_AGEMA_signal_13769, mcs1_mcs_mat1_5_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_15217, new_AGEMA_signal_15216, new_AGEMA_signal_15215, mcs1_mcs_mat1_5_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_8965, new_AGEMA_signal_8964, new_AGEMA_signal_8963, mcs1_mcs_mat1_5_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_12328, new_AGEMA_signal_12327, new_AGEMA_signal_12326, mcs1_mcs_mat1_5_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_13771, new_AGEMA_signal_13770, new_AGEMA_signal_13769, mcs1_mcs_mat1_5_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, new_AGEMA_signal_9824, mcs1_mcs_mat1_5_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .c ({new_AGEMA_signal_12325, new_AGEMA_signal_12324, new_AGEMA_signal_12323, mcs1_mcs_mat1_5_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5303], Fresh[5302], Fresh[5301], Fresh[5300], Fresh[5299], Fresh[5298]}), .c ({new_AGEMA_signal_12328, new_AGEMA_signal_12327, new_AGEMA_signal_12326, mcs1_mcs_mat1_5_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5309], Fresh[5308], Fresh[5307], Fresh[5306], Fresh[5305], Fresh[5304]}), .c ({new_AGEMA_signal_9826, new_AGEMA_signal_9825, new_AGEMA_signal_9824, mcs1_mcs_mat1_5_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5315], Fresh[5314], Fresh[5313], Fresh[5312], Fresh[5311], Fresh[5310]}), .c ({new_AGEMA_signal_11059, new_AGEMA_signal_11058, new_AGEMA_signal_11057, mcs1_mcs_mat1_5_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_20659, new_AGEMA_signal_20658, new_AGEMA_signal_20657, mcs1_mcs_mat1_5_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_17155, new_AGEMA_signal_17154, new_AGEMA_signal_17153, mcs1_mcs_mat1_5_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_21295, new_AGEMA_signal_21294, new_AGEMA_signal_21293, mcs1_mcs_mat1_5_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_19882, new_AGEMA_signal_19881, new_AGEMA_signal_19880, mcs1_mcs_mat1_5_mcs_out[99]}), .b ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .c ({new_AGEMA_signal_20659, new_AGEMA_signal_20658, new_AGEMA_signal_20657, mcs1_mcs_mat1_5_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_19159, new_AGEMA_signal_19158, new_AGEMA_signal_19157, mcs1_mcs_mat1_5_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .c ({new_AGEMA_signal_19882, new_AGEMA_signal_19881, new_AGEMA_signal_19880, mcs1_mcs_mat1_5_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_18487, new_AGEMA_signal_18486, new_AGEMA_signal_18485, mcs1_mcs_mat1_5_mcs_out[98]}), .b ({new_AGEMA_signal_15223, new_AGEMA_signal_15222, new_AGEMA_signal_15221, mcs1_mcs_mat1_5_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_19159, new_AGEMA_signal_19158, new_AGEMA_signal_19157, mcs1_mcs_mat1_5_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_15220, new_AGEMA_signal_15219, new_AGEMA_signal_15218, mcs1_mcs_mat1_5_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_17821, new_AGEMA_signal_17820, new_AGEMA_signal_17819, mcs1_mcs_mat1_5_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_18487, new_AGEMA_signal_18486, new_AGEMA_signal_18485, mcs1_mcs_mat1_5_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5321], Fresh[5320], Fresh[5319], Fresh[5318], Fresh[5317], Fresh[5316]}), .c ({new_AGEMA_signal_17821, new_AGEMA_signal_17820, new_AGEMA_signal_17819, mcs1_mcs_mat1_5_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5327], Fresh[5326], Fresh[5325], Fresh[5324], Fresh[5323], Fresh[5322]}), .c ({new_AGEMA_signal_15223, new_AGEMA_signal_15222, new_AGEMA_signal_15221, mcs1_mcs_mat1_5_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5333], Fresh[5332], Fresh[5331], Fresh[5330], Fresh[5329], Fresh[5328]}), .c ({new_AGEMA_signal_17155, new_AGEMA_signal_17154, new_AGEMA_signal_17153, mcs1_mcs_mat1_5_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_13777, new_AGEMA_signal_13776, new_AGEMA_signal_13775, mcs1_mcs_mat1_5_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_15226, new_AGEMA_signal_15225, new_AGEMA_signal_15224, mcs1_mcs_mat1_5_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_11065, new_AGEMA_signal_11064, new_AGEMA_signal_11063, mcs1_mcs_mat1_5_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_11068, new_AGEMA_signal_11067, new_AGEMA_signal_11066, mcs1_mcs_mat1_5_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_12334, new_AGEMA_signal_12333, new_AGEMA_signal_12332, mcs1_mcs_mat1_5_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_15229, new_AGEMA_signal_15228, new_AGEMA_signal_15227, mcs1_mcs_mat1_5_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_9829, new_AGEMA_signal_9828, new_AGEMA_signal_9827, mcs1_mcs_mat1_5_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_16318, new_AGEMA_signal_16317, new_AGEMA_signal_16316, mcs1_mcs_mat1_5_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_13777, new_AGEMA_signal_13776, new_AGEMA_signal_13775, mcs1_mcs_mat1_5_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .c ({new_AGEMA_signal_15229, new_AGEMA_signal_15228, new_AGEMA_signal_15227, mcs1_mcs_mat1_5_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_8968, new_AGEMA_signal_8967, new_AGEMA_signal_8966, mcs1_mcs_mat1_5_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_12337, new_AGEMA_signal_12336, new_AGEMA_signal_12335, mcs1_mcs_mat1_5_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_13777, new_AGEMA_signal_13776, new_AGEMA_signal_13775, mcs1_mcs_mat1_5_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5339], Fresh[5338], Fresh[5337], Fresh[5336], Fresh[5335], Fresh[5334]}), .c ({new_AGEMA_signal_12337, new_AGEMA_signal_12336, new_AGEMA_signal_12335, mcs1_mcs_mat1_5_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5345], Fresh[5344], Fresh[5343], Fresh[5342], Fresh[5341], Fresh[5340]}), .c ({new_AGEMA_signal_9829, new_AGEMA_signal_9828, new_AGEMA_signal_9827, mcs1_mcs_mat1_5_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5351], Fresh[5350], Fresh[5349], Fresh[5348], Fresh[5347], Fresh[5346]}), .c ({new_AGEMA_signal_11068, new_AGEMA_signal_11067, new_AGEMA_signal_11066, mcs1_mcs_mat1_5_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_17830, new_AGEMA_signal_17829, new_AGEMA_signal_17828, mcs1_mcs_mat1_5_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_17833, new_AGEMA_signal_17832, new_AGEMA_signal_17831, mcs1_mcs_mat1_5_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_18490, new_AGEMA_signal_18489, new_AGEMA_signal_18488, mcs1_mcs_mat1_5_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_17824, new_AGEMA_signal_17823, new_AGEMA_signal_17822, mcs1_mcs_mat1_5_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_13783, new_AGEMA_signal_13782, new_AGEMA_signal_13781, mcs1_mcs_mat1_5_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_18493, new_AGEMA_signal_18492, new_AGEMA_signal_18491, mcs1_mcs_mat1_5_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_17158, new_AGEMA_signal_17157, new_AGEMA_signal_17156, mcs1_mcs_mat1_5_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_17824, new_AGEMA_signal_17823, new_AGEMA_signal_17822, mcs1_mcs_mat1_5_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_17827, new_AGEMA_signal_17826, new_AGEMA_signal_17825, mcs1_mcs_mat1_5_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_18496, new_AGEMA_signal_18495, new_AGEMA_signal_18494, mcs1_mcs_mat1_5_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_15232, new_AGEMA_signal_15231, new_AGEMA_signal_15230, mcs1_mcs_mat1_5_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_17158, new_AGEMA_signal_17157, new_AGEMA_signal_17156, mcs1_mcs_mat1_5_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_17827, new_AGEMA_signal_17826, new_AGEMA_signal_17825, mcs1_mcs_mat1_5_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_18499, new_AGEMA_signal_18498, new_AGEMA_signal_18497, mcs1_mcs_mat1_5_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .c ({new_AGEMA_signal_19162, new_AGEMA_signal_19161, new_AGEMA_signal_19160, mcs1_mcs_mat1_5_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_17830, new_AGEMA_signal_17829, new_AGEMA_signal_17828, mcs1_mcs_mat1_5_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_15232, new_AGEMA_signal_15231, new_AGEMA_signal_15230, mcs1_mcs_mat1_5_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_18499, new_AGEMA_signal_18498, new_AGEMA_signal_18497, mcs1_mcs_mat1_5_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5357], Fresh[5356], Fresh[5355], Fresh[5354], Fresh[5353], Fresh[5352]}), .c ({new_AGEMA_signal_17833, new_AGEMA_signal_17832, new_AGEMA_signal_17831, mcs1_mcs_mat1_5_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5363], Fresh[5362], Fresh[5361], Fresh[5360], Fresh[5359], Fresh[5358]}), .c ({new_AGEMA_signal_15232, new_AGEMA_signal_15231, new_AGEMA_signal_15230, mcs1_mcs_mat1_5_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5369], Fresh[5368], Fresh[5367], Fresh[5366], Fresh[5365], Fresh[5364]}), .c ({new_AGEMA_signal_17158, new_AGEMA_signal_17157, new_AGEMA_signal_17156, mcs1_mcs_mat1_5_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_13786, new_AGEMA_signal_13785, new_AGEMA_signal_13784, mcs1_mcs_mat1_5_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_15235, new_AGEMA_signal_15234, new_AGEMA_signal_15233, mcs1_mcs_mat1_5_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_11077, new_AGEMA_signal_11076, new_AGEMA_signal_11075, mcs1_mcs_mat1_5_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_12343, new_AGEMA_signal_12342, new_AGEMA_signal_12341, mcs1_mcs_mat1_5_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_15238, new_AGEMA_signal_15237, new_AGEMA_signal_15236, mcs1_mcs_mat1_5_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_9835, new_AGEMA_signal_9834, new_AGEMA_signal_9833, mcs1_mcs_mat1_5_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_16321, new_AGEMA_signal_16320, new_AGEMA_signal_16319, mcs1_mcs_mat1_5_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_13786, new_AGEMA_signal_13785, new_AGEMA_signal_13784, mcs1_mcs_mat1_5_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .c ({new_AGEMA_signal_15238, new_AGEMA_signal_15237, new_AGEMA_signal_15236, mcs1_mcs_mat1_5_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_8971, new_AGEMA_signal_8970, new_AGEMA_signal_8969, mcs1_mcs_mat1_5_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_12346, new_AGEMA_signal_12345, new_AGEMA_signal_12344, mcs1_mcs_mat1_5_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_13786, new_AGEMA_signal_13785, new_AGEMA_signal_13784, mcs1_mcs_mat1_5_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5375], Fresh[5374], Fresh[5373], Fresh[5372], Fresh[5371], Fresh[5370]}), .c ({new_AGEMA_signal_12346, new_AGEMA_signal_12345, new_AGEMA_signal_12344, mcs1_mcs_mat1_5_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5381], Fresh[5380], Fresh[5379], Fresh[5378], Fresh[5377], Fresh[5376]}), .c ({new_AGEMA_signal_9835, new_AGEMA_signal_9834, new_AGEMA_signal_9833, mcs1_mcs_mat1_5_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5387], Fresh[5386], Fresh[5385], Fresh[5384], Fresh[5383], Fresh[5382]}), .c ({new_AGEMA_signal_11077, new_AGEMA_signal_11076, new_AGEMA_signal_11075, mcs1_mcs_mat1_5_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_15241, new_AGEMA_signal_15240, new_AGEMA_signal_15239, mcs1_mcs_mat1_5_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_16324, new_AGEMA_signal_16323, new_AGEMA_signal_16322, mcs1_mcs_mat1_5_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_13792, new_AGEMA_signal_13791, new_AGEMA_signal_13790, mcs1_mcs_mat1_5_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_12352, new_AGEMA_signal_12351, new_AGEMA_signal_12350, mcs1_mcs_mat1_5_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_15241, new_AGEMA_signal_15240, new_AGEMA_signal_15239, mcs1_mcs_mat1_5_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({new_AGEMA_signal_10333, new_AGEMA_signal_10332, new_AGEMA_signal_10331, mcs1_mcs_mat1_5_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_12349, new_AGEMA_signal_12348, new_AGEMA_signal_12347, mcs1_mcs_mat1_5_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_12352, new_AGEMA_signal_12351, new_AGEMA_signal_12350, mcs1_mcs_mat1_5_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_10333, new_AGEMA_signal_10332, new_AGEMA_signal_10331, mcs1_mcs_mat1_5_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_13789, new_AGEMA_signal_13788, new_AGEMA_signal_13787, mcs1_mcs_mat1_5_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_9838, new_AGEMA_signal_9837, new_AGEMA_signal_9836, mcs1_mcs_mat1_5_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_9841, new_AGEMA_signal_9840, new_AGEMA_signal_9839, mcs1_mcs_mat1_5_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_10333, new_AGEMA_signal_10332, new_AGEMA_signal_10331, mcs1_mcs_mat1_5_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_11080, new_AGEMA_signal_11079, new_AGEMA_signal_11078, mcs1_mcs_mat1_5_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .c ({new_AGEMA_signal_12352, new_AGEMA_signal_12351, new_AGEMA_signal_12350, mcs1_mcs_mat1_5_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_15244, new_AGEMA_signal_15243, new_AGEMA_signal_15242, mcs1_mcs_mat1_5_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_9838, new_AGEMA_signal_9837, new_AGEMA_signal_9836, mcs1_mcs_mat1_5_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_16327, new_AGEMA_signal_16326, new_AGEMA_signal_16325, mcs1_mcs_mat1_5_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_13792, new_AGEMA_signal_13791, new_AGEMA_signal_13790, mcs1_mcs_mat1_5_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_11080, new_AGEMA_signal_11079, new_AGEMA_signal_11078, mcs1_mcs_mat1_5_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_15244, new_AGEMA_signal_15243, new_AGEMA_signal_15242, mcs1_mcs_mat1_5_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .b ({new_AGEMA_signal_12355, new_AGEMA_signal_12354, new_AGEMA_signal_12353, mcs1_mcs_mat1_5_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_13792, new_AGEMA_signal_13791, new_AGEMA_signal_13790, mcs1_mcs_mat1_5_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5393], Fresh[5392], Fresh[5391], Fresh[5390], Fresh[5389], Fresh[5388]}), .c ({new_AGEMA_signal_12355, new_AGEMA_signal_12354, new_AGEMA_signal_12353, mcs1_mcs_mat1_5_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5399], Fresh[5398], Fresh[5397], Fresh[5396], Fresh[5395], Fresh[5394]}), .c ({new_AGEMA_signal_9841, new_AGEMA_signal_9840, new_AGEMA_signal_9839, mcs1_mcs_mat1_5_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5405], Fresh[5404], Fresh[5403], Fresh[5402], Fresh[5401], Fresh[5400]}), .c ({new_AGEMA_signal_11080, new_AGEMA_signal_11079, new_AGEMA_signal_11078, mcs1_mcs_mat1_5_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_13795, new_AGEMA_signal_13794, new_AGEMA_signal_13793, mcs1_mcs_mat1_5_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_11083, new_AGEMA_signal_11082, new_AGEMA_signal_11081, mcs1_mcs_mat1_5_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_15247, new_AGEMA_signal_15246, new_AGEMA_signal_15245, mcs1_mcs_mat1_5_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_12361, new_AGEMA_signal_12360, new_AGEMA_signal_12359, mcs1_mcs_mat1_5_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_15250, new_AGEMA_signal_15249, new_AGEMA_signal_15248, mcs1_mcs_mat1_5_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_16330, new_AGEMA_signal_16329, new_AGEMA_signal_16328, mcs1_mcs_mat1_5_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_13795, new_AGEMA_signal_13794, new_AGEMA_signal_13793, mcs1_mcs_mat1_5_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_15250, new_AGEMA_signal_15249, new_AGEMA_signal_15248, mcs1_mcs_mat1_5_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_16333, new_AGEMA_signal_16332, new_AGEMA_signal_16331, mcs1_mcs_mat1_5_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_11083, new_AGEMA_signal_11082, new_AGEMA_signal_11081, mcs1_mcs_mat1_5_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_13798, new_AGEMA_signal_13797, new_AGEMA_signal_13796, mcs1_mcs_mat1_5_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_15250, new_AGEMA_signal_15249, new_AGEMA_signal_15248, mcs1_mcs_mat1_5_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({new_AGEMA_signal_9844, new_AGEMA_signal_9843, new_AGEMA_signal_9842, mcs1_mcs_mat1_5_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_11083, new_AGEMA_signal_11082, new_AGEMA_signal_11081, mcs1_mcs_mat1_5_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_12358, new_AGEMA_signal_12357, new_AGEMA_signal_12356, mcs1_mcs_mat1_5_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .c ({new_AGEMA_signal_13795, new_AGEMA_signal_13794, new_AGEMA_signal_13793, mcs1_mcs_mat1_5_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_11086, new_AGEMA_signal_11085, new_AGEMA_signal_11084, mcs1_mcs_mat1_5_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8977, new_AGEMA_signal_8976, new_AGEMA_signal_8975, mcs1_mcs_mat1_5_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_12358, new_AGEMA_signal_12357, new_AGEMA_signal_12356, mcs1_mcs_mat1_5_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_13798, new_AGEMA_signal_13797, new_AGEMA_signal_13796, mcs1_mcs_mat1_5_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_12361, new_AGEMA_signal_12360, new_AGEMA_signal_12359, mcs1_mcs_mat1_5_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_15253, new_AGEMA_signal_15252, new_AGEMA_signal_15251, mcs1_mcs_mat1_5_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_11086, new_AGEMA_signal_11085, new_AGEMA_signal_11084, mcs1_mcs_mat1_5_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_12361, new_AGEMA_signal_12360, new_AGEMA_signal_12359, mcs1_mcs_mat1_5_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({new_AGEMA_signal_12364, new_AGEMA_signal_12363, new_AGEMA_signal_12362, mcs1_mcs_mat1_5_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_13798, new_AGEMA_signal_13797, new_AGEMA_signal_13796, mcs1_mcs_mat1_5_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5411], Fresh[5410], Fresh[5409], Fresh[5408], Fresh[5407], Fresh[5406]}), .c ({new_AGEMA_signal_12364, new_AGEMA_signal_12363, new_AGEMA_signal_12362, mcs1_mcs_mat1_5_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5417], Fresh[5416], Fresh[5415], Fresh[5414], Fresh[5413], Fresh[5412]}), .c ({new_AGEMA_signal_9844, new_AGEMA_signal_9843, new_AGEMA_signal_9842, mcs1_mcs_mat1_5_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5423], Fresh[5422], Fresh[5421], Fresh[5420], Fresh[5419], Fresh[5418]}), .c ({new_AGEMA_signal_11086, new_AGEMA_signal_11085, new_AGEMA_signal_11084, mcs1_mcs_mat1_5_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_19168, new_AGEMA_signal_19167, new_AGEMA_signal_19166, mcs1_mcs_mat1_5_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .c ({new_AGEMA_signal_19885, new_AGEMA_signal_19884, new_AGEMA_signal_19883, mcs1_mcs_mat1_5_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({new_AGEMA_signal_18502, new_AGEMA_signal_18501, new_AGEMA_signal_18500, mcs1_mcs_mat1_5_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_19165, new_AGEMA_signal_19164, new_AGEMA_signal_19163, mcs1_mcs_mat1_5_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_19888, new_AGEMA_signal_19887, new_AGEMA_signal_19886, mcs1_mcs_mat1_5_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_17161, new_AGEMA_signal_17160, new_AGEMA_signal_17159, mcs1_mcs_mat1_5_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_20662, new_AGEMA_signal_20661, new_AGEMA_signal_20660, mcs1_mcs_mat1_5_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_19168, new_AGEMA_signal_19167, new_AGEMA_signal_19166, mcs1_mcs_mat1_5_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .c ({new_AGEMA_signal_19888, new_AGEMA_signal_19887, new_AGEMA_signal_19886, mcs1_mcs_mat1_5_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_15256, new_AGEMA_signal_15255, new_AGEMA_signal_15254, mcs1_mcs_mat1_5_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_18502, new_AGEMA_signal_18501, new_AGEMA_signal_18500, mcs1_mcs_mat1_5_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_19168, new_AGEMA_signal_19167, new_AGEMA_signal_19166, mcs1_mcs_mat1_5_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_13801, new_AGEMA_signal_13800, new_AGEMA_signal_13799, mcs1_mcs_mat1_5_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_17839, new_AGEMA_signal_17838, new_AGEMA_signal_17837, mcs1_mcs_mat1_5_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_18502, new_AGEMA_signal_18501, new_AGEMA_signal_18500, mcs1_mcs_mat1_5_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5429], Fresh[5428], Fresh[5427], Fresh[5426], Fresh[5425], Fresh[5424]}), .c ({new_AGEMA_signal_17839, new_AGEMA_signal_17838, new_AGEMA_signal_17837, mcs1_mcs_mat1_5_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5435], Fresh[5434], Fresh[5433], Fresh[5432], Fresh[5431], Fresh[5430]}), .c ({new_AGEMA_signal_15256, new_AGEMA_signal_15255, new_AGEMA_signal_15254, mcs1_mcs_mat1_5_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5441], Fresh[5440], Fresh[5439], Fresh[5438], Fresh[5437], Fresh[5436]}), .c ({new_AGEMA_signal_17161, new_AGEMA_signal_17160, new_AGEMA_signal_17159, mcs1_mcs_mat1_5_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_13810, new_AGEMA_signal_13809, new_AGEMA_signal_13808, mcs1_mcs_mat1_5_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_11089, new_AGEMA_signal_11088, new_AGEMA_signal_11087, mcs1_mcs_mat1_5_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_15259, new_AGEMA_signal_15258, new_AGEMA_signal_15257, mcs1_mcs_mat1_5_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_9847, new_AGEMA_signal_9846, new_AGEMA_signal_9845, mcs1_mcs_mat1_5_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_12367, new_AGEMA_signal_12366, new_AGEMA_signal_12365, mcs1_mcs_mat1_5_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_13804, new_AGEMA_signal_13803, new_AGEMA_signal_13802, mcs1_mcs_mat1_5_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({new_AGEMA_signal_12370, new_AGEMA_signal_12369, new_AGEMA_signal_12368, mcs1_mcs_mat1_5_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_13807, new_AGEMA_signal_13806, new_AGEMA_signal_13805, mcs1_mcs_mat1_5_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5447], Fresh[5446], Fresh[5445], Fresh[5444], Fresh[5443], Fresh[5442]}), .c ({new_AGEMA_signal_12370, new_AGEMA_signal_12369, new_AGEMA_signal_12368, mcs1_mcs_mat1_5_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5453], Fresh[5452], Fresh[5451], Fresh[5450], Fresh[5449], Fresh[5448]}), .c ({new_AGEMA_signal_9847, new_AGEMA_signal_9846, new_AGEMA_signal_9845, mcs1_mcs_mat1_5_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5459], Fresh[5458], Fresh[5457], Fresh[5456], Fresh[5455], Fresh[5454]}), .c ({new_AGEMA_signal_11089, new_AGEMA_signal_11088, new_AGEMA_signal_11087, mcs1_mcs_mat1_5_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_9853, new_AGEMA_signal_9852, new_AGEMA_signal_9851, mcs1_mcs_mat1_5_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_11092, new_AGEMA_signal_11091, new_AGEMA_signal_11090, mcs1_mcs_mat1_5_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_12373, new_AGEMA_signal_12372, new_AGEMA_signal_12371, mcs1_mcs_mat1_5_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_9856, new_AGEMA_signal_9855, new_AGEMA_signal_9854, mcs1_mcs_mat1_5_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_12376, new_AGEMA_signal_12375, new_AGEMA_signal_12374, mcs1_mcs_mat1_5_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_13816, new_AGEMA_signal_13815, new_AGEMA_signal_13814, mcs1_mcs_mat1_5_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_13819, new_AGEMA_signal_13818, new_AGEMA_signal_13817, mcs1_mcs_mat1_5_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_12379, new_AGEMA_signal_12378, new_AGEMA_signal_12377, mcs1_mcs_mat1_5_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_15265, new_AGEMA_signal_15264, new_AGEMA_signal_15263, mcs1_mcs_mat1_5_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_12382, new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_5_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_13819, new_AGEMA_signal_13818, new_AGEMA_signal_13817, mcs1_mcs_mat1_5_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5465], Fresh[5464], Fresh[5463], Fresh[5462], Fresh[5461], Fresh[5460]}), .c ({new_AGEMA_signal_12382, new_AGEMA_signal_12381, new_AGEMA_signal_12380, mcs1_mcs_mat1_5_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5471], Fresh[5470], Fresh[5469], Fresh[5468], Fresh[5467], Fresh[5466]}), .c ({new_AGEMA_signal_9856, new_AGEMA_signal_9855, new_AGEMA_signal_9854, mcs1_mcs_mat1_5_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5477], Fresh[5476], Fresh[5475], Fresh[5474], Fresh[5473], Fresh[5472]}), .c ({new_AGEMA_signal_11092, new_AGEMA_signal_11091, new_AGEMA_signal_11090, mcs1_mcs_mat1_5_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_12388, new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_5_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_13822, new_AGEMA_signal_13821, new_AGEMA_signal_13820, mcs1_mcs_mat1_5_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_15268, new_AGEMA_signal_15267, new_AGEMA_signal_15266, mcs1_mcs_mat1_5_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_15271, new_AGEMA_signal_15270, new_AGEMA_signal_15269, mcs1_mcs_mat1_5_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, new_AGEMA_signal_12383, mcs1_mcs_mat1_5_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_16339, new_AGEMA_signal_16338, new_AGEMA_signal_16337, mcs1_mcs_mat1_5_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_11095, new_AGEMA_signal_11094, new_AGEMA_signal_11093, mcs1_mcs_mat1_5_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_12385, new_AGEMA_signal_12384, new_AGEMA_signal_12383, mcs1_mcs_mat1_5_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({new_AGEMA_signal_15271, new_AGEMA_signal_15270, new_AGEMA_signal_15269, mcs1_mcs_mat1_5_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_16342, new_AGEMA_signal_16341, new_AGEMA_signal_16340, mcs1_mcs_mat1_5_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_8986, new_AGEMA_signal_8985, new_AGEMA_signal_8984, mcs1_mcs_mat1_5_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_13822, new_AGEMA_signal_13821, new_AGEMA_signal_13820, mcs1_mcs_mat1_5_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_15271, new_AGEMA_signal_15270, new_AGEMA_signal_15269, mcs1_mcs_mat1_5_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_9859, new_AGEMA_signal_9858, new_AGEMA_signal_9857, mcs1_mcs_mat1_5_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_12394, new_AGEMA_signal_12393, new_AGEMA_signal_12392, mcs1_mcs_mat1_5_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_13822, new_AGEMA_signal_13821, new_AGEMA_signal_13820, mcs1_mcs_mat1_5_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_12391, new_AGEMA_signal_12390, new_AGEMA_signal_12389, mcs1_mcs_mat1_5_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_13825, new_AGEMA_signal_13824, new_AGEMA_signal_13823, mcs1_mcs_mat1_5_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_15274, new_AGEMA_signal_15273, new_AGEMA_signal_15272, mcs1_mcs_mat1_5_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_12388, new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_5_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_9859, new_AGEMA_signal_9858, new_AGEMA_signal_9857, mcs1_mcs_mat1_5_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_13825, new_AGEMA_signal_13824, new_AGEMA_signal_13823, mcs1_mcs_mat1_5_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_11095, new_AGEMA_signal_11094, new_AGEMA_signal_11093, mcs1_mcs_mat1_5_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_12388, new_AGEMA_signal_12387, new_AGEMA_signal_12386, mcs1_mcs_mat1_5_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5483], Fresh[5482], Fresh[5481], Fresh[5480], Fresh[5479], Fresh[5478]}), .c ({new_AGEMA_signal_12394, new_AGEMA_signal_12393, new_AGEMA_signal_12392, mcs1_mcs_mat1_5_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5489], Fresh[5488], Fresh[5487], Fresh[5486], Fresh[5485], Fresh[5484]}), .c ({new_AGEMA_signal_9859, new_AGEMA_signal_9858, new_AGEMA_signal_9857, mcs1_mcs_mat1_5_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5495], Fresh[5494], Fresh[5493], Fresh[5492], Fresh[5491], Fresh[5490]}), .c ({new_AGEMA_signal_11095, new_AGEMA_signal_11094, new_AGEMA_signal_11093, mcs1_mcs_mat1_5_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_11101, new_AGEMA_signal_11100, new_AGEMA_signal_11099, mcs1_mcs_mat1_5_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_12397, new_AGEMA_signal_12396, new_AGEMA_signal_12395, mcs1_mcs_mat1_5_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_16345, new_AGEMA_signal_16344, new_AGEMA_signal_16343, mcs1_mcs_mat1_5_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_9862, new_AGEMA_signal_9861, new_AGEMA_signal_9860, mcs1_mcs_mat1_5_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_17164, new_AGEMA_signal_17163, new_AGEMA_signal_17162, mcs1_mcs_mat1_5_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_15277, new_AGEMA_signal_15276, new_AGEMA_signal_15275, mcs1_mcs_mat1_5_mcs_out[47]}), .b ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .c ({new_AGEMA_signal_16345, new_AGEMA_signal_16344, new_AGEMA_signal_16343, mcs1_mcs_mat1_5_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_13828, new_AGEMA_signal_13827, new_AGEMA_signal_13826, mcs1_mcs_mat1_5_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .c ({new_AGEMA_signal_15277, new_AGEMA_signal_15276, new_AGEMA_signal_15275, mcs1_mcs_mat1_5_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_8989, new_AGEMA_signal_8988, new_AGEMA_signal_8987, mcs1_mcs_mat1_5_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_12400, new_AGEMA_signal_12399, new_AGEMA_signal_12398, mcs1_mcs_mat1_5_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_13828, new_AGEMA_signal_13827, new_AGEMA_signal_13826, mcs1_mcs_mat1_5_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5501], Fresh[5500], Fresh[5499], Fresh[5498], Fresh[5497], Fresh[5496]}), .c ({new_AGEMA_signal_12400, new_AGEMA_signal_12399, new_AGEMA_signal_12398, mcs1_mcs_mat1_5_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5507], Fresh[5506], Fresh[5505], Fresh[5504], Fresh[5503], Fresh[5502]}), .c ({new_AGEMA_signal_9862, new_AGEMA_signal_9861, new_AGEMA_signal_9860, mcs1_mcs_mat1_5_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5513], Fresh[5512], Fresh[5511], Fresh[5510], Fresh[5509], Fresh[5508]}), .c ({new_AGEMA_signal_11101, new_AGEMA_signal_11100, new_AGEMA_signal_11099, mcs1_mcs_mat1_5_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_13831, new_AGEMA_signal_13830, new_AGEMA_signal_13829, mcs1_mcs_mat1_5_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_11104, new_AGEMA_signal_11103, new_AGEMA_signal_11102, mcs1_mcs_mat1_5_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_15280, new_AGEMA_signal_15279, new_AGEMA_signal_15278, mcs1_mcs_mat1_5_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_12403, new_AGEMA_signal_12402, new_AGEMA_signal_12401, mcs1_mcs_mat1_5_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9865, new_AGEMA_signal_9864, new_AGEMA_signal_9863, mcs1_mcs_mat1_5_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_13831, new_AGEMA_signal_13830, new_AGEMA_signal_13829, mcs1_mcs_mat1_5_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_13834, new_AGEMA_signal_13833, new_AGEMA_signal_13832, mcs1_mcs_mat1_5_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_12409, new_AGEMA_signal_12408, new_AGEMA_signal_12407, mcs1_mcs_mat1_5_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_15283, new_AGEMA_signal_15282, new_AGEMA_signal_15281, mcs1_mcs_mat1_5_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_13837, new_AGEMA_signal_13836, new_AGEMA_signal_13835, mcs1_mcs_mat1_5_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_8992, new_AGEMA_signal_8991, new_AGEMA_signal_8990, mcs1_mcs_mat1_5_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_15286, new_AGEMA_signal_15285, new_AGEMA_signal_15284, mcs1_mcs_mat1_5_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_12403, new_AGEMA_signal_12402, new_AGEMA_signal_12401, mcs1_mcs_mat1_5_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_11107, new_AGEMA_signal_11106, new_AGEMA_signal_11105, mcs1_mcs_mat1_5_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_13837, new_AGEMA_signal_13836, new_AGEMA_signal_13835, mcs1_mcs_mat1_5_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_12406, new_AGEMA_signal_12405, new_AGEMA_signal_12404, mcs1_mcs_mat1_5_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_11107, new_AGEMA_signal_11106, new_AGEMA_signal_11105, mcs1_mcs_mat1_5_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_13840, new_AGEMA_signal_13839, new_AGEMA_signal_13838, mcs1_mcs_mat1_5_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5519], Fresh[5518], Fresh[5517], Fresh[5516], Fresh[5515], Fresh[5514]}), .c ({new_AGEMA_signal_12409, new_AGEMA_signal_12408, new_AGEMA_signal_12407, mcs1_mcs_mat1_5_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5525], Fresh[5524], Fresh[5523], Fresh[5522], Fresh[5521], Fresh[5520]}), .c ({new_AGEMA_signal_9865, new_AGEMA_signal_9864, new_AGEMA_signal_9863, mcs1_mcs_mat1_5_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5531], Fresh[5530], Fresh[5529], Fresh[5528], Fresh[5527], Fresh[5526]}), .c ({new_AGEMA_signal_11107, new_AGEMA_signal_11106, new_AGEMA_signal_11105, mcs1_mcs_mat1_5_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_15289, new_AGEMA_signal_15288, new_AGEMA_signal_15287, mcs1_mcs_mat1_5_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_8995, new_AGEMA_signal_8994, new_AGEMA_signal_8993, mcs1_mcs_mat1_5_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_16348, new_AGEMA_signal_16347, new_AGEMA_signal_16346, mcs1_mcs_mat1_5_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_11113, new_AGEMA_signal_11112, new_AGEMA_signal_11111, mcs1_mcs_mat1_5_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_11110, new_AGEMA_signal_11109, new_AGEMA_signal_11108, mcs1_mcs_mat1_5_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_12412, new_AGEMA_signal_12411, new_AGEMA_signal_12410, mcs1_mcs_mat1_5_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({new_AGEMA_signal_15289, new_AGEMA_signal_15288, new_AGEMA_signal_15287, mcs1_mcs_mat1_5_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_16351, new_AGEMA_signal_16350, new_AGEMA_signal_16349, mcs1_mcs_mat1_5_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_12415, new_AGEMA_signal_12414, new_AGEMA_signal_12413, mcs1_mcs_mat1_5_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_13843, new_AGEMA_signal_13842, new_AGEMA_signal_13841, mcs1_mcs_mat1_5_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_15289, new_AGEMA_signal_15288, new_AGEMA_signal_15287, mcs1_mcs_mat1_5_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_12418, new_AGEMA_signal_12417, new_AGEMA_signal_12416, mcs1_mcs_mat1_5_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_11116, new_AGEMA_signal_11115, new_AGEMA_signal_11114, mcs1_mcs_mat1_5_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_13843, new_AGEMA_signal_13842, new_AGEMA_signal_13841, mcs1_mcs_mat1_5_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_12418, new_AGEMA_signal_12417, new_AGEMA_signal_12416, mcs1_mcs_mat1_5_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_11113, new_AGEMA_signal_11112, new_AGEMA_signal_11111, mcs1_mcs_mat1_5_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_13846, new_AGEMA_signal_13845, new_AGEMA_signal_13844, mcs1_mcs_mat1_5_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .b ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, new_AGEMA_signal_10334, mcs1_mcs_mat1_5_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_11113, new_AGEMA_signal_11112, new_AGEMA_signal_11111, mcs1_mcs_mat1_5_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({new_AGEMA_signal_9868, new_AGEMA_signal_9867, new_AGEMA_signal_9866, mcs1_mcs_mat1_5_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_10336, new_AGEMA_signal_10335, new_AGEMA_signal_10334, mcs1_mcs_mat1_5_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5537], Fresh[5536], Fresh[5535], Fresh[5534], Fresh[5533], Fresh[5532]}), .c ({new_AGEMA_signal_12418, new_AGEMA_signal_12417, new_AGEMA_signal_12416, mcs1_mcs_mat1_5_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5543], Fresh[5542], Fresh[5541], Fresh[5540], Fresh[5539], Fresh[5538]}), .c ({new_AGEMA_signal_9868, new_AGEMA_signal_9867, new_AGEMA_signal_9866, mcs1_mcs_mat1_5_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5549], Fresh[5548], Fresh[5547], Fresh[5546], Fresh[5545], Fresh[5544]}), .c ({new_AGEMA_signal_11116, new_AGEMA_signal_11115, new_AGEMA_signal_11114, mcs1_mcs_mat1_5_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_17845, new_AGEMA_signal_17844, new_AGEMA_signal_17843, mcs1_mcs_mat1_5_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_17167, new_AGEMA_signal_17166, new_AGEMA_signal_17165, mcs1_mcs_mat1_5_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_18508, new_AGEMA_signal_18507, new_AGEMA_signal_18506, mcs1_mcs_mat1_5_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_15292, new_AGEMA_signal_15291, new_AGEMA_signal_15290, mcs1_mcs_mat1_5_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_16354, new_AGEMA_signal_16353, new_AGEMA_signal_16352, mcs1_mcs_mat1_5_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_19891, new_AGEMA_signal_19890, new_AGEMA_signal_19889, mcs1_mcs_mat1_5_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_17848, new_AGEMA_signal_17847, new_AGEMA_signal_17846, mcs1_mcs_mat1_5_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_20665, new_AGEMA_signal_20664, new_AGEMA_signal_20663, mcs1_mcs_mat1_5_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5555], Fresh[5554], Fresh[5553], Fresh[5552], Fresh[5551], Fresh[5550]}), .c ({new_AGEMA_signal_17848, new_AGEMA_signal_17847, new_AGEMA_signal_17846, mcs1_mcs_mat1_5_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5561], Fresh[5560], Fresh[5559], Fresh[5558], Fresh[5557], Fresh[5556]}), .c ({new_AGEMA_signal_15292, new_AGEMA_signal_15291, new_AGEMA_signal_15290, mcs1_mcs_mat1_5_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5567], Fresh[5566], Fresh[5565], Fresh[5564], Fresh[5563], Fresh[5562]}), .c ({new_AGEMA_signal_17167, new_AGEMA_signal_17166, new_AGEMA_signal_17165, mcs1_mcs_mat1_5_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_15295, new_AGEMA_signal_15294, new_AGEMA_signal_15293, mcs1_mcs_mat1_5_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_13852, new_AGEMA_signal_13851, new_AGEMA_signal_13850, mcs1_mcs_mat1_5_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_16357, new_AGEMA_signal_16356, new_AGEMA_signal_16355, mcs1_mcs_mat1_5_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_9874, new_AGEMA_signal_9873, new_AGEMA_signal_9872, mcs1_mcs_mat1_5_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_13855, new_AGEMA_signal_13854, new_AGEMA_signal_13853, mcs1_mcs_mat1_5_mcs_out[29]}), .c ({new_AGEMA_signal_15295, new_AGEMA_signal_15294, new_AGEMA_signal_15293, mcs1_mcs_mat1_5_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_9871, new_AGEMA_signal_9870, new_AGEMA_signal_9869, mcs1_mcs_mat1_5_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_13852, new_AGEMA_signal_13851, new_AGEMA_signal_13850, mcs1_mcs_mat1_5_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_15298, new_AGEMA_signal_15297, new_AGEMA_signal_15296, mcs1_mcs_mat1_5_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_12427, new_AGEMA_signal_12426, new_AGEMA_signal_12425, mcs1_mcs_mat1_5_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .c ({new_AGEMA_signal_13852, new_AGEMA_signal_13851, new_AGEMA_signal_13850, mcs1_mcs_mat1_5_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_15301, new_AGEMA_signal_15300, new_AGEMA_signal_15299, mcs1_mcs_mat1_5_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_12421, new_AGEMA_signal_12420, new_AGEMA_signal_12419, mcs1_mcs_mat1_5_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_16360, new_AGEMA_signal_16359, new_AGEMA_signal_16358, mcs1_mcs_mat1_5_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_13858, new_AGEMA_signal_13857, new_AGEMA_signal_13856, mcs1_mcs_mat1_5_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_12424, new_AGEMA_signal_12423, new_AGEMA_signal_12422, mcs1_mcs_mat1_5_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_15301, new_AGEMA_signal_15300, new_AGEMA_signal_15299, mcs1_mcs_mat1_5_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_11119, new_AGEMA_signal_11118, new_AGEMA_signal_11117, mcs1_mcs_mat1_5_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_12424, new_AGEMA_signal_12423, new_AGEMA_signal_12422, mcs1_mcs_mat1_5_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_12427, new_AGEMA_signal_12426, new_AGEMA_signal_12425, mcs1_mcs_mat1_5_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_9874, new_AGEMA_signal_9873, new_AGEMA_signal_9872, mcs1_mcs_mat1_5_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_13858, new_AGEMA_signal_13857, new_AGEMA_signal_13856, mcs1_mcs_mat1_5_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5573], Fresh[5572], Fresh[5571], Fresh[5570], Fresh[5569], Fresh[5568]}), .c ({new_AGEMA_signal_12427, new_AGEMA_signal_12426, new_AGEMA_signal_12425, mcs1_mcs_mat1_5_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5579], Fresh[5578], Fresh[5577], Fresh[5576], Fresh[5575], Fresh[5574]}), .c ({new_AGEMA_signal_9874, new_AGEMA_signal_9873, new_AGEMA_signal_9872, mcs1_mcs_mat1_5_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5585], Fresh[5584], Fresh[5583], Fresh[5582], Fresh[5581], Fresh[5580]}), .c ({new_AGEMA_signal_11119, new_AGEMA_signal_11118, new_AGEMA_signal_11117, mcs1_mcs_mat1_5_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_12430, new_AGEMA_signal_12429, new_AGEMA_signal_12428, mcs1_mcs_mat1_5_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_13861, new_AGEMA_signal_13860, new_AGEMA_signal_13859, mcs1_mcs_mat1_5_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_11122, new_AGEMA_signal_11121, new_AGEMA_signal_11120, mcs1_mcs_mat1_5_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_9877, new_AGEMA_signal_9876, new_AGEMA_signal_9875, mcs1_mcs_mat1_5_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_12430, new_AGEMA_signal_12429, new_AGEMA_signal_12428, mcs1_mcs_mat1_5_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_13864, new_AGEMA_signal_13863, new_AGEMA_signal_13862, mcs1_mcs_mat1_5_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_15304, new_AGEMA_signal_15303, new_AGEMA_signal_15302, mcs1_mcs_mat1_5_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_12436, new_AGEMA_signal_12435, new_AGEMA_signal_12434, mcs1_mcs_mat1_5_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_9877, new_AGEMA_signal_9876, new_AGEMA_signal_9875, mcs1_mcs_mat1_5_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_13864, new_AGEMA_signal_13863, new_AGEMA_signal_13862, mcs1_mcs_mat1_5_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_15307, new_AGEMA_signal_15306, new_AGEMA_signal_15305, mcs1_mcs_mat1_5_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .c ({new_AGEMA_signal_16363, new_AGEMA_signal_16362, new_AGEMA_signal_16361, mcs1_mcs_mat1_5_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_12436, new_AGEMA_signal_12435, new_AGEMA_signal_12434, mcs1_mcs_mat1_5_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_13867, new_AGEMA_signal_13866, new_AGEMA_signal_13865, mcs1_mcs_mat1_5_mcs_out[24]}), .c ({new_AGEMA_signal_15307, new_AGEMA_signal_15306, new_AGEMA_signal_15305, mcs1_mcs_mat1_5_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_12433, new_AGEMA_signal_12432, new_AGEMA_signal_12431, mcs1_mcs_mat1_5_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .c ({new_AGEMA_signal_13867, new_AGEMA_signal_13866, new_AGEMA_signal_13865, mcs1_mcs_mat1_5_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_11122, new_AGEMA_signal_11121, new_AGEMA_signal_11120, mcs1_mcs_mat1_5_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_9001, new_AGEMA_signal_9000, new_AGEMA_signal_8999, mcs1_mcs_mat1_5_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_12433, new_AGEMA_signal_12432, new_AGEMA_signal_12431, mcs1_mcs_mat1_5_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5591], Fresh[5590], Fresh[5589], Fresh[5588], Fresh[5587], Fresh[5586]}), .c ({new_AGEMA_signal_12436, new_AGEMA_signal_12435, new_AGEMA_signal_12434, mcs1_mcs_mat1_5_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5597], Fresh[5596], Fresh[5595], Fresh[5594], Fresh[5593], Fresh[5592]}), .c ({new_AGEMA_signal_9877, new_AGEMA_signal_9876, new_AGEMA_signal_9875, mcs1_mcs_mat1_5_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5603], Fresh[5602], Fresh[5601], Fresh[5600], Fresh[5599], Fresh[5598]}), .c ({new_AGEMA_signal_11122, new_AGEMA_signal_11121, new_AGEMA_signal_11120, mcs1_mcs_mat1_5_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_12439, new_AGEMA_signal_12438, new_AGEMA_signal_12437, mcs1_mcs_mat1_5_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .c ({new_AGEMA_signal_13870, new_AGEMA_signal_13869, new_AGEMA_signal_13868, mcs1_mcs_mat1_5_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_11125, new_AGEMA_signal_11124, new_AGEMA_signal_11123, mcs1_mcs_mat1_5_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_9880, new_AGEMA_signal_9879, new_AGEMA_signal_9878, mcs1_mcs_mat1_5_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_12439, new_AGEMA_signal_12438, new_AGEMA_signal_12437, mcs1_mcs_mat1_5_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_13873, new_AGEMA_signal_13872, new_AGEMA_signal_13871, mcs1_mcs_mat1_5_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .c ({new_AGEMA_signal_15310, new_AGEMA_signal_15309, new_AGEMA_signal_15308, mcs1_mcs_mat1_5_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_12445, new_AGEMA_signal_12444, new_AGEMA_signal_12443, mcs1_mcs_mat1_5_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_9880, new_AGEMA_signal_9879, new_AGEMA_signal_9878, mcs1_mcs_mat1_5_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_13873, new_AGEMA_signal_13872, new_AGEMA_signal_13871, mcs1_mcs_mat1_5_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_15313, new_AGEMA_signal_15312, new_AGEMA_signal_15311, mcs1_mcs_mat1_5_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_8401, new_AGEMA_signal_8400, new_AGEMA_signal_8399, mcs1_mcs_mat1_5_mcs_out[86]}), .c ({new_AGEMA_signal_16366, new_AGEMA_signal_16365, new_AGEMA_signal_16364, mcs1_mcs_mat1_5_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_12445, new_AGEMA_signal_12444, new_AGEMA_signal_12443, mcs1_mcs_mat1_5_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_13876, new_AGEMA_signal_13875, new_AGEMA_signal_13874, mcs1_mcs_mat1_5_mcs_out[20]}), .c ({new_AGEMA_signal_15313, new_AGEMA_signal_15312, new_AGEMA_signal_15311, mcs1_mcs_mat1_5_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_12442, new_AGEMA_signal_12441, new_AGEMA_signal_12440, mcs1_mcs_mat1_5_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .c ({new_AGEMA_signal_13876, new_AGEMA_signal_13875, new_AGEMA_signal_13874, mcs1_mcs_mat1_5_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_11125, new_AGEMA_signal_11124, new_AGEMA_signal_11123, mcs1_mcs_mat1_5_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_9004, new_AGEMA_signal_9003, new_AGEMA_signal_9002, mcs1_mcs_mat1_5_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_12442, new_AGEMA_signal_12441, new_AGEMA_signal_12440, mcs1_mcs_mat1_5_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5609], Fresh[5608], Fresh[5607], Fresh[5606], Fresh[5605], Fresh[5604]}), .c ({new_AGEMA_signal_12445, new_AGEMA_signal_12444, new_AGEMA_signal_12443, mcs1_mcs_mat1_5_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5615], Fresh[5614], Fresh[5613], Fresh[5612], Fresh[5611], Fresh[5610]}), .c ({new_AGEMA_signal_9880, new_AGEMA_signal_9879, new_AGEMA_signal_9878, mcs1_mcs_mat1_5_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5621], Fresh[5620], Fresh[5619], Fresh[5618], Fresh[5617], Fresh[5616]}), .c ({new_AGEMA_signal_11125, new_AGEMA_signal_11124, new_AGEMA_signal_11123, mcs1_mcs_mat1_5_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_17851, new_AGEMA_signal_17850, new_AGEMA_signal_17849, mcs1_mcs_mat1_5_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_17860, new_AGEMA_signal_17859, new_AGEMA_signal_17858, mcs1_mcs_mat1_5_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_18514, new_AGEMA_signal_18513, new_AGEMA_signal_18512, mcs1_mcs_mat1_5_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_18517, new_AGEMA_signal_18516, new_AGEMA_signal_18515, mcs1_mcs_mat1_5_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_13879, new_AGEMA_signal_13878, new_AGEMA_signal_13877, mcs1_mcs_mat1_5_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_19174, new_AGEMA_signal_19173, new_AGEMA_signal_19172, mcs1_mcs_mat1_5_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_19177, new_AGEMA_signal_19176, new_AGEMA_signal_19175, mcs1_mcs_mat1_5_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_15316, new_AGEMA_signal_15315, new_AGEMA_signal_15314, mcs1_mcs_mat1_5_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_19894, new_AGEMA_signal_19893, new_AGEMA_signal_19892, mcs1_mcs_mat1_5_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_11398, new_AGEMA_signal_11397, new_AGEMA_signal_11396, mcs1_mcs_mat1_5_mcs_out[50]}), .b ({new_AGEMA_signal_18517, new_AGEMA_signal_18516, new_AGEMA_signal_18515, mcs1_mcs_mat1_5_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_19177, new_AGEMA_signal_19176, new_AGEMA_signal_19175, mcs1_mcs_mat1_5_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_17854, new_AGEMA_signal_17853, new_AGEMA_signal_17852, mcs1_mcs_mat1_5_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .c ({new_AGEMA_signal_18517, new_AGEMA_signal_18516, new_AGEMA_signal_18515, mcs1_mcs_mat1_5_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_17170, new_AGEMA_signal_17169, new_AGEMA_signal_17168, mcs1_mcs_mat1_5_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_17173, new_AGEMA_signal_17172, new_AGEMA_signal_17171, mcs1_mcs_mat1_5_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_17854, new_AGEMA_signal_17853, new_AGEMA_signal_17852, mcs1_mcs_mat1_5_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_17857, new_AGEMA_signal_17856, new_AGEMA_signal_17855, mcs1_mcs_mat1_5_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_15316, new_AGEMA_signal_15315, new_AGEMA_signal_15314, mcs1_mcs_mat1_5_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_18520, new_AGEMA_signal_18519, new_AGEMA_signal_18518, mcs1_mcs_mat1_5_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5627], Fresh[5626], Fresh[5625], Fresh[5624], Fresh[5623], Fresh[5622]}), .c ({new_AGEMA_signal_17860, new_AGEMA_signal_17859, new_AGEMA_signal_17858, mcs1_mcs_mat1_5_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5633], Fresh[5632], Fresh[5631], Fresh[5630], Fresh[5629], Fresh[5628]}), .c ({new_AGEMA_signal_15316, new_AGEMA_signal_15315, new_AGEMA_signal_15314, mcs1_mcs_mat1_5_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5639], Fresh[5638], Fresh[5637], Fresh[5636], Fresh[5635], Fresh[5634]}), .c ({new_AGEMA_signal_17173, new_AGEMA_signal_17172, new_AGEMA_signal_17171, mcs1_mcs_mat1_5_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_15325, new_AGEMA_signal_15324, new_AGEMA_signal_15323, mcs1_mcs_mat1_5_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_10339, new_AGEMA_signal_10338, new_AGEMA_signal_10337, mcs1_mcs_mat1_5_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_16369, new_AGEMA_signal_16368, new_AGEMA_signal_16367, mcs1_mcs_mat1_5_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_13888, new_AGEMA_signal_13887, new_AGEMA_signal_13886, mcs1_mcs_mat1_5_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_13882, new_AGEMA_signal_13881, new_AGEMA_signal_13880, mcs1_mcs_mat1_5_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_15319, new_AGEMA_signal_15318, new_AGEMA_signal_15317, mcs1_mcs_mat1_5_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_12451, new_AGEMA_signal_12450, new_AGEMA_signal_12449, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_9883, new_AGEMA_signal_9882, new_AGEMA_signal_9881, mcs1_mcs_mat1_5_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_13882, new_AGEMA_signal_13881, new_AGEMA_signal_13880, mcs1_mcs_mat1_5_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_10339, new_AGEMA_signal_10338, new_AGEMA_signal_10337, mcs1_mcs_mat1_5_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_13885, new_AGEMA_signal_13884, new_AGEMA_signal_13883, mcs1_mcs_mat1_5_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_15322, new_AGEMA_signal_15321, new_AGEMA_signal_15320, mcs1_mcs_mat1_5_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_12448, new_AGEMA_signal_12447, new_AGEMA_signal_12446, mcs1_mcs_mat1_5_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_12451, new_AGEMA_signal_12450, new_AGEMA_signal_12449, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_13885, new_AGEMA_signal_13884, new_AGEMA_signal_13883, mcs1_mcs_mat1_5_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_9007, new_AGEMA_signal_9006, new_AGEMA_signal_9005, mcs1_mcs_mat1_5_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_9883, new_AGEMA_signal_9882, new_AGEMA_signal_9881, mcs1_mcs_mat1_5_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_10339, new_AGEMA_signal_10338, new_AGEMA_signal_10337, mcs1_mcs_mat1_5_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_16372, new_AGEMA_signal_16371, new_AGEMA_signal_16370, mcs1_mcs_mat1_5_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .c ({new_AGEMA_signal_17176, new_AGEMA_signal_17175, new_AGEMA_signal_17174, mcs1_mcs_mat1_5_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_15325, new_AGEMA_signal_15324, new_AGEMA_signal_15323, mcs1_mcs_mat1_5_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_12451, new_AGEMA_signal_12450, new_AGEMA_signal_12449, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_16372, new_AGEMA_signal_16371, new_AGEMA_signal_16370, mcs1_mcs_mat1_5_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({new_AGEMA_signal_13888, new_AGEMA_signal_13887, new_AGEMA_signal_13886, mcs1_mcs_mat1_5_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_15325, new_AGEMA_signal_15324, new_AGEMA_signal_15323, mcs1_mcs_mat1_5_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({new_AGEMA_signal_12448, new_AGEMA_signal_12447, new_AGEMA_signal_12446, mcs1_mcs_mat1_5_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_13888, new_AGEMA_signal_13887, new_AGEMA_signal_13886, mcs1_mcs_mat1_5_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_8368, new_AGEMA_signal_8367, new_AGEMA_signal_8366, shiftr_out[104]}), .b ({new_AGEMA_signal_11128, new_AGEMA_signal_11127, new_AGEMA_signal_11126, mcs1_mcs_mat1_5_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_12448, new_AGEMA_signal_12447, new_AGEMA_signal_12446, mcs1_mcs_mat1_5_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10408, new_AGEMA_signal_10407, new_AGEMA_signal_10406, mcs1_mcs_mat1_5_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5645], Fresh[5644], Fresh[5643], Fresh[5642], Fresh[5641], Fresh[5640]}), .c ({new_AGEMA_signal_12451, new_AGEMA_signal_12450, new_AGEMA_signal_12449, mcs1_mcs_mat1_5_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8572, new_AGEMA_signal_8571, new_AGEMA_signal_8570, mcs1_mcs_mat1_5_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5651], Fresh[5650], Fresh[5649], Fresh[5648], Fresh[5647], Fresh[5646]}), .c ({new_AGEMA_signal_9883, new_AGEMA_signal_9882, new_AGEMA_signal_9881, mcs1_mcs_mat1_5_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10210, new_AGEMA_signal_10209, new_AGEMA_signal_10208, mcs1_mcs_mat1_5_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5657], Fresh[5656], Fresh[5655], Fresh[5654], Fresh[5653], Fresh[5652]}), .c ({new_AGEMA_signal_11128, new_AGEMA_signal_11127, new_AGEMA_signal_11126, mcs1_mcs_mat1_5_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, new_AGEMA_signal_10340, mcs1_mcs_mat1_5_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .c ({new_AGEMA_signal_11131, new_AGEMA_signal_11130, new_AGEMA_signal_11129, mcs1_mcs_mat1_5_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_13894, new_AGEMA_signal_13893, new_AGEMA_signal_13892, mcs1_mcs_mat1_5_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .c ({new_AGEMA_signal_15328, new_AGEMA_signal_15327, new_AGEMA_signal_15326, mcs1_mcs_mat1_5_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_12454, new_AGEMA_signal_12453, new_AGEMA_signal_12452, mcs1_mcs_mat1_5_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .c ({new_AGEMA_signal_13891, new_AGEMA_signal_13890, new_AGEMA_signal_13889, mcs1_mcs_mat1_5_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_11134, new_AGEMA_signal_11133, new_AGEMA_signal_11132, mcs1_mcs_mat1_5_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, new_AGEMA_signal_10340, mcs1_mcs_mat1_5_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_12454, new_AGEMA_signal_12453, new_AGEMA_signal_12452, mcs1_mcs_mat1_5_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_9010, new_AGEMA_signal_9009, new_AGEMA_signal_9008, mcs1_mcs_mat1_5_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_9886, new_AGEMA_signal_9885, new_AGEMA_signal_9884, mcs1_mcs_mat1_5_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_10342, new_AGEMA_signal_10341, new_AGEMA_signal_10340, mcs1_mcs_mat1_5_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_15331, new_AGEMA_signal_15330, new_AGEMA_signal_15329, mcs1_mcs_mat1_5_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_8383, new_AGEMA_signal_8382, new_AGEMA_signal_8381, shiftr_out[72]}), .c ({new_AGEMA_signal_16375, new_AGEMA_signal_16374, new_AGEMA_signal_16373, mcs1_mcs_mat1_5_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_9010, new_AGEMA_signal_9009, new_AGEMA_signal_9008, mcs1_mcs_mat1_5_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_13894, new_AGEMA_signal_13893, new_AGEMA_signal_13892, mcs1_mcs_mat1_5_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_15331, new_AGEMA_signal_15330, new_AGEMA_signal_15329, mcs1_mcs_mat1_5_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_12457, new_AGEMA_signal_12456, new_AGEMA_signal_12455, mcs1_mcs_mat1_5_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_11134, new_AGEMA_signal_11133, new_AGEMA_signal_11132, mcs1_mcs_mat1_5_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_13894, new_AGEMA_signal_13893, new_AGEMA_signal_13892, mcs1_mcs_mat1_5_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10423, new_AGEMA_signal_10422, new_AGEMA_signal_10421, mcs1_mcs_mat1_5_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5663], Fresh[5662], Fresh[5661], Fresh[5660], Fresh[5659], Fresh[5658]}), .c ({new_AGEMA_signal_12457, new_AGEMA_signal_12456, new_AGEMA_signal_12455, mcs1_mcs_mat1_5_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8587, new_AGEMA_signal_8586, new_AGEMA_signal_8585, mcs1_mcs_mat1_5_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5669], Fresh[5668], Fresh[5667], Fresh[5666], Fresh[5665], Fresh[5664]}), .c ({new_AGEMA_signal_9886, new_AGEMA_signal_9885, new_AGEMA_signal_9884, mcs1_mcs_mat1_5_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10224, new_AGEMA_signal_10223, shiftr_out[75]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5675], Fresh[5674], Fresh[5673], Fresh[5672], Fresh[5671], Fresh[5670]}), .c ({new_AGEMA_signal_11134, new_AGEMA_signal_11133, new_AGEMA_signal_11132, mcs1_mcs_mat1_5_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_17179, new_AGEMA_signal_17178, new_AGEMA_signal_17177, mcs1_mcs_mat1_5_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_11140, new_AGEMA_signal_11139, new_AGEMA_signal_11138, mcs1_mcs_mat1_5_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_17863, new_AGEMA_signal_17862, new_AGEMA_signal_17861, mcs1_mcs_mat1_5_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_16378, new_AGEMA_signal_16377, new_AGEMA_signal_16376, mcs1_mcs_mat1_5_mcs_out[7]}), .b ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .c ({new_AGEMA_signal_17179, new_AGEMA_signal_17178, new_AGEMA_signal_17177, mcs1_mcs_mat1_5_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_15334, new_AGEMA_signal_15333, new_AGEMA_signal_15332, mcs1_mcs_mat1_5_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .c ({new_AGEMA_signal_16378, new_AGEMA_signal_16377, new_AGEMA_signal_16376, mcs1_mcs_mat1_5_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_13897, new_AGEMA_signal_13896, new_AGEMA_signal_13895, mcs1_mcs_mat1_5_mcs_out[6]}), .b ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, new_AGEMA_signal_9890, mcs1_mcs_mat1_5_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_15334, new_AGEMA_signal_15333, new_AGEMA_signal_15332, mcs1_mcs_mat1_5_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_9889, new_AGEMA_signal_9888, new_AGEMA_signal_9887, mcs1_mcs_mat1_5_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_12460, new_AGEMA_signal_12459, new_AGEMA_signal_12458, mcs1_mcs_mat1_5_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_13897, new_AGEMA_signal_13896, new_AGEMA_signal_13895, mcs1_mcs_mat1_5_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10440, new_AGEMA_signal_10439, shiftr_out[41]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5681], Fresh[5680], Fresh[5679], Fresh[5678], Fresh[5677], Fresh[5676]}), .c ({new_AGEMA_signal_12460, new_AGEMA_signal_12459, new_AGEMA_signal_12458, mcs1_mcs_mat1_5_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8604, new_AGEMA_signal_8603, shiftr_out[42]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5687], Fresh[5686], Fresh[5685], Fresh[5684], Fresh[5683], Fresh[5682]}), .c ({new_AGEMA_signal_9892, new_AGEMA_signal_9891, new_AGEMA_signal_9890, mcs1_mcs_mat1_5_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10243, new_AGEMA_signal_10242, new_AGEMA_signal_10241, mcs1_mcs_mat1_5_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5693], Fresh[5692], Fresh[5691], Fresh[5690], Fresh[5689], Fresh[5688]}), .c ({new_AGEMA_signal_11140, new_AGEMA_signal_11139, new_AGEMA_signal_11138, mcs1_mcs_mat1_5_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_17182, new_AGEMA_signal_17181, new_AGEMA_signal_17180, mcs1_mcs_mat1_5_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_17866, new_AGEMA_signal_17865, new_AGEMA_signal_17864, mcs1_mcs_mat1_5_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_18526, new_AGEMA_signal_18525, new_AGEMA_signal_18524, mcs1_mcs_mat1_5_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .b ({new_AGEMA_signal_17185, new_AGEMA_signal_17184, new_AGEMA_signal_17183, mcs1_mcs_mat1_5_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_17866, new_AGEMA_signal_17865, new_AGEMA_signal_17864, mcs1_mcs_mat1_5_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_18529, new_AGEMA_signal_18528, new_AGEMA_signal_18527, mcs1_mcs_mat1_5_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_15337, new_AGEMA_signal_15336, new_AGEMA_signal_15335, mcs1_mcs_mat1_5_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_19180, new_AGEMA_signal_19179, new_AGEMA_signal_19178, mcs1_mcs_mat1_5_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_18532, new_AGEMA_signal_18531, new_AGEMA_signal_18530, mcs1_mcs_mat1_5_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_17872, new_AGEMA_signal_17871, new_AGEMA_signal_17870, mcs1_mcs_mat1_5_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_19183, new_AGEMA_signal_19182, new_AGEMA_signal_19181, mcs1_mcs_mat1_5_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_17875, new_AGEMA_signal_17874, new_AGEMA_signal_17873, mcs1_mcs_mat1_5_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_13900, new_AGEMA_signal_13899, new_AGEMA_signal_13898, mcs1_mcs_mat1_5_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_18532, new_AGEMA_signal_18531, new_AGEMA_signal_18530, mcs1_mcs_mat1_5_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16624, new_AGEMA_signal_16623, new_AGEMA_signal_16622, shiftr_out[9]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5699], Fresh[5698], Fresh[5697], Fresh[5696], Fresh[5695], Fresh[5694]}), .c ({new_AGEMA_signal_17875, new_AGEMA_signal_17874, new_AGEMA_signal_17873, mcs1_mcs_mat1_5_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12838, new_AGEMA_signal_12837, new_AGEMA_signal_12836, shiftr_out[10]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5705], Fresh[5704], Fresh[5703], Fresh[5702], Fresh[5701], Fresh[5700]}), .c ({new_AGEMA_signal_15337, new_AGEMA_signal_15336, new_AGEMA_signal_15335, mcs1_mcs_mat1_5_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_5_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15712, new_AGEMA_signal_15711, new_AGEMA_signal_15710, mcs1_mcs_mat1_5_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5711], Fresh[5710], Fresh[5709], Fresh[5708], Fresh[5707], Fresh[5706]}), .c ({new_AGEMA_signal_17185, new_AGEMA_signal_17184, new_AGEMA_signal_17183, mcs1_mcs_mat1_5_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U96 ( .a ({new_AGEMA_signal_20668, new_AGEMA_signal_20667, new_AGEMA_signal_20666, mcs1_mcs_mat1_6_n128}), .b ({new_AGEMA_signal_16381, new_AGEMA_signal_16380, new_AGEMA_signal_16379, mcs1_mcs_mat1_6_n127}), .c ({temp_next_s3[69], temp_next_s2[69], temp_next_s1[69], temp_next_s0[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U95 ( .a ({new_AGEMA_signal_15445, new_AGEMA_signal_15444, new_AGEMA_signal_15443, mcs1_mcs_mat1_6_mcs_out[41]}), .b ({new_AGEMA_signal_12556, new_AGEMA_signal_12555, new_AGEMA_signal_12554, mcs1_mcs_mat1_6_mcs_out[45]}), .c ({new_AGEMA_signal_16381, new_AGEMA_signal_16380, new_AGEMA_signal_16379, mcs1_mcs_mat1_6_n127}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U94 ( .a ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, new_AGEMA_signal_10346, mcs1_mcs_mat1_6_mcs_out[33]}), .b ({new_AGEMA_signal_19963, new_AGEMA_signal_19962, new_AGEMA_signal_19961, mcs1_mcs_mat1_6_mcs_out[37]}), .c ({new_AGEMA_signal_20668, new_AGEMA_signal_20667, new_AGEMA_signal_20666, mcs1_mcs_mat1_6_n128}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U93 ( .a ({new_AGEMA_signal_19186, new_AGEMA_signal_19185, new_AGEMA_signal_19184, mcs1_mcs_mat1_6_n126}), .b ({new_AGEMA_signal_17878, new_AGEMA_signal_17877, new_AGEMA_signal_17876, mcs1_mcs_mat1_6_n125}), .c ({temp_next_s3[68], temp_next_s2[68], temp_next_s1[68], temp_next_s0[68]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U92 ( .a ({new_AGEMA_signal_14014, new_AGEMA_signal_14013, new_AGEMA_signal_14012, mcs1_mcs_mat1_6_mcs_out[40]}), .b ({new_AGEMA_signal_17260, new_AGEMA_signal_17259, new_AGEMA_signal_17258, mcs1_mcs_mat1_6_mcs_out[44]}), .c ({new_AGEMA_signal_17878, new_AGEMA_signal_17877, new_AGEMA_signal_17876, mcs1_mcs_mat1_6_n125}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U91 ( .a ({new_AGEMA_signal_17272, new_AGEMA_signal_17271, new_AGEMA_signal_17270, mcs1_mcs_mat1_6_mcs_out[32]}), .b ({new_AGEMA_signal_18583, new_AGEMA_signal_18582, new_AGEMA_signal_18581, mcs1_mcs_mat1_6_mcs_out[36]}), .c ({new_AGEMA_signal_19186, new_AGEMA_signal_19185, new_AGEMA_signal_19184, mcs1_mcs_mat1_6_n126}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U90 ( .a ({new_AGEMA_signal_19189, new_AGEMA_signal_19188, new_AGEMA_signal_19187, mcs1_mcs_mat1_6_n124}), .b ({new_AGEMA_signal_17188, new_AGEMA_signal_17187, new_AGEMA_signal_17186, mcs1_mcs_mat1_6_n123}), .c ({temp_next_s3[39], temp_next_s2[39], temp_next_s1[39], temp_next_s0[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U89 ( .a ({new_AGEMA_signal_14035, new_AGEMA_signal_14034, new_AGEMA_signal_14033, mcs1_mcs_mat1_6_mcs_out[27]}), .b ({new_AGEMA_signal_16471, new_AGEMA_signal_16470, new_AGEMA_signal_16469, mcs1_mcs_mat1_6_mcs_out[31]}), .c ({new_AGEMA_signal_17188, new_AGEMA_signal_17187, new_AGEMA_signal_17186, mcs1_mcs_mat1_6_n123}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U88 ( .a ({new_AGEMA_signal_14047, new_AGEMA_signal_14046, new_AGEMA_signal_14045, mcs1_mcs_mat1_6_mcs_out[19]}), .b ({new_AGEMA_signal_18586, new_AGEMA_signal_18585, new_AGEMA_signal_18584, mcs1_mcs_mat1_6_mcs_out[23]}), .c ({new_AGEMA_signal_19189, new_AGEMA_signal_19188, new_AGEMA_signal_19187, mcs1_mcs_mat1_6_n124}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U87 ( .a ({new_AGEMA_signal_19903, new_AGEMA_signal_19902, new_AGEMA_signal_19901, mcs1_mcs_mat1_6_n122}), .b ({new_AGEMA_signal_16384, new_AGEMA_signal_16383, new_AGEMA_signal_16382, mcs1_mcs_mat1_6_n121}), .c ({temp_next_s3[38], temp_next_s2[38], temp_next_s1[38], temp_next_s0[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U86 ( .a ({new_AGEMA_signal_15463, new_AGEMA_signal_15462, new_AGEMA_signal_15461, mcs1_mcs_mat1_6_mcs_out[26]}), .b ({new_AGEMA_signal_15457, new_AGEMA_signal_15456, new_AGEMA_signal_15455, mcs1_mcs_mat1_6_mcs_out[30]}), .c ({new_AGEMA_signal_16384, new_AGEMA_signal_16383, new_AGEMA_signal_16382, mcs1_mcs_mat1_6_n121}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U85 ( .a ({new_AGEMA_signal_15472, new_AGEMA_signal_15471, new_AGEMA_signal_15470, mcs1_mcs_mat1_6_mcs_out[18]}), .b ({new_AGEMA_signal_19252, new_AGEMA_signal_19251, new_AGEMA_signal_19250, mcs1_mcs_mat1_6_mcs_out[22]}), .c ({new_AGEMA_signal_19903, new_AGEMA_signal_19902, new_AGEMA_signal_19901, mcs1_mcs_mat1_6_n122}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U84 ( .a ({new_AGEMA_signal_20674, new_AGEMA_signal_20673, new_AGEMA_signal_20672, mcs1_mcs_mat1_6_n120}), .b ({new_AGEMA_signal_17191, new_AGEMA_signal_17190, new_AGEMA_signal_17189, mcs1_mcs_mat1_6_n119}), .c ({temp_next_s3[37], temp_next_s2[37], temp_next_s1[37], temp_next_s0[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U83 ( .a ({new_AGEMA_signal_16477, new_AGEMA_signal_16476, new_AGEMA_signal_16475, mcs1_mcs_mat1_6_mcs_out[25]}), .b ({new_AGEMA_signal_14029, new_AGEMA_signal_14028, new_AGEMA_signal_14027, mcs1_mcs_mat1_6_mcs_out[29]}), .c ({new_AGEMA_signal_17191, new_AGEMA_signal_17190, new_AGEMA_signal_17189, mcs1_mcs_mat1_6_n119}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U82 ( .a ({new_AGEMA_signal_16480, new_AGEMA_signal_16479, new_AGEMA_signal_16478, mcs1_mcs_mat1_6_mcs_out[17]}), .b ({new_AGEMA_signal_19966, new_AGEMA_signal_19965, new_AGEMA_signal_19964, mcs1_mcs_mat1_6_mcs_out[21]}), .c ({new_AGEMA_signal_20674, new_AGEMA_signal_20673, new_AGEMA_signal_20672, mcs1_mcs_mat1_6_n120}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U81 ( .a ({new_AGEMA_signal_19192, new_AGEMA_signal_19191, new_AGEMA_signal_19190, mcs1_mcs_mat1_6_n118}), .b ({new_AGEMA_signal_17194, new_AGEMA_signal_17193, new_AGEMA_signal_17192, mcs1_mcs_mat1_6_n117}), .c ({temp_next_s3[36], temp_next_s2[36], temp_next_s1[36], temp_next_s0[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U80 ( .a ({new_AGEMA_signal_14041, new_AGEMA_signal_14040, new_AGEMA_signal_14039, mcs1_mcs_mat1_6_mcs_out[24]}), .b ({new_AGEMA_signal_16474, new_AGEMA_signal_16473, new_AGEMA_signal_16472, mcs1_mcs_mat1_6_mcs_out[28]}), .c ({new_AGEMA_signal_17194, new_AGEMA_signal_17193, new_AGEMA_signal_17192, mcs1_mcs_mat1_6_n117}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U79 ( .a ({new_AGEMA_signal_14053, new_AGEMA_signal_14052, new_AGEMA_signal_14051, mcs1_mcs_mat1_6_mcs_out[16]}), .b ({new_AGEMA_signal_18592, new_AGEMA_signal_18591, new_AGEMA_signal_18590, mcs1_mcs_mat1_6_mcs_out[20]}), .c ({new_AGEMA_signal_19192, new_AGEMA_signal_19191, new_AGEMA_signal_19190, mcs1_mcs_mat1_6_n118}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U78 ( .a ({new_AGEMA_signal_17197, new_AGEMA_signal_17196, new_AGEMA_signal_17195, mcs1_mcs_mat1_6_n116}), .b ({new_AGEMA_signal_20677, new_AGEMA_signal_20676, new_AGEMA_signal_20675, mcs1_mcs_mat1_6_n115}), .c ({temp_next_s3[7], temp_next_s2[7], temp_next_s1[7], temp_next_s0[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U77 ( .a ({new_AGEMA_signal_14074, new_AGEMA_signal_14073, new_AGEMA_signal_14072, mcs1_mcs_mat1_6_mcs_out[3]}), .b ({new_AGEMA_signal_19969, new_AGEMA_signal_19968, new_AGEMA_signal_19967, mcs1_mcs_mat1_6_mcs_out[7]}), .c ({new_AGEMA_signal_20677, new_AGEMA_signal_20676, new_AGEMA_signal_20675, mcs1_mcs_mat1_6_n115}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U76 ( .a ({new_AGEMA_signal_11236, new_AGEMA_signal_11235, new_AGEMA_signal_11234, mcs1_mcs_mat1_6_mcs_out[11]}), .b ({new_AGEMA_signal_16483, new_AGEMA_signal_16482, new_AGEMA_signal_16481, mcs1_mcs_mat1_6_mcs_out[15]}), .c ({new_AGEMA_signal_17197, new_AGEMA_signal_17196, new_AGEMA_signal_17195, mcs1_mcs_mat1_6_n116}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U75 ( .a ({new_AGEMA_signal_20680, new_AGEMA_signal_20679, new_AGEMA_signal_20678, mcs1_mcs_mat1_6_n114}), .b ({new_AGEMA_signal_17200, new_AGEMA_signal_17199, new_AGEMA_signal_17198, mcs1_mcs_mat1_6_n113}), .c ({new_AGEMA_signal_21307, new_AGEMA_signal_21306, new_AGEMA_signal_21305, mcs_out[231]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U74 ( .a ({new_AGEMA_signal_16414, new_AGEMA_signal_16413, new_AGEMA_signal_16412, mcs1_mcs_mat1_6_mcs_out[123]}), .b ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_17200, new_AGEMA_signal_17199, new_AGEMA_signal_17198, mcs1_mcs_mat1_6_n113}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U73 ( .a ({new_AGEMA_signal_15364, new_AGEMA_signal_15363, new_AGEMA_signal_15362, mcs1_mcs_mat1_6_mcs_out[115]}), .b ({new_AGEMA_signal_19942, new_AGEMA_signal_19941, new_AGEMA_signal_19940, mcs1_mcs_mat1_6_mcs_out[119]}), .c ({new_AGEMA_signal_20680, new_AGEMA_signal_20679, new_AGEMA_signal_20678, mcs1_mcs_mat1_6_n114}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U72 ( .a ({new_AGEMA_signal_20683, new_AGEMA_signal_20682, new_AGEMA_signal_20681, mcs1_mcs_mat1_6_n112}), .b ({new_AGEMA_signal_13903, new_AGEMA_signal_13902, new_AGEMA_signal_13901, mcs1_mcs_mat1_6_n111}), .c ({new_AGEMA_signal_21310, new_AGEMA_signal_21309, new_AGEMA_signal_21308, mcs_out[230]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U71 ( .a ({new_AGEMA_signal_12463, new_AGEMA_signal_12462, new_AGEMA_signal_12461, mcs1_mcs_mat1_6_mcs_out[122]}), .b ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_13903, new_AGEMA_signal_13902, new_AGEMA_signal_13901, mcs1_mcs_mat1_6_n111}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U70 ( .a ({new_AGEMA_signal_13921, new_AGEMA_signal_13920, new_AGEMA_signal_13919, mcs1_mcs_mat1_6_mcs_out[114]}), .b ({new_AGEMA_signal_19945, new_AGEMA_signal_19944, new_AGEMA_signal_19943, mcs1_mcs_mat1_6_mcs_out[118]}), .c ({new_AGEMA_signal_20683, new_AGEMA_signal_20682, new_AGEMA_signal_20681, mcs1_mcs_mat1_6_n112}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U69 ( .a ({new_AGEMA_signal_16387, new_AGEMA_signal_16386, new_AGEMA_signal_16385, mcs1_mcs_mat1_6_n110}), .b ({new_AGEMA_signal_19195, new_AGEMA_signal_19194, new_AGEMA_signal_19193, mcs1_mcs_mat1_6_n109}), .c ({temp_next_s3[6], temp_next_s2[6], temp_next_s1[6], temp_next_s0[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U68 ( .a ({new_AGEMA_signal_14077, new_AGEMA_signal_14076, new_AGEMA_signal_14075, mcs1_mcs_mat1_6_mcs_out[2]}), .b ({new_AGEMA_signal_18595, new_AGEMA_signal_18594, new_AGEMA_signal_18593, mcs1_mcs_mat1_6_mcs_out[6]}), .c ({new_AGEMA_signal_19195, new_AGEMA_signal_19194, new_AGEMA_signal_19193, mcs1_mcs_mat1_6_n109}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U67 ( .a ({new_AGEMA_signal_15487, new_AGEMA_signal_15486, new_AGEMA_signal_15485, mcs1_mcs_mat1_6_mcs_out[10]}), .b ({new_AGEMA_signal_15478, new_AGEMA_signal_15477, new_AGEMA_signal_15476, mcs1_mcs_mat1_6_mcs_out[14]}), .c ({new_AGEMA_signal_16387, new_AGEMA_signal_16386, new_AGEMA_signal_16385, mcs1_mcs_mat1_6_n110}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U66 ( .a ({new_AGEMA_signal_19912, new_AGEMA_signal_19911, new_AGEMA_signal_19910, mcs1_mcs_mat1_6_n108}), .b ({new_AGEMA_signal_17203, new_AGEMA_signal_17202, new_AGEMA_signal_17201, mcs1_mcs_mat1_6_n107}), .c ({new_AGEMA_signal_20686, new_AGEMA_signal_20685, new_AGEMA_signal_20684, mcs_out[229]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U65 ( .a ({new_AGEMA_signal_16417, new_AGEMA_signal_16416, new_AGEMA_signal_16415, mcs1_mcs_mat1_6_mcs_out[121]}), .b ({new_AGEMA_signal_11143, new_AGEMA_signal_11142, new_AGEMA_signal_11141, mcs1_mcs_mat1_6_mcs_out[125]}), .c ({new_AGEMA_signal_17203, new_AGEMA_signal_17202, new_AGEMA_signal_17201, mcs1_mcs_mat1_6_n107}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U64 ( .a ({new_AGEMA_signal_12469, new_AGEMA_signal_12468, new_AGEMA_signal_12467, mcs1_mcs_mat1_6_mcs_out[113]}), .b ({new_AGEMA_signal_19222, new_AGEMA_signal_19221, new_AGEMA_signal_19220, mcs1_mcs_mat1_6_mcs_out[117]}), .c ({new_AGEMA_signal_19912, new_AGEMA_signal_19911, new_AGEMA_signal_19910, mcs1_mcs_mat1_6_n108}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U63 ( .a ({new_AGEMA_signal_19198, new_AGEMA_signal_19197, new_AGEMA_signal_19196, mcs1_mcs_mat1_6_n106}), .b ({new_AGEMA_signal_16390, new_AGEMA_signal_16389, new_AGEMA_signal_16388, mcs1_mcs_mat1_6_n105}), .c ({new_AGEMA_signal_19915, new_AGEMA_signal_19914, new_AGEMA_signal_19913, mcs_out[228]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U62 ( .a ({new_AGEMA_signal_15358, new_AGEMA_signal_15357, new_AGEMA_signal_15356, mcs1_mcs_mat1_6_mcs_out[120]}), .b ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_16390, new_AGEMA_signal_16389, new_AGEMA_signal_16388, mcs1_mcs_mat1_6_n105}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U61 ( .a ({new_AGEMA_signal_16420, new_AGEMA_signal_16419, new_AGEMA_signal_16418, mcs1_mcs_mat1_6_mcs_out[112]}), .b ({new_AGEMA_signal_18553, new_AGEMA_signal_18552, new_AGEMA_signal_18551, mcs1_mcs_mat1_6_mcs_out[116]}), .c ({new_AGEMA_signal_19198, new_AGEMA_signal_19197, new_AGEMA_signal_19196, mcs1_mcs_mat1_6_n106}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U60 ( .a ({new_AGEMA_signal_19918, new_AGEMA_signal_19917, new_AGEMA_signal_19916, mcs1_mcs_mat1_6_n104}), .b ({new_AGEMA_signal_17206, new_AGEMA_signal_17205, new_AGEMA_signal_17204, mcs1_mcs_mat1_6_n103}), .c ({new_AGEMA_signal_20689, new_AGEMA_signal_20688, new_AGEMA_signal_20687, mcs_out[199]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U59 ( .a ({new_AGEMA_signal_16423, new_AGEMA_signal_16422, new_AGEMA_signal_16421, mcs1_mcs_mat1_6_mcs_out[111]}), .b ({new_AGEMA_signal_16438, new_AGEMA_signal_16437, new_AGEMA_signal_16436, mcs1_mcs_mat1_6_mcs_out[99]}), .c ({new_AGEMA_signal_17206, new_AGEMA_signal_17205, new_AGEMA_signal_17204, mcs1_mcs_mat1_6_n103}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U58 ( .a ({new_AGEMA_signal_19225, new_AGEMA_signal_19224, new_AGEMA_signal_19223, mcs1_mcs_mat1_6_mcs_out[103]}), .b ({new_AGEMA_signal_15376, new_AGEMA_signal_15375, new_AGEMA_signal_15374, mcs1_mcs_mat1_6_mcs_out[107]}), .c ({new_AGEMA_signal_19918, new_AGEMA_signal_19917, new_AGEMA_signal_19916, mcs1_mcs_mat1_6_n104}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U57 ( .a ({new_AGEMA_signal_18535, new_AGEMA_signal_18534, new_AGEMA_signal_18533, mcs1_mcs_mat1_6_n102}), .b ({new_AGEMA_signal_17209, new_AGEMA_signal_17208, new_AGEMA_signal_17207, mcs1_mcs_mat1_6_n101}), .c ({new_AGEMA_signal_19201, new_AGEMA_signal_19200, new_AGEMA_signal_19199, mcs_out[198]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U56 ( .a ({new_AGEMA_signal_16426, new_AGEMA_signal_16425, new_AGEMA_signal_16424, mcs1_mcs_mat1_6_mcs_out[110]}), .b ({new_AGEMA_signal_13945, new_AGEMA_signal_13944, new_AGEMA_signal_13943, mcs1_mcs_mat1_6_mcs_out[98]}), .c ({new_AGEMA_signal_17209, new_AGEMA_signal_17208, new_AGEMA_signal_17207, mcs1_mcs_mat1_6_n101}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U55 ( .a ({new_AGEMA_signal_17899, new_AGEMA_signal_17898, new_AGEMA_signal_17897, mcs1_mcs_mat1_6_mcs_out[102]}), .b ({new_AGEMA_signal_15379, new_AGEMA_signal_15378, new_AGEMA_signal_15377, mcs1_mcs_mat1_6_mcs_out[106]}), .c ({new_AGEMA_signal_18535, new_AGEMA_signal_18534, new_AGEMA_signal_18533, mcs1_mcs_mat1_6_n102}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U54 ( .a ({new_AGEMA_signal_19204, new_AGEMA_signal_19203, new_AGEMA_signal_19202, mcs1_mcs_mat1_6_n100}), .b ({new_AGEMA_signal_17212, new_AGEMA_signal_17211, new_AGEMA_signal_17210, mcs1_mcs_mat1_6_n99}), .c ({new_AGEMA_signal_19921, new_AGEMA_signal_19920, new_AGEMA_signal_19919, mcs_out[197]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U53 ( .a ({new_AGEMA_signal_16429, new_AGEMA_signal_16428, new_AGEMA_signal_16427, mcs1_mcs_mat1_6_mcs_out[109]}), .b ({new_AGEMA_signal_11167, new_AGEMA_signal_11166, new_AGEMA_signal_11165, mcs1_mcs_mat1_6_mcs_out[97]}), .c ({new_AGEMA_signal_17212, new_AGEMA_signal_17211, new_AGEMA_signal_17210, mcs1_mcs_mat1_6_n99}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U52 ( .a ({new_AGEMA_signal_18559, new_AGEMA_signal_18558, new_AGEMA_signal_18557, mcs1_mcs_mat1_6_mcs_out[101]}), .b ({new_AGEMA_signal_15382, new_AGEMA_signal_15381, new_AGEMA_signal_15380, mcs1_mcs_mat1_6_mcs_out[105]}), .c ({new_AGEMA_signal_19204, new_AGEMA_signal_19203, new_AGEMA_signal_19202, mcs1_mcs_mat1_6_n100}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U51 ( .a ({new_AGEMA_signal_19924, new_AGEMA_signal_19923, new_AGEMA_signal_19922, mcs1_mcs_mat1_6_n98}), .b ({new_AGEMA_signal_18538, new_AGEMA_signal_18537, new_AGEMA_signal_18536, mcs1_mcs_mat1_6_n97}), .c ({new_AGEMA_signal_20692, new_AGEMA_signal_20691, new_AGEMA_signal_20690, mcs_out[196]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U50 ( .a ({new_AGEMA_signal_16432, new_AGEMA_signal_16431, new_AGEMA_signal_16430, mcs1_mcs_mat1_6_mcs_out[108]}), .b ({new_AGEMA_signal_17911, new_AGEMA_signal_17910, new_AGEMA_signal_17909, mcs1_mcs_mat1_6_mcs_out[96]}), .c ({new_AGEMA_signal_18538, new_AGEMA_signal_18537, new_AGEMA_signal_18536, mcs1_mcs_mat1_6_n97}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U49 ( .a ({new_AGEMA_signal_19228, new_AGEMA_signal_19227, new_AGEMA_signal_19226, mcs1_mcs_mat1_6_mcs_out[100]}), .b ({new_AGEMA_signal_16435, new_AGEMA_signal_16434, new_AGEMA_signal_16433, mcs1_mcs_mat1_6_mcs_out[104]}), .c ({new_AGEMA_signal_19924, new_AGEMA_signal_19923, new_AGEMA_signal_19922, mcs1_mcs_mat1_6_n98}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U48 ( .a ({new_AGEMA_signal_18541, new_AGEMA_signal_18540, new_AGEMA_signal_18539, mcs1_mcs_mat1_6_n96}), .b ({new_AGEMA_signal_16393, new_AGEMA_signal_16392, new_AGEMA_signal_16391, mcs1_mcs_mat1_6_n95}), .c ({new_AGEMA_signal_19207, new_AGEMA_signal_19206, new_AGEMA_signal_19205, mcs_out[167]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U47 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_15394, new_AGEMA_signal_15393, new_AGEMA_signal_15392, mcs1_mcs_mat1_6_mcs_out[95]}), .c ({new_AGEMA_signal_16393, new_AGEMA_signal_16392, new_AGEMA_signal_16391, mcs1_mcs_mat1_6_n95}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U46 ( .a ({new_AGEMA_signal_13951, new_AGEMA_signal_13950, new_AGEMA_signal_13949, mcs1_mcs_mat1_6_mcs_out[83]}), .b ({new_AGEMA_signal_17914, new_AGEMA_signal_17913, new_AGEMA_signal_17912, mcs1_mcs_mat1_6_mcs_out[87]}), .c ({new_AGEMA_signal_18541, new_AGEMA_signal_18540, new_AGEMA_signal_18539, mcs1_mcs_mat1_6_n96}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U45 ( .a ({new_AGEMA_signal_15340, new_AGEMA_signal_15339, new_AGEMA_signal_15338, mcs1_mcs_mat1_6_n94}), .b ({new_AGEMA_signal_13906, new_AGEMA_signal_13905, new_AGEMA_signal_13904, mcs1_mcs_mat1_6_n93}), .c ({new_AGEMA_signal_16396, new_AGEMA_signal_16395, new_AGEMA_signal_16394, mcs_out[166]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U43 ( .a ({new_AGEMA_signal_13954, new_AGEMA_signal_13953, new_AGEMA_signal_13952, mcs1_mcs_mat1_6_mcs_out[82]}), .b ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_15340, new_AGEMA_signal_15339, new_AGEMA_signal_15338, mcs1_mcs_mat1_6_n94}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U42 ( .a ({new_AGEMA_signal_17215, new_AGEMA_signal_17214, new_AGEMA_signal_17213, mcs1_mcs_mat1_6_n92}), .b ({new_AGEMA_signal_13909, new_AGEMA_signal_13908, new_AGEMA_signal_13907, mcs1_mcs_mat1_6_n91}), .c ({new_AGEMA_signal_17881, new_AGEMA_signal_17880, new_AGEMA_signal_17879, mcs_out[165]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U41 ( .a ({new_AGEMA_signal_11185, new_AGEMA_signal_11184, new_AGEMA_signal_11183, mcs1_mcs_mat1_6_mcs_out[89]}), .b ({new_AGEMA_signal_12496, new_AGEMA_signal_12495, new_AGEMA_signal_12494, mcs1_mcs_mat1_6_mcs_out[93]}), .c ({new_AGEMA_signal_13909, new_AGEMA_signal_13908, new_AGEMA_signal_13907, mcs1_mcs_mat1_6_n91}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U40 ( .a ({new_AGEMA_signal_13957, new_AGEMA_signal_13956, new_AGEMA_signal_13955, mcs1_mcs_mat1_6_mcs_out[81]}), .b ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_17215, new_AGEMA_signal_17214, new_AGEMA_signal_17213, mcs1_mcs_mat1_6_n92}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U39 ( .a ({new_AGEMA_signal_19210, new_AGEMA_signal_19209, new_AGEMA_signal_19208, mcs1_mcs_mat1_6_n90}), .b ({new_AGEMA_signal_17218, new_AGEMA_signal_17217, new_AGEMA_signal_17216, mcs1_mcs_mat1_6_n89}), .c ({new_AGEMA_signal_19927, new_AGEMA_signal_19926, new_AGEMA_signal_19925, mcs_out[164]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U38 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_16441, new_AGEMA_signal_16440, new_AGEMA_signal_16439, mcs1_mcs_mat1_6_mcs_out[92]}), .c ({new_AGEMA_signal_17218, new_AGEMA_signal_17217, new_AGEMA_signal_17216, mcs1_mcs_mat1_6_n89}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U37 ( .a ({new_AGEMA_signal_15400, new_AGEMA_signal_15399, new_AGEMA_signal_15398, mcs1_mcs_mat1_6_mcs_out[80]}), .b ({new_AGEMA_signal_18565, new_AGEMA_signal_18564, new_AGEMA_signal_18563, mcs1_mcs_mat1_6_mcs_out[84]}), .c ({new_AGEMA_signal_19210, new_AGEMA_signal_19209, new_AGEMA_signal_19208, mcs1_mcs_mat1_6_n90}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U36 ( .a ({new_AGEMA_signal_16399, new_AGEMA_signal_16398, new_AGEMA_signal_16397, mcs1_mcs_mat1_6_n88}), .b ({new_AGEMA_signal_17884, new_AGEMA_signal_17883, new_AGEMA_signal_17882, mcs1_mcs_mat1_6_n87}), .c ({temp_next_s3[5], temp_next_s2[5], temp_next_s1[5], temp_next_s0[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U35 ( .a ({new_AGEMA_signal_17281, new_AGEMA_signal_17280, new_AGEMA_signal_17279, mcs1_mcs_mat1_6_mcs_out[5]}), .b ({new_AGEMA_signal_14065, new_AGEMA_signal_14064, new_AGEMA_signal_14063, mcs1_mcs_mat1_6_mcs_out[9]}), .c ({new_AGEMA_signal_17884, new_AGEMA_signal_17883, new_AGEMA_signal_17882, mcs1_mcs_mat1_6_n87}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U34 ( .a ({new_AGEMA_signal_15481, new_AGEMA_signal_15480, new_AGEMA_signal_15479, mcs1_mcs_mat1_6_mcs_out[13]}), .b ({new_AGEMA_signal_15499, new_AGEMA_signal_15498, new_AGEMA_signal_15497, mcs1_mcs_mat1_6_mcs_out[1]}), .c ({new_AGEMA_signal_16399, new_AGEMA_signal_16398, new_AGEMA_signal_16397, mcs1_mcs_mat1_6_n88}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U33 ( .a ({new_AGEMA_signal_19930, new_AGEMA_signal_19929, new_AGEMA_signal_19928, mcs1_mcs_mat1_6_n86}), .b ({new_AGEMA_signal_16402, new_AGEMA_signal_16401, new_AGEMA_signal_16400, mcs1_mcs_mat1_6_n85}), .c ({new_AGEMA_signal_20695, new_AGEMA_signal_20694, new_AGEMA_signal_20693, mcs_out[135]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U32 ( .a ({new_AGEMA_signal_12520, new_AGEMA_signal_12519, new_AGEMA_signal_12518, mcs1_mcs_mat1_6_mcs_out[75]}), .b ({new_AGEMA_signal_15403, new_AGEMA_signal_15402, new_AGEMA_signal_15401, mcs1_mcs_mat1_6_mcs_out[79]}), .c ({new_AGEMA_signal_16402, new_AGEMA_signal_16401, new_AGEMA_signal_16400, mcs1_mcs_mat1_6_n85}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U31 ( .a ({new_AGEMA_signal_16453, new_AGEMA_signal_16452, new_AGEMA_signal_16451, mcs1_mcs_mat1_6_mcs_out[67]}), .b ({new_AGEMA_signal_19231, new_AGEMA_signal_19230, new_AGEMA_signal_19229, mcs1_mcs_mat1_6_mcs_out[71]}), .c ({new_AGEMA_signal_19930, new_AGEMA_signal_19929, new_AGEMA_signal_19928, mcs1_mcs_mat1_6_n86}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U30 ( .a ({new_AGEMA_signal_20698, new_AGEMA_signal_20697, new_AGEMA_signal_20696, mcs1_mcs_mat1_6_n84}), .b ({new_AGEMA_signal_17221, new_AGEMA_signal_17220, new_AGEMA_signal_17219, mcs1_mcs_mat1_6_n83}), .c ({new_AGEMA_signal_21313, new_AGEMA_signal_21312, new_AGEMA_signal_21311, mcs_out[134]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U29 ( .a ({new_AGEMA_signal_16447, new_AGEMA_signal_16446, new_AGEMA_signal_16445, mcs1_mcs_mat1_6_mcs_out[74]}), .b ({new_AGEMA_signal_9925, new_AGEMA_signal_9924, new_AGEMA_signal_9923, mcs1_mcs_mat1_6_mcs_out[78]}), .c ({new_AGEMA_signal_17221, new_AGEMA_signal_17220, new_AGEMA_signal_17219, mcs1_mcs_mat1_6_n83}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U28 ( .a ({new_AGEMA_signal_15418, new_AGEMA_signal_15417, new_AGEMA_signal_15416, mcs1_mcs_mat1_6_mcs_out[66]}), .b ({new_AGEMA_signal_19948, new_AGEMA_signal_19947, new_AGEMA_signal_19946, mcs1_mcs_mat1_6_mcs_out[70]}), .c ({new_AGEMA_signal_20698, new_AGEMA_signal_20697, new_AGEMA_signal_20696, mcs1_mcs_mat1_6_n84}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U27 ( .a ({new_AGEMA_signal_20701, new_AGEMA_signal_20700, new_AGEMA_signal_20699, mcs1_mcs_mat1_6_n82}), .b ({new_AGEMA_signal_15343, new_AGEMA_signal_15342, new_AGEMA_signal_15341, mcs1_mcs_mat1_6_n81}), .c ({new_AGEMA_signal_21316, new_AGEMA_signal_21315, new_AGEMA_signal_21314, mcs_out[133]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U26 ( .a ({new_AGEMA_signal_13966, new_AGEMA_signal_13965, new_AGEMA_signal_13964, mcs1_mcs_mat1_6_mcs_out[73]}), .b ({new_AGEMA_signal_12514, new_AGEMA_signal_12513, new_AGEMA_signal_12512, mcs1_mcs_mat1_6_mcs_out[77]}), .c ({new_AGEMA_signal_15343, new_AGEMA_signal_15342, new_AGEMA_signal_15341, mcs1_mcs_mat1_6_n81}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U25 ( .a ({new_AGEMA_signal_12529, new_AGEMA_signal_12528, new_AGEMA_signal_12527, mcs1_mcs_mat1_6_mcs_out[65]}), .b ({new_AGEMA_signal_19951, new_AGEMA_signal_19950, new_AGEMA_signal_19949, mcs1_mcs_mat1_6_mcs_out[69]}), .c ({new_AGEMA_signal_20701, new_AGEMA_signal_20700, new_AGEMA_signal_20699, mcs1_mcs_mat1_6_n82}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U24 ( .a ({new_AGEMA_signal_19933, new_AGEMA_signal_19932, new_AGEMA_signal_19931, mcs1_mcs_mat1_6_n80}), .b ({new_AGEMA_signal_17224, new_AGEMA_signal_17223, new_AGEMA_signal_17222, mcs1_mcs_mat1_6_n79}), .c ({new_AGEMA_signal_20704, new_AGEMA_signal_20703, new_AGEMA_signal_20702, mcs_out[132]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U23 ( .a ({new_AGEMA_signal_16450, new_AGEMA_signal_16449, new_AGEMA_signal_16448, mcs1_mcs_mat1_6_mcs_out[72]}), .b ({new_AGEMA_signal_16444, new_AGEMA_signal_16443, new_AGEMA_signal_16442, mcs1_mcs_mat1_6_mcs_out[76]}), .c ({new_AGEMA_signal_17224, new_AGEMA_signal_17223, new_AGEMA_signal_17222, mcs1_mcs_mat1_6_n79}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U22 ( .a ({new_AGEMA_signal_17254, new_AGEMA_signal_17253, new_AGEMA_signal_17252, mcs1_mcs_mat1_6_mcs_out[64]}), .b ({new_AGEMA_signal_19237, new_AGEMA_signal_19236, new_AGEMA_signal_19235, mcs1_mcs_mat1_6_mcs_out[68]}), .c ({new_AGEMA_signal_19933, new_AGEMA_signal_19932, new_AGEMA_signal_19931, mcs1_mcs_mat1_6_n80}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U21 ( .a ({new_AGEMA_signal_19936, new_AGEMA_signal_19935, new_AGEMA_signal_19934, mcs1_mcs_mat1_6_n78}), .b ({new_AGEMA_signal_16405, new_AGEMA_signal_16404, new_AGEMA_signal_16403, mcs1_mcs_mat1_6_n77}), .c ({temp_next_s3[103], temp_next_s2[103], temp_next_s1[103], temp_next_s0[103]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U20 ( .a ({new_AGEMA_signal_13987, new_AGEMA_signal_13986, new_AGEMA_signal_13985, mcs1_mcs_mat1_6_mcs_out[59]}), .b ({new_AGEMA_signal_15424, new_AGEMA_signal_15423, new_AGEMA_signal_15422, mcs1_mcs_mat1_6_mcs_out[63]}), .c ({new_AGEMA_signal_16405, new_AGEMA_signal_16404, new_AGEMA_signal_16403, mcs1_mcs_mat1_6_n77}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U19 ( .a ({new_AGEMA_signal_12553, new_AGEMA_signal_12552, new_AGEMA_signal_12551, mcs1_mcs_mat1_6_mcs_out[51]}), .b ({new_AGEMA_signal_19240, new_AGEMA_signal_19239, new_AGEMA_signal_19238, mcs1_mcs_mat1_6_mcs_out[55]}), .c ({new_AGEMA_signal_19936, new_AGEMA_signal_19935, new_AGEMA_signal_19934, mcs1_mcs_mat1_6_n78}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U18 ( .a ({new_AGEMA_signal_20710, new_AGEMA_signal_20709, new_AGEMA_signal_20708, mcs1_mcs_mat1_6_n76}), .b ({new_AGEMA_signal_15346, new_AGEMA_signal_15345, new_AGEMA_signal_15344, mcs1_mcs_mat1_6_n75}), .c ({temp_next_s3[102], temp_next_s2[102], temp_next_s1[102], temp_next_s0[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U17 ( .a ({new_AGEMA_signal_12541, new_AGEMA_signal_12540, new_AGEMA_signal_12539, mcs1_mcs_mat1_6_mcs_out[58]}), .b ({new_AGEMA_signal_13978, new_AGEMA_signal_13977, new_AGEMA_signal_13976, mcs1_mcs_mat1_6_mcs_out[62]}), .c ({new_AGEMA_signal_15346, new_AGEMA_signal_15345, new_AGEMA_signal_15344, mcs1_mcs_mat1_6_n75}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U16 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_19954, new_AGEMA_signal_19953, new_AGEMA_signal_19952, mcs1_mcs_mat1_6_mcs_out[54]}), .c ({new_AGEMA_signal_20710, new_AGEMA_signal_20709, new_AGEMA_signal_20708, mcs1_mcs_mat1_6_n76}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U15 ( .a ({new_AGEMA_signal_20713, new_AGEMA_signal_20712, new_AGEMA_signal_20711, mcs1_mcs_mat1_6_n74}), .b ({new_AGEMA_signal_15349, new_AGEMA_signal_15348, new_AGEMA_signal_15347, mcs1_mcs_mat1_6_n73}), .c ({temp_next_s3[101], temp_next_s2[101], temp_next_s1[101], temp_next_s0[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U14 ( .a ({new_AGEMA_signal_13990, new_AGEMA_signal_13989, new_AGEMA_signal_13988, mcs1_mcs_mat1_6_mcs_out[57]}), .b ({new_AGEMA_signal_13981, new_AGEMA_signal_13980, new_AGEMA_signal_13979, mcs1_mcs_mat1_6_mcs_out[61]}), .c ({new_AGEMA_signal_15349, new_AGEMA_signal_15348, new_AGEMA_signal_15347, mcs1_mcs_mat1_6_n73}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U13 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({new_AGEMA_signal_19957, new_AGEMA_signal_19956, new_AGEMA_signal_19955, mcs1_mcs_mat1_6_mcs_out[53]}), .c ({new_AGEMA_signal_20713, new_AGEMA_signal_20712, new_AGEMA_signal_20711, mcs1_mcs_mat1_6_n74}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U12 ( .a ({new_AGEMA_signal_19939, new_AGEMA_signal_19938, new_AGEMA_signal_19937, mcs1_mcs_mat1_6_n72}), .b ({new_AGEMA_signal_17227, new_AGEMA_signal_17226, new_AGEMA_signal_17225, mcs1_mcs_mat1_6_n71}), .c ({temp_next_s3[100], temp_next_s2[100], temp_next_s1[100], temp_next_s0[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U11 ( .a ({new_AGEMA_signal_15430, new_AGEMA_signal_15429, new_AGEMA_signal_15428, mcs1_mcs_mat1_6_mcs_out[56]}), .b ({new_AGEMA_signal_16459, new_AGEMA_signal_16458, new_AGEMA_signal_16457, mcs1_mcs_mat1_6_mcs_out[60]}), .c ({new_AGEMA_signal_17227, new_AGEMA_signal_17226, new_AGEMA_signal_17225, mcs1_mcs_mat1_6_n71}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U10 ( .a ({new_AGEMA_signal_13999, new_AGEMA_signal_13998, new_AGEMA_signal_13997, mcs1_mcs_mat1_6_mcs_out[48]}), .b ({new_AGEMA_signal_19246, new_AGEMA_signal_19245, new_AGEMA_signal_19244, mcs1_mcs_mat1_6_mcs_out[52]}), .c ({new_AGEMA_signal_19939, new_AGEMA_signal_19938, new_AGEMA_signal_19937, mcs1_mcs_mat1_6_n72}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U9 ( .a ({new_AGEMA_signal_20719, new_AGEMA_signal_20718, new_AGEMA_signal_20717, mcs1_mcs_mat1_6_n70}), .b ({new_AGEMA_signal_16408, new_AGEMA_signal_16407, new_AGEMA_signal_16406, mcs1_mcs_mat1_6_n69}), .c ({temp_next_s3[71], temp_next_s2[71], temp_next_s1[71], temp_next_s0[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U8 ( .a ({new_AGEMA_signal_15439, new_AGEMA_signal_15438, new_AGEMA_signal_15437, mcs1_mcs_mat1_6_mcs_out[43]}), .b ({new_AGEMA_signal_15436, new_AGEMA_signal_15435, new_AGEMA_signal_15434, mcs1_mcs_mat1_6_mcs_out[47]}), .c ({new_AGEMA_signal_16408, new_AGEMA_signal_16407, new_AGEMA_signal_16406, mcs1_mcs_mat1_6_n69}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U7 ( .a ({new_AGEMA_signal_15451, new_AGEMA_signal_15450, new_AGEMA_signal_15449, mcs1_mcs_mat1_6_mcs_out[35]}), .b ({new_AGEMA_signal_19960, new_AGEMA_signal_19959, new_AGEMA_signal_19958, mcs1_mcs_mat1_6_mcs_out[39]}), .c ({new_AGEMA_signal_20719, new_AGEMA_signal_20718, new_AGEMA_signal_20717, mcs1_mcs_mat1_6_n70}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U6 ( .a ({new_AGEMA_signal_18547, new_AGEMA_signal_18546, new_AGEMA_signal_18545, mcs1_mcs_mat1_6_n68}), .b ({new_AGEMA_signal_16411, new_AGEMA_signal_16410, new_AGEMA_signal_16409, mcs1_mcs_mat1_6_n67}), .c ({temp_next_s3[70], temp_next_s2[70], temp_next_s1[70], temp_next_s0[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U5 ( .a ({new_AGEMA_signal_15442, new_AGEMA_signal_15441, new_AGEMA_signal_15440, mcs1_mcs_mat1_6_mcs_out[42]}), .b ({new_AGEMA_signal_11206, new_AGEMA_signal_11205, new_AGEMA_signal_11204, mcs1_mcs_mat1_6_mcs_out[46]}), .c ({new_AGEMA_signal_16411, new_AGEMA_signal_16410, new_AGEMA_signal_16409, mcs1_mcs_mat1_6_n67}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U4 ( .a ({new_AGEMA_signal_14020, new_AGEMA_signal_14019, new_AGEMA_signal_14018, mcs1_mcs_mat1_6_mcs_out[34]}), .b ({new_AGEMA_signal_17938, new_AGEMA_signal_17937, new_AGEMA_signal_17936, mcs1_mcs_mat1_6_mcs_out[38]}), .c ({new_AGEMA_signal_18547, new_AGEMA_signal_18546, new_AGEMA_signal_18545, mcs1_mcs_mat1_6_n68}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U3 ( .a ({new_AGEMA_signal_17887, new_AGEMA_signal_17886, new_AGEMA_signal_17885, mcs1_mcs_mat1_6_n66}), .b ({new_AGEMA_signal_21703, new_AGEMA_signal_21702, new_AGEMA_signal_21701, mcs1_mcs_mat1_6_n65}), .c ({temp_next_s3[4], temp_next_s2[4], temp_next_s1[4], temp_next_s0[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U2 ( .a ({new_AGEMA_signal_21328, new_AGEMA_signal_21327, new_AGEMA_signal_21326, mcs1_mcs_mat1_6_mcs_out[4]}), .b ({new_AGEMA_signal_16489, new_AGEMA_signal_16488, new_AGEMA_signal_16487, mcs1_mcs_mat1_6_mcs_out[8]}), .c ({new_AGEMA_signal_21703, new_AGEMA_signal_21702, new_AGEMA_signal_21701, mcs1_mcs_mat1_6_n65}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_U1 ( .a ({new_AGEMA_signal_15502, new_AGEMA_signal_15501, new_AGEMA_signal_15500, mcs1_mcs_mat1_6_mcs_out[0]}), .b ({new_AGEMA_signal_17278, new_AGEMA_signal_17277, new_AGEMA_signal_17276, mcs1_mcs_mat1_6_mcs_out[12]}), .c ({new_AGEMA_signal_17887, new_AGEMA_signal_17886, new_AGEMA_signal_17885, mcs1_mcs_mat1_6_n66}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_15352, new_AGEMA_signal_15351, new_AGEMA_signal_15350, mcs1_mcs_mat1_6_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_16414, new_AGEMA_signal_16413, new_AGEMA_signal_16412, mcs1_mcs_mat1_6_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_13912, new_AGEMA_signal_13911, new_AGEMA_signal_13910, mcs1_mcs_mat1_6_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_9016, new_AGEMA_signal_9015, new_AGEMA_signal_9014, mcs1_mcs_mat1_6_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_15352, new_AGEMA_signal_15351, new_AGEMA_signal_15350, mcs1_mcs_mat1_6_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_9895, new_AGEMA_signal_9894, new_AGEMA_signal_9893, mcs1_mcs_mat1_6_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_11146, new_AGEMA_signal_11145, new_AGEMA_signal_11144, mcs1_mcs_mat1_6_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_12463, new_AGEMA_signal_12462, new_AGEMA_signal_12461, mcs1_mcs_mat1_6_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_9898, new_AGEMA_signal_9897, new_AGEMA_signal_9896, mcs1_mcs_mat1_6_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .c ({new_AGEMA_signal_11146, new_AGEMA_signal_11145, new_AGEMA_signal_11144, mcs1_mcs_mat1_6_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_15355, new_AGEMA_signal_15354, new_AGEMA_signal_15353, mcs1_mcs_mat1_6_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .c ({new_AGEMA_signal_16417, new_AGEMA_signal_16416, new_AGEMA_signal_16415, mcs1_mcs_mat1_6_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_13912, new_AGEMA_signal_13911, new_AGEMA_signal_13910, mcs1_mcs_mat1_6_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_15355, new_AGEMA_signal_15354, new_AGEMA_signal_15353, mcs1_mcs_mat1_6_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_12466, new_AGEMA_signal_12465, new_AGEMA_signal_12464, mcs1_mcs_mat1_6_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_11149, new_AGEMA_signal_11148, new_AGEMA_signal_11147, mcs1_mcs_mat1_6_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_13912, new_AGEMA_signal_13911, new_AGEMA_signal_13910, mcs1_mcs_mat1_6_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_13915, new_AGEMA_signal_13914, new_AGEMA_signal_13913, mcs1_mcs_mat1_6_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_15358, new_AGEMA_signal_15357, new_AGEMA_signal_15356, mcs1_mcs_mat1_6_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_12466, new_AGEMA_signal_12465, new_AGEMA_signal_12464, mcs1_mcs_mat1_6_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_9898, new_AGEMA_signal_9897, new_AGEMA_signal_9896, mcs1_mcs_mat1_6_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_13915, new_AGEMA_signal_13914, new_AGEMA_signal_13913, mcs1_mcs_mat1_6_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5717], Fresh[5716], Fresh[5715], Fresh[5714], Fresh[5713], Fresh[5712]}), .c ({new_AGEMA_signal_12466, new_AGEMA_signal_12465, new_AGEMA_signal_12464, mcs1_mcs_mat1_6_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5723], Fresh[5722], Fresh[5721], Fresh[5720], Fresh[5719], Fresh[5718]}), .c ({new_AGEMA_signal_9898, new_AGEMA_signal_9897, new_AGEMA_signal_9896, mcs1_mcs_mat1_6_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5729], Fresh[5728], Fresh[5727], Fresh[5726], Fresh[5725], Fresh[5724]}), .c ({new_AGEMA_signal_11149, new_AGEMA_signal_11148, new_AGEMA_signal_11147, mcs1_mcs_mat1_6_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_19216, new_AGEMA_signal_19215, new_AGEMA_signal_19214, mcs1_mcs_mat1_6_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .c ({new_AGEMA_signal_19942, new_AGEMA_signal_19941, new_AGEMA_signal_19940, mcs1_mcs_mat1_6_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_18550, new_AGEMA_signal_18549, new_AGEMA_signal_18548, mcs1_mcs_mat1_6_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_17236, new_AGEMA_signal_17235, new_AGEMA_signal_17234, mcs1_mcs_mat1_6_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_19216, new_AGEMA_signal_19215, new_AGEMA_signal_19214, mcs1_mcs_mat1_6_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_19219, new_AGEMA_signal_19218, new_AGEMA_signal_19217, mcs1_mcs_mat1_6_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_17893, new_AGEMA_signal_17892, new_AGEMA_signal_17891, mcs1_mcs_mat1_6_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_19945, new_AGEMA_signal_19944, new_AGEMA_signal_19943, mcs1_mcs_mat1_6_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_18550, new_AGEMA_signal_18549, new_AGEMA_signal_18548, mcs1_mcs_mat1_6_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .c ({new_AGEMA_signal_19219, new_AGEMA_signal_19218, new_AGEMA_signal_19217, mcs1_mcs_mat1_6_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_18550, new_AGEMA_signal_18549, new_AGEMA_signal_18548, mcs1_mcs_mat1_6_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_17890, new_AGEMA_signal_17889, new_AGEMA_signal_17888, mcs1_mcs_mat1_6_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_19222, new_AGEMA_signal_19221, new_AGEMA_signal_19220, mcs1_mcs_mat1_6_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_17896, new_AGEMA_signal_17895, new_AGEMA_signal_17894, mcs1_mcs_mat1_6_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_15361, new_AGEMA_signal_15360, new_AGEMA_signal_15359, mcs1_mcs_mat1_6_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_18550, new_AGEMA_signal_18549, new_AGEMA_signal_18548, mcs1_mcs_mat1_6_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_17233, new_AGEMA_signal_17232, new_AGEMA_signal_17231, mcs1_mcs_mat1_6_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_17893, new_AGEMA_signal_17892, new_AGEMA_signal_17891, mcs1_mcs_mat1_6_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_18553, new_AGEMA_signal_18552, new_AGEMA_signal_18551, mcs1_mcs_mat1_6_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_13918, new_AGEMA_signal_13917, new_AGEMA_signal_13916, mcs1_mcs_mat1_6_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_17236, new_AGEMA_signal_17235, new_AGEMA_signal_17234, mcs1_mcs_mat1_6_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_17893, new_AGEMA_signal_17892, new_AGEMA_signal_17891, mcs1_mcs_mat1_6_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_15361, new_AGEMA_signal_15360, new_AGEMA_signal_15359, mcs1_mcs_mat1_6_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_17233, new_AGEMA_signal_17232, new_AGEMA_signal_17231, mcs1_mcs_mat1_6_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5735], Fresh[5734], Fresh[5733], Fresh[5732], Fresh[5731], Fresh[5730]}), .c ({new_AGEMA_signal_17896, new_AGEMA_signal_17895, new_AGEMA_signal_17894, mcs1_mcs_mat1_6_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5741], Fresh[5740], Fresh[5739], Fresh[5738], Fresh[5737], Fresh[5736]}), .c ({new_AGEMA_signal_15361, new_AGEMA_signal_15360, new_AGEMA_signal_15359, mcs1_mcs_mat1_6_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5747], Fresh[5746], Fresh[5745], Fresh[5744], Fresh[5743], Fresh[5742]}), .c ({new_AGEMA_signal_17236, new_AGEMA_signal_17235, new_AGEMA_signal_17234, mcs1_mcs_mat1_6_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_13924, new_AGEMA_signal_13923, new_AGEMA_signal_13922, mcs1_mcs_mat1_6_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_9901, new_AGEMA_signal_9900, new_AGEMA_signal_9899, mcs1_mcs_mat1_6_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_15364, new_AGEMA_signal_15363, new_AGEMA_signal_15362, mcs1_mcs_mat1_6_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_11152, new_AGEMA_signal_11151, new_AGEMA_signal_11150, mcs1_mcs_mat1_6_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_11155, new_AGEMA_signal_11154, new_AGEMA_signal_11153, mcs1_mcs_mat1_6_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_12469, new_AGEMA_signal_12468, new_AGEMA_signal_12467, mcs1_mcs_mat1_6_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_13927, new_AGEMA_signal_13926, new_AGEMA_signal_13925, mcs1_mcs_mat1_6_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_15367, new_AGEMA_signal_15366, new_AGEMA_signal_15365, mcs1_mcs_mat1_6_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_16420, new_AGEMA_signal_16419, new_AGEMA_signal_16418, mcs1_mcs_mat1_6_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_13924, new_AGEMA_signal_13923, new_AGEMA_signal_13922, mcs1_mcs_mat1_6_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_15367, new_AGEMA_signal_15366, new_AGEMA_signal_15365, mcs1_mcs_mat1_6_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_9019, new_AGEMA_signal_9018, new_AGEMA_signal_9017, mcs1_mcs_mat1_6_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_12475, new_AGEMA_signal_12474, new_AGEMA_signal_12473, mcs1_mcs_mat1_6_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_13924, new_AGEMA_signal_13923, new_AGEMA_signal_13922, mcs1_mcs_mat1_6_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_9904, new_AGEMA_signal_9903, new_AGEMA_signal_9902, mcs1_mcs_mat1_6_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_12472, new_AGEMA_signal_12471, new_AGEMA_signal_12470, mcs1_mcs_mat1_6_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_13927, new_AGEMA_signal_13926, new_AGEMA_signal_13925, mcs1_mcs_mat1_6_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5753], Fresh[5752], Fresh[5751], Fresh[5750], Fresh[5749], Fresh[5748]}), .c ({new_AGEMA_signal_12475, new_AGEMA_signal_12474, new_AGEMA_signal_12473, mcs1_mcs_mat1_6_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5759], Fresh[5758], Fresh[5757], Fresh[5756], Fresh[5755], Fresh[5754]}), .c ({new_AGEMA_signal_9904, new_AGEMA_signal_9903, new_AGEMA_signal_9902, mcs1_mcs_mat1_6_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5765], Fresh[5764], Fresh[5763], Fresh[5762], Fresh[5761], Fresh[5760]}), .c ({new_AGEMA_signal_11155, new_AGEMA_signal_11154, new_AGEMA_signal_11153, mcs1_mcs_mat1_6_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({new_AGEMA_signal_15370, new_AGEMA_signal_15369, new_AGEMA_signal_15368, mcs1_mcs_mat1_6_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_16423, new_AGEMA_signal_16422, new_AGEMA_signal_16421, mcs1_mcs_mat1_6_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({new_AGEMA_signal_15373, new_AGEMA_signal_15372, new_AGEMA_signal_15371, mcs1_mcs_mat1_6_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_16426, new_AGEMA_signal_16425, new_AGEMA_signal_16424, mcs1_mcs_mat1_6_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_11158, new_AGEMA_signal_11157, new_AGEMA_signal_11156, mcs1_mcs_mat1_6_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_15370, new_AGEMA_signal_15369, new_AGEMA_signal_15368, mcs1_mcs_mat1_6_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_16429, new_AGEMA_signal_16428, new_AGEMA_signal_16427, mcs1_mcs_mat1_6_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_9907, new_AGEMA_signal_9906, new_AGEMA_signal_9905, mcs1_mcs_mat1_6_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_13930, new_AGEMA_signal_13929, new_AGEMA_signal_13928, mcs1_mcs_mat1_6_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_15370, new_AGEMA_signal_15369, new_AGEMA_signal_15368, mcs1_mcs_mat1_6_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_12478, new_AGEMA_signal_12477, new_AGEMA_signal_12476, mcs1_mcs_mat1_6_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_15373, new_AGEMA_signal_15372, new_AGEMA_signal_15371, mcs1_mcs_mat1_6_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_16432, new_AGEMA_signal_16431, new_AGEMA_signal_16430, mcs1_mcs_mat1_6_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_13933, new_AGEMA_signal_13932, new_AGEMA_signal_13931, mcs1_mcs_mat1_6_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_15373, new_AGEMA_signal_15372, new_AGEMA_signal_15371, mcs1_mcs_mat1_6_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_11158, new_AGEMA_signal_11157, new_AGEMA_signal_11156, mcs1_mcs_mat1_6_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_12481, new_AGEMA_signal_12480, new_AGEMA_signal_12479, mcs1_mcs_mat1_6_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_13933, new_AGEMA_signal_13932, new_AGEMA_signal_13931, mcs1_mcs_mat1_6_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5771], Fresh[5770], Fresh[5769], Fresh[5768], Fresh[5767], Fresh[5766]}), .c ({new_AGEMA_signal_12481, new_AGEMA_signal_12480, new_AGEMA_signal_12479, mcs1_mcs_mat1_6_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5777], Fresh[5776], Fresh[5775], Fresh[5774], Fresh[5773], Fresh[5772]}), .c ({new_AGEMA_signal_9907, new_AGEMA_signal_9906, new_AGEMA_signal_9905, mcs1_mcs_mat1_6_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5783], Fresh[5782], Fresh[5781], Fresh[5780], Fresh[5779], Fresh[5778]}), .c ({new_AGEMA_signal_11158, new_AGEMA_signal_11157, new_AGEMA_signal_11156, mcs1_mcs_mat1_6_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_13939, new_AGEMA_signal_13938, new_AGEMA_signal_13937, mcs1_mcs_mat1_6_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_13936, new_AGEMA_signal_13935, new_AGEMA_signal_13934, mcs1_mcs_mat1_6_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_15376, new_AGEMA_signal_15375, new_AGEMA_signal_15374, mcs1_mcs_mat1_6_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_13936, new_AGEMA_signal_13935, new_AGEMA_signal_13934, mcs1_mcs_mat1_6_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_11161, new_AGEMA_signal_11160, new_AGEMA_signal_11159, mcs1_mcs_mat1_6_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_15379, new_AGEMA_signal_15378, new_AGEMA_signal_15377, mcs1_mcs_mat1_6_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_9910, new_AGEMA_signal_9909, new_AGEMA_signal_9908, mcs1_mcs_mat1_6_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .c ({new_AGEMA_signal_11161, new_AGEMA_signal_11160, new_AGEMA_signal_11159, mcs1_mcs_mat1_6_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({new_AGEMA_signal_13936, new_AGEMA_signal_13935, new_AGEMA_signal_13934, mcs1_mcs_mat1_6_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_15382, new_AGEMA_signal_15381, new_AGEMA_signal_15380, mcs1_mcs_mat1_6_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_12487, new_AGEMA_signal_12486, new_AGEMA_signal_12485, mcs1_mcs_mat1_6_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_9025, new_AGEMA_signal_9024, new_AGEMA_signal_9023, mcs1_mcs_mat1_6_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_13936, new_AGEMA_signal_13935, new_AGEMA_signal_13934, mcs1_mcs_mat1_6_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_15385, new_AGEMA_signal_15384, new_AGEMA_signal_15383, mcs1_mcs_mat1_6_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_16435, new_AGEMA_signal_16434, new_AGEMA_signal_16433, mcs1_mcs_mat1_6_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_13939, new_AGEMA_signal_13938, new_AGEMA_signal_13937, mcs1_mcs_mat1_6_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_12487, new_AGEMA_signal_12486, new_AGEMA_signal_12485, mcs1_mcs_mat1_6_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_15385, new_AGEMA_signal_15384, new_AGEMA_signal_15383, mcs1_mcs_mat1_6_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_12484, new_AGEMA_signal_12483, new_AGEMA_signal_12482, mcs1_mcs_mat1_6_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .c ({new_AGEMA_signal_13939, new_AGEMA_signal_13938, new_AGEMA_signal_13937, mcs1_mcs_mat1_6_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_9910, new_AGEMA_signal_9909, new_AGEMA_signal_9908, mcs1_mcs_mat1_6_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_11164, new_AGEMA_signal_11163, new_AGEMA_signal_11162, mcs1_mcs_mat1_6_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_12484, new_AGEMA_signal_12483, new_AGEMA_signal_12482, mcs1_mcs_mat1_6_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5789], Fresh[5788], Fresh[5787], Fresh[5786], Fresh[5785], Fresh[5784]}), .c ({new_AGEMA_signal_12487, new_AGEMA_signal_12486, new_AGEMA_signal_12485, mcs1_mcs_mat1_6_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5795], Fresh[5794], Fresh[5793], Fresh[5792], Fresh[5791], Fresh[5790]}), .c ({new_AGEMA_signal_9910, new_AGEMA_signal_9909, new_AGEMA_signal_9908, mcs1_mcs_mat1_6_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5801], Fresh[5800], Fresh[5799], Fresh[5798], Fresh[5797], Fresh[5796]}), .c ({new_AGEMA_signal_11164, new_AGEMA_signal_11163, new_AGEMA_signal_11162, mcs1_mcs_mat1_6_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_17239, new_AGEMA_signal_17238, new_AGEMA_signal_17237, mcs1_mcs_mat1_6_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_18556, new_AGEMA_signal_18555, new_AGEMA_signal_18554, mcs1_mcs_mat1_6_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_19225, new_AGEMA_signal_19224, new_AGEMA_signal_19223, mcs1_mcs_mat1_6_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_17908, new_AGEMA_signal_17907, new_AGEMA_signal_17906, mcs1_mcs_mat1_6_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_18556, new_AGEMA_signal_18555, new_AGEMA_signal_18554, mcs1_mcs_mat1_6_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_17902, new_AGEMA_signal_17901, new_AGEMA_signal_17900, mcs1_mcs_mat1_6_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_17242, new_AGEMA_signal_17241, new_AGEMA_signal_17240, mcs1_mcs_mat1_6_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_18559, new_AGEMA_signal_18558, new_AGEMA_signal_18557, mcs1_mcs_mat1_6_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_17905, new_AGEMA_signal_17904, new_AGEMA_signal_17903, mcs1_mcs_mat1_6_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_18562, new_AGEMA_signal_18561, new_AGEMA_signal_18560, mcs1_mcs_mat1_6_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_19228, new_AGEMA_signal_19227, new_AGEMA_signal_19226, mcs1_mcs_mat1_6_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_13942, new_AGEMA_signal_13941, new_AGEMA_signal_13940, mcs1_mcs_mat1_6_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_17908, new_AGEMA_signal_17907, new_AGEMA_signal_17906, mcs1_mcs_mat1_6_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_18562, new_AGEMA_signal_18561, new_AGEMA_signal_18560, mcs1_mcs_mat1_6_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_15388, new_AGEMA_signal_15387, new_AGEMA_signal_15386, mcs1_mcs_mat1_6_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .c ({new_AGEMA_signal_17905, new_AGEMA_signal_17904, new_AGEMA_signal_17903, mcs1_mcs_mat1_6_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5807], Fresh[5806], Fresh[5805], Fresh[5804], Fresh[5803], Fresh[5802]}), .c ({new_AGEMA_signal_17908, new_AGEMA_signal_17907, new_AGEMA_signal_17906, mcs1_mcs_mat1_6_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5813], Fresh[5812], Fresh[5811], Fresh[5810], Fresh[5809], Fresh[5808]}), .c ({new_AGEMA_signal_15388, new_AGEMA_signal_15387, new_AGEMA_signal_15386, mcs1_mcs_mat1_6_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5819], Fresh[5818], Fresh[5817], Fresh[5816], Fresh[5815], Fresh[5814]}), .c ({new_AGEMA_signal_17242, new_AGEMA_signal_17241, new_AGEMA_signal_17240, mcs1_mcs_mat1_6_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_17245, new_AGEMA_signal_17244, new_AGEMA_signal_17243, mcs1_mcs_mat1_6_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_11170, new_AGEMA_signal_11169, new_AGEMA_signal_11168, mcs1_mcs_mat1_6_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_17911, new_AGEMA_signal_17910, new_AGEMA_signal_17909, mcs1_mcs_mat1_6_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_16438, new_AGEMA_signal_16437, new_AGEMA_signal_16436, mcs1_mcs_mat1_6_mcs_out[99]}), .b ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .c ({new_AGEMA_signal_17245, new_AGEMA_signal_17244, new_AGEMA_signal_17243, mcs1_mcs_mat1_6_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_15391, new_AGEMA_signal_15390, new_AGEMA_signal_15389, mcs1_mcs_mat1_6_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .c ({new_AGEMA_signal_16438, new_AGEMA_signal_16437, new_AGEMA_signal_16436, mcs1_mcs_mat1_6_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_13945, new_AGEMA_signal_13944, new_AGEMA_signal_13943, mcs1_mcs_mat1_6_mcs_out[98]}), .b ({new_AGEMA_signal_9916, new_AGEMA_signal_9915, new_AGEMA_signal_9914, mcs1_mcs_mat1_6_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_15391, new_AGEMA_signal_15390, new_AGEMA_signal_15389, mcs1_mcs_mat1_6_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_9913, new_AGEMA_signal_9912, new_AGEMA_signal_9911, mcs1_mcs_mat1_6_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_12490, new_AGEMA_signal_12489, new_AGEMA_signal_12488, mcs1_mcs_mat1_6_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_13945, new_AGEMA_signal_13944, new_AGEMA_signal_13943, mcs1_mcs_mat1_6_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5825], Fresh[5824], Fresh[5823], Fresh[5822], Fresh[5821], Fresh[5820]}), .c ({new_AGEMA_signal_12490, new_AGEMA_signal_12489, new_AGEMA_signal_12488, mcs1_mcs_mat1_6_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5831], Fresh[5830], Fresh[5829], Fresh[5828], Fresh[5827], Fresh[5826]}), .c ({new_AGEMA_signal_9916, new_AGEMA_signal_9915, new_AGEMA_signal_9914, mcs1_mcs_mat1_6_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5837], Fresh[5836], Fresh[5835], Fresh[5834], Fresh[5833], Fresh[5832]}), .c ({new_AGEMA_signal_11170, new_AGEMA_signal_11169, new_AGEMA_signal_11168, mcs1_mcs_mat1_6_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_13948, new_AGEMA_signal_13947, new_AGEMA_signal_13946, mcs1_mcs_mat1_6_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_15394, new_AGEMA_signal_15393, new_AGEMA_signal_15392, mcs1_mcs_mat1_6_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_11176, new_AGEMA_signal_11175, new_AGEMA_signal_11174, mcs1_mcs_mat1_6_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_11179, new_AGEMA_signal_11178, new_AGEMA_signal_11177, mcs1_mcs_mat1_6_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_12496, new_AGEMA_signal_12495, new_AGEMA_signal_12494, mcs1_mcs_mat1_6_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_15397, new_AGEMA_signal_15396, new_AGEMA_signal_15395, mcs1_mcs_mat1_6_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_9919, new_AGEMA_signal_9918, new_AGEMA_signal_9917, mcs1_mcs_mat1_6_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_16441, new_AGEMA_signal_16440, new_AGEMA_signal_16439, mcs1_mcs_mat1_6_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_13948, new_AGEMA_signal_13947, new_AGEMA_signal_13946, mcs1_mcs_mat1_6_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .c ({new_AGEMA_signal_15397, new_AGEMA_signal_15396, new_AGEMA_signal_15395, mcs1_mcs_mat1_6_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_9031, new_AGEMA_signal_9030, new_AGEMA_signal_9029, mcs1_mcs_mat1_6_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_12499, new_AGEMA_signal_12498, new_AGEMA_signal_12497, mcs1_mcs_mat1_6_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_13948, new_AGEMA_signal_13947, new_AGEMA_signal_13946, mcs1_mcs_mat1_6_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5843], Fresh[5842], Fresh[5841], Fresh[5840], Fresh[5839], Fresh[5838]}), .c ({new_AGEMA_signal_12499, new_AGEMA_signal_12498, new_AGEMA_signal_12497, mcs1_mcs_mat1_6_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5849], Fresh[5848], Fresh[5847], Fresh[5846], Fresh[5845], Fresh[5844]}), .c ({new_AGEMA_signal_9919, new_AGEMA_signal_9918, new_AGEMA_signal_9917, mcs1_mcs_mat1_6_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5855], Fresh[5854], Fresh[5853], Fresh[5852], Fresh[5851], Fresh[5850]}), .c ({new_AGEMA_signal_11179, new_AGEMA_signal_11178, new_AGEMA_signal_11177, mcs1_mcs_mat1_6_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_12508, new_AGEMA_signal_12507, new_AGEMA_signal_12506, mcs1_mcs_mat1_6_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_12511, new_AGEMA_signal_12510, new_AGEMA_signal_12509, mcs1_mcs_mat1_6_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_13951, new_AGEMA_signal_13950, new_AGEMA_signal_13949, mcs1_mcs_mat1_6_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_12502, new_AGEMA_signal_12501, new_AGEMA_signal_12500, mcs1_mcs_mat1_6_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_9034, new_AGEMA_signal_9033, new_AGEMA_signal_9032, mcs1_mcs_mat1_6_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_13954, new_AGEMA_signal_13953, new_AGEMA_signal_13952, mcs1_mcs_mat1_6_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_11188, new_AGEMA_signal_11187, new_AGEMA_signal_11186, mcs1_mcs_mat1_6_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_12502, new_AGEMA_signal_12501, new_AGEMA_signal_12500, mcs1_mcs_mat1_6_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_12505, new_AGEMA_signal_12504, new_AGEMA_signal_12503, mcs1_mcs_mat1_6_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_13957, new_AGEMA_signal_13956, new_AGEMA_signal_13955, mcs1_mcs_mat1_6_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_9922, new_AGEMA_signal_9921, new_AGEMA_signal_9920, mcs1_mcs_mat1_6_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_11188, new_AGEMA_signal_11187, new_AGEMA_signal_11186, mcs1_mcs_mat1_6_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_12505, new_AGEMA_signal_12504, new_AGEMA_signal_12503, mcs1_mcs_mat1_6_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_13960, new_AGEMA_signal_13959, new_AGEMA_signal_13958, mcs1_mcs_mat1_6_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .c ({new_AGEMA_signal_15400, new_AGEMA_signal_15399, new_AGEMA_signal_15398, mcs1_mcs_mat1_6_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_12508, new_AGEMA_signal_12507, new_AGEMA_signal_12506, mcs1_mcs_mat1_6_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_9922, new_AGEMA_signal_9921, new_AGEMA_signal_9920, mcs1_mcs_mat1_6_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_13960, new_AGEMA_signal_13959, new_AGEMA_signal_13958, mcs1_mcs_mat1_6_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5861], Fresh[5860], Fresh[5859], Fresh[5858], Fresh[5857], Fresh[5856]}), .c ({new_AGEMA_signal_12511, new_AGEMA_signal_12510, new_AGEMA_signal_12509, mcs1_mcs_mat1_6_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5867], Fresh[5866], Fresh[5865], Fresh[5864], Fresh[5863], Fresh[5862]}), .c ({new_AGEMA_signal_9922, new_AGEMA_signal_9921, new_AGEMA_signal_9920, mcs1_mcs_mat1_6_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5873], Fresh[5872], Fresh[5871], Fresh[5870], Fresh[5869], Fresh[5868]}), .c ({new_AGEMA_signal_11188, new_AGEMA_signal_11187, new_AGEMA_signal_11186, mcs1_mcs_mat1_6_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_13963, new_AGEMA_signal_13962, new_AGEMA_signal_13961, mcs1_mcs_mat1_6_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_15403, new_AGEMA_signal_15402, new_AGEMA_signal_15401, mcs1_mcs_mat1_6_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_11191, new_AGEMA_signal_11190, new_AGEMA_signal_11189, mcs1_mcs_mat1_6_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_12514, new_AGEMA_signal_12513, new_AGEMA_signal_12512, mcs1_mcs_mat1_6_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_15406, new_AGEMA_signal_15405, new_AGEMA_signal_15404, mcs1_mcs_mat1_6_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_9928, new_AGEMA_signal_9927, new_AGEMA_signal_9926, mcs1_mcs_mat1_6_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_16444, new_AGEMA_signal_16443, new_AGEMA_signal_16442, mcs1_mcs_mat1_6_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_13963, new_AGEMA_signal_13962, new_AGEMA_signal_13961, mcs1_mcs_mat1_6_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .c ({new_AGEMA_signal_15406, new_AGEMA_signal_15405, new_AGEMA_signal_15404, mcs1_mcs_mat1_6_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_9037, new_AGEMA_signal_9036, new_AGEMA_signal_9035, mcs1_mcs_mat1_6_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_12517, new_AGEMA_signal_12516, new_AGEMA_signal_12515, mcs1_mcs_mat1_6_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_13963, new_AGEMA_signal_13962, new_AGEMA_signal_13961, mcs1_mcs_mat1_6_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5879], Fresh[5878], Fresh[5877], Fresh[5876], Fresh[5875], Fresh[5874]}), .c ({new_AGEMA_signal_12517, new_AGEMA_signal_12516, new_AGEMA_signal_12515, mcs1_mcs_mat1_6_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5885], Fresh[5884], Fresh[5883], Fresh[5882], Fresh[5881], Fresh[5880]}), .c ({new_AGEMA_signal_9928, new_AGEMA_signal_9927, new_AGEMA_signal_9926, mcs1_mcs_mat1_6_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5891], Fresh[5890], Fresh[5889], Fresh[5888], Fresh[5887], Fresh[5886]}), .c ({new_AGEMA_signal_11191, new_AGEMA_signal_11190, new_AGEMA_signal_11189, mcs1_mcs_mat1_6_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_15409, new_AGEMA_signal_15408, new_AGEMA_signal_15407, mcs1_mcs_mat1_6_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_16447, new_AGEMA_signal_16446, new_AGEMA_signal_16445, mcs1_mcs_mat1_6_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_13969, new_AGEMA_signal_13968, new_AGEMA_signal_13967, mcs1_mcs_mat1_6_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_12523, new_AGEMA_signal_12522, new_AGEMA_signal_12521, mcs1_mcs_mat1_6_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_15409, new_AGEMA_signal_15408, new_AGEMA_signal_15407, mcs1_mcs_mat1_6_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({new_AGEMA_signal_10345, new_AGEMA_signal_10344, new_AGEMA_signal_10343, mcs1_mcs_mat1_6_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_12520, new_AGEMA_signal_12519, new_AGEMA_signal_12518, mcs1_mcs_mat1_6_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_12523, new_AGEMA_signal_12522, new_AGEMA_signal_12521, mcs1_mcs_mat1_6_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_10345, new_AGEMA_signal_10344, new_AGEMA_signal_10343, mcs1_mcs_mat1_6_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_13966, new_AGEMA_signal_13965, new_AGEMA_signal_13964, mcs1_mcs_mat1_6_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_9931, new_AGEMA_signal_9930, new_AGEMA_signal_9929, mcs1_mcs_mat1_6_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_9934, new_AGEMA_signal_9933, new_AGEMA_signal_9932, mcs1_mcs_mat1_6_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_10345, new_AGEMA_signal_10344, new_AGEMA_signal_10343, mcs1_mcs_mat1_6_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_11194, new_AGEMA_signal_11193, new_AGEMA_signal_11192, mcs1_mcs_mat1_6_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .c ({new_AGEMA_signal_12523, new_AGEMA_signal_12522, new_AGEMA_signal_12521, mcs1_mcs_mat1_6_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_15412, new_AGEMA_signal_15411, new_AGEMA_signal_15410, mcs1_mcs_mat1_6_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_9931, new_AGEMA_signal_9930, new_AGEMA_signal_9929, mcs1_mcs_mat1_6_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_16450, new_AGEMA_signal_16449, new_AGEMA_signal_16448, mcs1_mcs_mat1_6_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_13969, new_AGEMA_signal_13968, new_AGEMA_signal_13967, mcs1_mcs_mat1_6_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_11194, new_AGEMA_signal_11193, new_AGEMA_signal_11192, mcs1_mcs_mat1_6_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_15412, new_AGEMA_signal_15411, new_AGEMA_signal_15410, mcs1_mcs_mat1_6_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .b ({new_AGEMA_signal_12526, new_AGEMA_signal_12525, new_AGEMA_signal_12524, mcs1_mcs_mat1_6_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_13969, new_AGEMA_signal_13968, new_AGEMA_signal_13967, mcs1_mcs_mat1_6_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5897], Fresh[5896], Fresh[5895], Fresh[5894], Fresh[5893], Fresh[5892]}), .c ({new_AGEMA_signal_12526, new_AGEMA_signal_12525, new_AGEMA_signal_12524, mcs1_mcs_mat1_6_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5903], Fresh[5902], Fresh[5901], Fresh[5900], Fresh[5899], Fresh[5898]}), .c ({new_AGEMA_signal_9934, new_AGEMA_signal_9933, new_AGEMA_signal_9932, mcs1_mcs_mat1_6_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5909], Fresh[5908], Fresh[5907], Fresh[5906], Fresh[5905], Fresh[5904]}), .c ({new_AGEMA_signal_11194, new_AGEMA_signal_11193, new_AGEMA_signal_11192, mcs1_mcs_mat1_6_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_18568, new_AGEMA_signal_18567, new_AGEMA_signal_18566, mcs1_mcs_mat1_6_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_17248, new_AGEMA_signal_17247, new_AGEMA_signal_17246, mcs1_mcs_mat1_6_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_19231, new_AGEMA_signal_19230, new_AGEMA_signal_19229, mcs1_mcs_mat1_6_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_17920, new_AGEMA_signal_17919, new_AGEMA_signal_17918, mcs1_mcs_mat1_6_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_19234, new_AGEMA_signal_19233, new_AGEMA_signal_19232, mcs1_mcs_mat1_6_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_19948, new_AGEMA_signal_19947, new_AGEMA_signal_19946, mcs1_mcs_mat1_6_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_18568, new_AGEMA_signal_18567, new_AGEMA_signal_18566, mcs1_mcs_mat1_6_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_19234, new_AGEMA_signal_19233, new_AGEMA_signal_19232, mcs1_mcs_mat1_6_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_19951, new_AGEMA_signal_19950, new_AGEMA_signal_19949, mcs1_mcs_mat1_6_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_17248, new_AGEMA_signal_17247, new_AGEMA_signal_17246, mcs1_mcs_mat1_6_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_18571, new_AGEMA_signal_18570, new_AGEMA_signal_18569, mcs1_mcs_mat1_6_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_19234, new_AGEMA_signal_19233, new_AGEMA_signal_19232, mcs1_mcs_mat1_6_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({new_AGEMA_signal_15415, new_AGEMA_signal_15414, new_AGEMA_signal_15413, mcs1_mcs_mat1_6_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_17248, new_AGEMA_signal_17247, new_AGEMA_signal_17246, mcs1_mcs_mat1_6_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_17917, new_AGEMA_signal_17916, new_AGEMA_signal_17915, mcs1_mcs_mat1_6_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .c ({new_AGEMA_signal_18568, new_AGEMA_signal_18567, new_AGEMA_signal_18566, mcs1_mcs_mat1_6_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_17251, new_AGEMA_signal_17250, new_AGEMA_signal_17249, mcs1_mcs_mat1_6_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_13972, new_AGEMA_signal_13971, new_AGEMA_signal_13970, mcs1_mcs_mat1_6_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_17917, new_AGEMA_signal_17916, new_AGEMA_signal_17915, mcs1_mcs_mat1_6_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_18571, new_AGEMA_signal_18570, new_AGEMA_signal_18569, mcs1_mcs_mat1_6_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_17920, new_AGEMA_signal_17919, new_AGEMA_signal_17918, mcs1_mcs_mat1_6_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_19237, new_AGEMA_signal_19236, new_AGEMA_signal_19235, mcs1_mcs_mat1_6_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_17251, new_AGEMA_signal_17250, new_AGEMA_signal_17249, mcs1_mcs_mat1_6_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_17920, new_AGEMA_signal_17919, new_AGEMA_signal_17918, mcs1_mcs_mat1_6_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({new_AGEMA_signal_17923, new_AGEMA_signal_17922, new_AGEMA_signal_17921, mcs1_mcs_mat1_6_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_18571, new_AGEMA_signal_18570, new_AGEMA_signal_18569, mcs1_mcs_mat1_6_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5915], Fresh[5914], Fresh[5913], Fresh[5912], Fresh[5911], Fresh[5910]}), .c ({new_AGEMA_signal_17923, new_AGEMA_signal_17922, new_AGEMA_signal_17921, mcs1_mcs_mat1_6_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5921], Fresh[5920], Fresh[5919], Fresh[5918], Fresh[5917], Fresh[5916]}), .c ({new_AGEMA_signal_15415, new_AGEMA_signal_15414, new_AGEMA_signal_15413, mcs1_mcs_mat1_6_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5927], Fresh[5926], Fresh[5925], Fresh[5924], Fresh[5923], Fresh[5922]}), .c ({new_AGEMA_signal_17251, new_AGEMA_signal_17250, new_AGEMA_signal_17249, mcs1_mcs_mat1_6_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_15421, new_AGEMA_signal_15420, new_AGEMA_signal_15419, mcs1_mcs_mat1_6_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .c ({new_AGEMA_signal_16453, new_AGEMA_signal_16452, new_AGEMA_signal_16451, mcs1_mcs_mat1_6_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({new_AGEMA_signal_13975, new_AGEMA_signal_13974, new_AGEMA_signal_13973, mcs1_mcs_mat1_6_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_15418, new_AGEMA_signal_15417, new_AGEMA_signal_15416, mcs1_mcs_mat1_6_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_16456, new_AGEMA_signal_16455, new_AGEMA_signal_16454, mcs1_mcs_mat1_6_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_11197, new_AGEMA_signal_11196, new_AGEMA_signal_11195, mcs1_mcs_mat1_6_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_17254, new_AGEMA_signal_17253, new_AGEMA_signal_17252, mcs1_mcs_mat1_6_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_15421, new_AGEMA_signal_15420, new_AGEMA_signal_15419, mcs1_mcs_mat1_6_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .c ({new_AGEMA_signal_16456, new_AGEMA_signal_16455, new_AGEMA_signal_16454, mcs1_mcs_mat1_6_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_9937, new_AGEMA_signal_9936, new_AGEMA_signal_9935, mcs1_mcs_mat1_6_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_13975, new_AGEMA_signal_13974, new_AGEMA_signal_13973, mcs1_mcs_mat1_6_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_15421, new_AGEMA_signal_15420, new_AGEMA_signal_15419, mcs1_mcs_mat1_6_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_9043, new_AGEMA_signal_9042, new_AGEMA_signal_9041, mcs1_mcs_mat1_6_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_12532, new_AGEMA_signal_12531, new_AGEMA_signal_12530, mcs1_mcs_mat1_6_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_13975, new_AGEMA_signal_13974, new_AGEMA_signal_13973, mcs1_mcs_mat1_6_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5933], Fresh[5932], Fresh[5931], Fresh[5930], Fresh[5929], Fresh[5928]}), .c ({new_AGEMA_signal_12532, new_AGEMA_signal_12531, new_AGEMA_signal_12530, mcs1_mcs_mat1_6_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5939], Fresh[5938], Fresh[5937], Fresh[5936], Fresh[5935], Fresh[5934]}), .c ({new_AGEMA_signal_9937, new_AGEMA_signal_9936, new_AGEMA_signal_9935, mcs1_mcs_mat1_6_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5945], Fresh[5944], Fresh[5943], Fresh[5942], Fresh[5941], Fresh[5940]}), .c ({new_AGEMA_signal_11197, new_AGEMA_signal_11196, new_AGEMA_signal_11195, mcs1_mcs_mat1_6_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_13984, new_AGEMA_signal_13983, new_AGEMA_signal_13982, mcs1_mcs_mat1_6_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_11200, new_AGEMA_signal_11199, new_AGEMA_signal_11198, mcs1_mcs_mat1_6_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_15424, new_AGEMA_signal_15423, new_AGEMA_signal_15422, mcs1_mcs_mat1_6_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_9940, new_AGEMA_signal_9939, new_AGEMA_signal_9938, mcs1_mcs_mat1_6_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_12535, new_AGEMA_signal_12534, new_AGEMA_signal_12533, mcs1_mcs_mat1_6_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_13978, new_AGEMA_signal_13977, new_AGEMA_signal_13976, mcs1_mcs_mat1_6_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({new_AGEMA_signal_12538, new_AGEMA_signal_12537, new_AGEMA_signal_12536, mcs1_mcs_mat1_6_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_13981, new_AGEMA_signal_13980, new_AGEMA_signal_13979, mcs1_mcs_mat1_6_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5951], Fresh[5950], Fresh[5949], Fresh[5948], Fresh[5947], Fresh[5946]}), .c ({new_AGEMA_signal_12538, new_AGEMA_signal_12537, new_AGEMA_signal_12536, mcs1_mcs_mat1_6_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5957], Fresh[5956], Fresh[5955], Fresh[5954], Fresh[5953], Fresh[5952]}), .c ({new_AGEMA_signal_9940, new_AGEMA_signal_9939, new_AGEMA_signal_9938, mcs1_mcs_mat1_6_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5963], Fresh[5962], Fresh[5961], Fresh[5960], Fresh[5959], Fresh[5958]}), .c ({new_AGEMA_signal_11200, new_AGEMA_signal_11199, new_AGEMA_signal_11198, mcs1_mcs_mat1_6_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_9946, new_AGEMA_signal_9945, new_AGEMA_signal_9944, mcs1_mcs_mat1_6_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_11203, new_AGEMA_signal_11202, new_AGEMA_signal_11201, mcs1_mcs_mat1_6_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_12541, new_AGEMA_signal_12540, new_AGEMA_signal_12539, mcs1_mcs_mat1_6_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_9949, new_AGEMA_signal_9948, new_AGEMA_signal_9947, mcs1_mcs_mat1_6_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_12544, new_AGEMA_signal_12543, new_AGEMA_signal_12542, mcs1_mcs_mat1_6_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_13990, new_AGEMA_signal_13989, new_AGEMA_signal_13988, mcs1_mcs_mat1_6_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_13993, new_AGEMA_signal_13992, new_AGEMA_signal_13991, mcs1_mcs_mat1_6_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_12547, new_AGEMA_signal_12546, new_AGEMA_signal_12545, mcs1_mcs_mat1_6_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_15430, new_AGEMA_signal_15429, new_AGEMA_signal_15428, mcs1_mcs_mat1_6_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_12550, new_AGEMA_signal_12549, new_AGEMA_signal_12548, mcs1_mcs_mat1_6_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_13993, new_AGEMA_signal_13992, new_AGEMA_signal_13991, mcs1_mcs_mat1_6_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5969], Fresh[5968], Fresh[5967], Fresh[5966], Fresh[5965], Fresh[5964]}), .c ({new_AGEMA_signal_12550, new_AGEMA_signal_12549, new_AGEMA_signal_12548, mcs1_mcs_mat1_6_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5975], Fresh[5974], Fresh[5973], Fresh[5972], Fresh[5971], Fresh[5970]}), .c ({new_AGEMA_signal_9949, new_AGEMA_signal_9948, new_AGEMA_signal_9947, mcs1_mcs_mat1_6_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5981], Fresh[5980], Fresh[5979], Fresh[5978], Fresh[5977], Fresh[5976]}), .c ({new_AGEMA_signal_11203, new_AGEMA_signal_11202, new_AGEMA_signal_11201, mcs1_mcs_mat1_6_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_17929, new_AGEMA_signal_17928, new_AGEMA_signal_17927, mcs1_mcs_mat1_6_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_18574, new_AGEMA_signal_18573, new_AGEMA_signal_18572, mcs1_mcs_mat1_6_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_19240, new_AGEMA_signal_19239, new_AGEMA_signal_19238, mcs1_mcs_mat1_6_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_19243, new_AGEMA_signal_19242, new_AGEMA_signal_19241, mcs1_mcs_mat1_6_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_17926, new_AGEMA_signal_17925, new_AGEMA_signal_17924, mcs1_mcs_mat1_6_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_19954, new_AGEMA_signal_19953, new_AGEMA_signal_19952, mcs1_mcs_mat1_6_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_17257, new_AGEMA_signal_17256, new_AGEMA_signal_17255, mcs1_mcs_mat1_6_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_17926, new_AGEMA_signal_17925, new_AGEMA_signal_17924, mcs1_mcs_mat1_6_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({new_AGEMA_signal_19243, new_AGEMA_signal_19242, new_AGEMA_signal_19241, mcs1_mcs_mat1_6_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_19957, new_AGEMA_signal_19956, new_AGEMA_signal_19955, mcs1_mcs_mat1_6_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_13996, new_AGEMA_signal_13995, new_AGEMA_signal_13994, mcs1_mcs_mat1_6_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_18574, new_AGEMA_signal_18573, new_AGEMA_signal_18572, mcs1_mcs_mat1_6_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_19243, new_AGEMA_signal_19242, new_AGEMA_signal_19241, mcs1_mcs_mat1_6_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_15433, new_AGEMA_signal_15432, new_AGEMA_signal_15431, mcs1_mcs_mat1_6_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_17935, new_AGEMA_signal_17934, new_AGEMA_signal_17933, mcs1_mcs_mat1_6_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_18574, new_AGEMA_signal_18573, new_AGEMA_signal_18572, mcs1_mcs_mat1_6_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_17932, new_AGEMA_signal_17931, new_AGEMA_signal_17930, mcs1_mcs_mat1_6_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_18577, new_AGEMA_signal_18576, new_AGEMA_signal_18575, mcs1_mcs_mat1_6_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_19246, new_AGEMA_signal_19245, new_AGEMA_signal_19244, mcs1_mcs_mat1_6_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_17929, new_AGEMA_signal_17928, new_AGEMA_signal_17927, mcs1_mcs_mat1_6_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_15433, new_AGEMA_signal_15432, new_AGEMA_signal_15431, mcs1_mcs_mat1_6_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_18577, new_AGEMA_signal_18576, new_AGEMA_signal_18575, mcs1_mcs_mat1_6_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_17257, new_AGEMA_signal_17256, new_AGEMA_signal_17255, mcs1_mcs_mat1_6_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_17929, new_AGEMA_signal_17928, new_AGEMA_signal_17927, mcs1_mcs_mat1_6_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5987], Fresh[5986], Fresh[5985], Fresh[5984], Fresh[5983], Fresh[5982]}), .c ({new_AGEMA_signal_17935, new_AGEMA_signal_17934, new_AGEMA_signal_17933, mcs1_mcs_mat1_6_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5993], Fresh[5992], Fresh[5991], Fresh[5990], Fresh[5989], Fresh[5988]}), .c ({new_AGEMA_signal_15433, new_AGEMA_signal_15432, new_AGEMA_signal_15431, mcs1_mcs_mat1_6_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[5999], Fresh[5998], Fresh[5997], Fresh[5996], Fresh[5995], Fresh[5994]}), .c ({new_AGEMA_signal_17257, new_AGEMA_signal_17256, new_AGEMA_signal_17255, mcs1_mcs_mat1_6_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_11209, new_AGEMA_signal_11208, new_AGEMA_signal_11207, mcs1_mcs_mat1_6_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_12556, new_AGEMA_signal_12555, new_AGEMA_signal_12554, mcs1_mcs_mat1_6_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_16462, new_AGEMA_signal_16461, new_AGEMA_signal_16460, mcs1_mcs_mat1_6_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_9952, new_AGEMA_signal_9951, new_AGEMA_signal_9950, mcs1_mcs_mat1_6_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_17260, new_AGEMA_signal_17259, new_AGEMA_signal_17258, mcs1_mcs_mat1_6_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_15436, new_AGEMA_signal_15435, new_AGEMA_signal_15434, mcs1_mcs_mat1_6_mcs_out[47]}), .b ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .c ({new_AGEMA_signal_16462, new_AGEMA_signal_16461, new_AGEMA_signal_16460, mcs1_mcs_mat1_6_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_14002, new_AGEMA_signal_14001, new_AGEMA_signal_14000, mcs1_mcs_mat1_6_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .c ({new_AGEMA_signal_15436, new_AGEMA_signal_15435, new_AGEMA_signal_15434, mcs1_mcs_mat1_6_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_9052, new_AGEMA_signal_9051, new_AGEMA_signal_9050, mcs1_mcs_mat1_6_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_12559, new_AGEMA_signal_12558, new_AGEMA_signal_12557, mcs1_mcs_mat1_6_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_14002, new_AGEMA_signal_14001, new_AGEMA_signal_14000, mcs1_mcs_mat1_6_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6005], Fresh[6004], Fresh[6003], Fresh[6002], Fresh[6001], Fresh[6000]}), .c ({new_AGEMA_signal_12559, new_AGEMA_signal_12558, new_AGEMA_signal_12557, mcs1_mcs_mat1_6_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6011], Fresh[6010], Fresh[6009], Fresh[6008], Fresh[6007], Fresh[6006]}), .c ({new_AGEMA_signal_9952, new_AGEMA_signal_9951, new_AGEMA_signal_9950, mcs1_mcs_mat1_6_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6017], Fresh[6016], Fresh[6015], Fresh[6014], Fresh[6013], Fresh[6012]}), .c ({new_AGEMA_signal_11209, new_AGEMA_signal_11208, new_AGEMA_signal_11207, mcs1_mcs_mat1_6_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_14005, new_AGEMA_signal_14004, new_AGEMA_signal_14003, mcs1_mcs_mat1_6_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_11212, new_AGEMA_signal_11211, new_AGEMA_signal_11210, mcs1_mcs_mat1_6_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_15439, new_AGEMA_signal_15438, new_AGEMA_signal_15437, mcs1_mcs_mat1_6_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_12562, new_AGEMA_signal_12561, new_AGEMA_signal_12560, mcs1_mcs_mat1_6_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_9955, new_AGEMA_signal_9954, new_AGEMA_signal_9953, mcs1_mcs_mat1_6_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_14005, new_AGEMA_signal_14004, new_AGEMA_signal_14003, mcs1_mcs_mat1_6_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_14008, new_AGEMA_signal_14007, new_AGEMA_signal_14006, mcs1_mcs_mat1_6_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_12568, new_AGEMA_signal_12567, new_AGEMA_signal_12566, mcs1_mcs_mat1_6_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_15442, new_AGEMA_signal_15441, new_AGEMA_signal_15440, mcs1_mcs_mat1_6_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_14011, new_AGEMA_signal_14010, new_AGEMA_signal_14009, mcs1_mcs_mat1_6_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_9055, new_AGEMA_signal_9054, new_AGEMA_signal_9053, mcs1_mcs_mat1_6_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_15445, new_AGEMA_signal_15444, new_AGEMA_signal_15443, mcs1_mcs_mat1_6_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_12562, new_AGEMA_signal_12561, new_AGEMA_signal_12560, mcs1_mcs_mat1_6_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_11215, new_AGEMA_signal_11214, new_AGEMA_signal_11213, mcs1_mcs_mat1_6_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_14011, new_AGEMA_signal_14010, new_AGEMA_signal_14009, mcs1_mcs_mat1_6_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_12565, new_AGEMA_signal_12564, new_AGEMA_signal_12563, mcs1_mcs_mat1_6_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_11215, new_AGEMA_signal_11214, new_AGEMA_signal_11213, mcs1_mcs_mat1_6_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_14014, new_AGEMA_signal_14013, new_AGEMA_signal_14012, mcs1_mcs_mat1_6_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6023], Fresh[6022], Fresh[6021], Fresh[6020], Fresh[6019], Fresh[6018]}), .c ({new_AGEMA_signal_12568, new_AGEMA_signal_12567, new_AGEMA_signal_12566, mcs1_mcs_mat1_6_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6029], Fresh[6028], Fresh[6027], Fresh[6026], Fresh[6025], Fresh[6024]}), .c ({new_AGEMA_signal_9955, new_AGEMA_signal_9954, new_AGEMA_signal_9953, mcs1_mcs_mat1_6_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6035], Fresh[6034], Fresh[6033], Fresh[6032], Fresh[6031], Fresh[6030]}), .c ({new_AGEMA_signal_11215, new_AGEMA_signal_11214, new_AGEMA_signal_11213, mcs1_mcs_mat1_6_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_19249, new_AGEMA_signal_19248, new_AGEMA_signal_19247, mcs1_mcs_mat1_6_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_14017, new_AGEMA_signal_14016, new_AGEMA_signal_14015, mcs1_mcs_mat1_6_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_19960, new_AGEMA_signal_19959, new_AGEMA_signal_19958, mcs1_mcs_mat1_6_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_17266, new_AGEMA_signal_17265, new_AGEMA_signal_17264, mcs1_mcs_mat1_6_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_17263, new_AGEMA_signal_17262, new_AGEMA_signal_17261, mcs1_mcs_mat1_6_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_17938, new_AGEMA_signal_17937, new_AGEMA_signal_17936, mcs1_mcs_mat1_6_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({new_AGEMA_signal_19249, new_AGEMA_signal_19248, new_AGEMA_signal_19247, mcs1_mcs_mat1_6_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_19963, new_AGEMA_signal_19962, new_AGEMA_signal_19961, mcs1_mcs_mat1_6_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_17941, new_AGEMA_signal_17940, new_AGEMA_signal_17939, mcs1_mcs_mat1_6_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_18580, new_AGEMA_signal_18579, new_AGEMA_signal_18578, mcs1_mcs_mat1_6_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_19249, new_AGEMA_signal_19248, new_AGEMA_signal_19247, mcs1_mcs_mat1_6_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_17944, new_AGEMA_signal_17943, new_AGEMA_signal_17942, mcs1_mcs_mat1_6_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_17269, new_AGEMA_signal_17268, new_AGEMA_signal_17267, mcs1_mcs_mat1_6_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_18580, new_AGEMA_signal_18579, new_AGEMA_signal_18578, mcs1_mcs_mat1_6_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_17944, new_AGEMA_signal_17943, new_AGEMA_signal_17942, mcs1_mcs_mat1_6_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_17266, new_AGEMA_signal_17265, new_AGEMA_signal_17264, mcs1_mcs_mat1_6_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_18583, new_AGEMA_signal_18582, new_AGEMA_signal_18581, mcs1_mcs_mat1_6_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .b ({new_AGEMA_signal_16465, new_AGEMA_signal_16464, new_AGEMA_signal_16463, mcs1_mcs_mat1_6_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_17266, new_AGEMA_signal_17265, new_AGEMA_signal_17264, mcs1_mcs_mat1_6_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({new_AGEMA_signal_15448, new_AGEMA_signal_15447, new_AGEMA_signal_15446, mcs1_mcs_mat1_6_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_16465, new_AGEMA_signal_16464, new_AGEMA_signal_16463, mcs1_mcs_mat1_6_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6041], Fresh[6040], Fresh[6039], Fresh[6038], Fresh[6037], Fresh[6036]}), .c ({new_AGEMA_signal_17944, new_AGEMA_signal_17943, new_AGEMA_signal_17942, mcs1_mcs_mat1_6_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6047], Fresh[6046], Fresh[6045], Fresh[6044], Fresh[6043], Fresh[6042]}), .c ({new_AGEMA_signal_15448, new_AGEMA_signal_15447, new_AGEMA_signal_15446, mcs1_mcs_mat1_6_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6053], Fresh[6052], Fresh[6051], Fresh[6050], Fresh[6049], Fresh[6048]}), .c ({new_AGEMA_signal_17269, new_AGEMA_signal_17268, new_AGEMA_signal_17267, mcs1_mcs_mat1_6_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_12571, new_AGEMA_signal_12570, new_AGEMA_signal_12569, mcs1_mcs_mat1_6_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_11218, new_AGEMA_signal_11217, new_AGEMA_signal_11216, mcs1_mcs_mat1_6_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_14020, new_AGEMA_signal_14019, new_AGEMA_signal_14018, mcs1_mcs_mat1_6_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, new_AGEMA_signal_9956, mcs1_mcs_mat1_6_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_10348, new_AGEMA_signal_10347, new_AGEMA_signal_10346, mcs1_mcs_mat1_6_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_16468, new_AGEMA_signal_16467, new_AGEMA_signal_16466, mcs1_mcs_mat1_6_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_12574, new_AGEMA_signal_12573, new_AGEMA_signal_12572, mcs1_mcs_mat1_6_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_17272, new_AGEMA_signal_17271, new_AGEMA_signal_17270, mcs1_mcs_mat1_6_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6059], Fresh[6058], Fresh[6057], Fresh[6056], Fresh[6055], Fresh[6054]}), .c ({new_AGEMA_signal_12574, new_AGEMA_signal_12573, new_AGEMA_signal_12572, mcs1_mcs_mat1_6_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6065], Fresh[6064], Fresh[6063], Fresh[6062], Fresh[6061], Fresh[6060]}), .c ({new_AGEMA_signal_9958, new_AGEMA_signal_9957, new_AGEMA_signal_9956, mcs1_mcs_mat1_6_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6071], Fresh[6070], Fresh[6069], Fresh[6068], Fresh[6067], Fresh[6066]}), .c ({new_AGEMA_signal_11218, new_AGEMA_signal_11217, new_AGEMA_signal_11216, mcs1_mcs_mat1_6_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_15454, new_AGEMA_signal_15453, new_AGEMA_signal_15452, mcs1_mcs_mat1_6_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_14026, new_AGEMA_signal_14025, new_AGEMA_signal_14024, mcs1_mcs_mat1_6_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_16471, new_AGEMA_signal_16470, new_AGEMA_signal_16469, mcs1_mcs_mat1_6_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_9964, new_AGEMA_signal_9963, new_AGEMA_signal_9962, mcs1_mcs_mat1_6_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_14029, new_AGEMA_signal_14028, new_AGEMA_signal_14027, mcs1_mcs_mat1_6_mcs_out[29]}), .c ({new_AGEMA_signal_15454, new_AGEMA_signal_15453, new_AGEMA_signal_15452, mcs1_mcs_mat1_6_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_9961, new_AGEMA_signal_9960, new_AGEMA_signal_9959, mcs1_mcs_mat1_6_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_14026, new_AGEMA_signal_14025, new_AGEMA_signal_14024, mcs1_mcs_mat1_6_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_15457, new_AGEMA_signal_15456, new_AGEMA_signal_15455, mcs1_mcs_mat1_6_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_12583, new_AGEMA_signal_12582, new_AGEMA_signal_12581, mcs1_mcs_mat1_6_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .c ({new_AGEMA_signal_14026, new_AGEMA_signal_14025, new_AGEMA_signal_14024, mcs1_mcs_mat1_6_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_15460, new_AGEMA_signal_15459, new_AGEMA_signal_15458, mcs1_mcs_mat1_6_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_12577, new_AGEMA_signal_12576, new_AGEMA_signal_12575, mcs1_mcs_mat1_6_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_16474, new_AGEMA_signal_16473, new_AGEMA_signal_16472, mcs1_mcs_mat1_6_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_14032, new_AGEMA_signal_14031, new_AGEMA_signal_14030, mcs1_mcs_mat1_6_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_12580, new_AGEMA_signal_12579, new_AGEMA_signal_12578, mcs1_mcs_mat1_6_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_15460, new_AGEMA_signal_15459, new_AGEMA_signal_15458, mcs1_mcs_mat1_6_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_11221, new_AGEMA_signal_11220, new_AGEMA_signal_11219, mcs1_mcs_mat1_6_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_12580, new_AGEMA_signal_12579, new_AGEMA_signal_12578, mcs1_mcs_mat1_6_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_12583, new_AGEMA_signal_12582, new_AGEMA_signal_12581, mcs1_mcs_mat1_6_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_9964, new_AGEMA_signal_9963, new_AGEMA_signal_9962, mcs1_mcs_mat1_6_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_14032, new_AGEMA_signal_14031, new_AGEMA_signal_14030, mcs1_mcs_mat1_6_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6077], Fresh[6076], Fresh[6075], Fresh[6074], Fresh[6073], Fresh[6072]}), .c ({new_AGEMA_signal_12583, new_AGEMA_signal_12582, new_AGEMA_signal_12581, mcs1_mcs_mat1_6_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6083], Fresh[6082], Fresh[6081], Fresh[6080], Fresh[6079], Fresh[6078]}), .c ({new_AGEMA_signal_9964, new_AGEMA_signal_9963, new_AGEMA_signal_9962, mcs1_mcs_mat1_6_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6089], Fresh[6088], Fresh[6087], Fresh[6086], Fresh[6085], Fresh[6084]}), .c ({new_AGEMA_signal_11221, new_AGEMA_signal_11220, new_AGEMA_signal_11219, mcs1_mcs_mat1_6_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_12586, new_AGEMA_signal_12585, new_AGEMA_signal_12584, mcs1_mcs_mat1_6_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_14035, new_AGEMA_signal_14034, new_AGEMA_signal_14033, mcs1_mcs_mat1_6_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_11224, new_AGEMA_signal_11223, new_AGEMA_signal_11222, mcs1_mcs_mat1_6_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_9967, new_AGEMA_signal_9966, new_AGEMA_signal_9965, mcs1_mcs_mat1_6_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_12586, new_AGEMA_signal_12585, new_AGEMA_signal_12584, mcs1_mcs_mat1_6_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_14038, new_AGEMA_signal_14037, new_AGEMA_signal_14036, mcs1_mcs_mat1_6_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_15463, new_AGEMA_signal_15462, new_AGEMA_signal_15461, mcs1_mcs_mat1_6_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_12592, new_AGEMA_signal_12591, new_AGEMA_signal_12590, mcs1_mcs_mat1_6_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_9967, new_AGEMA_signal_9966, new_AGEMA_signal_9965, mcs1_mcs_mat1_6_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_14038, new_AGEMA_signal_14037, new_AGEMA_signal_14036, mcs1_mcs_mat1_6_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_15466, new_AGEMA_signal_15465, new_AGEMA_signal_15464, mcs1_mcs_mat1_6_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .c ({new_AGEMA_signal_16477, new_AGEMA_signal_16476, new_AGEMA_signal_16475, mcs1_mcs_mat1_6_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_12592, new_AGEMA_signal_12591, new_AGEMA_signal_12590, mcs1_mcs_mat1_6_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_14041, new_AGEMA_signal_14040, new_AGEMA_signal_14039, mcs1_mcs_mat1_6_mcs_out[24]}), .c ({new_AGEMA_signal_15466, new_AGEMA_signal_15465, new_AGEMA_signal_15464, mcs1_mcs_mat1_6_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_12589, new_AGEMA_signal_12588, new_AGEMA_signal_12587, mcs1_mcs_mat1_6_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .c ({new_AGEMA_signal_14041, new_AGEMA_signal_14040, new_AGEMA_signal_14039, mcs1_mcs_mat1_6_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_11224, new_AGEMA_signal_11223, new_AGEMA_signal_11222, mcs1_mcs_mat1_6_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_9064, new_AGEMA_signal_9063, new_AGEMA_signal_9062, mcs1_mcs_mat1_6_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_12589, new_AGEMA_signal_12588, new_AGEMA_signal_12587, mcs1_mcs_mat1_6_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6095], Fresh[6094], Fresh[6093], Fresh[6092], Fresh[6091], Fresh[6090]}), .c ({new_AGEMA_signal_12592, new_AGEMA_signal_12591, new_AGEMA_signal_12590, mcs1_mcs_mat1_6_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6101], Fresh[6100], Fresh[6099], Fresh[6098], Fresh[6097], Fresh[6096]}), .c ({new_AGEMA_signal_9967, new_AGEMA_signal_9966, new_AGEMA_signal_9965, mcs1_mcs_mat1_6_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6107], Fresh[6106], Fresh[6105], Fresh[6104], Fresh[6103], Fresh[6102]}), .c ({new_AGEMA_signal_11224, new_AGEMA_signal_11223, new_AGEMA_signal_11222, mcs1_mcs_mat1_6_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_17947, new_AGEMA_signal_17946, new_AGEMA_signal_17945, mcs1_mcs_mat1_6_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .c ({new_AGEMA_signal_18586, new_AGEMA_signal_18585, new_AGEMA_signal_18584, mcs1_mcs_mat1_6_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_17275, new_AGEMA_signal_17274, new_AGEMA_signal_17273, mcs1_mcs_mat1_6_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_15469, new_AGEMA_signal_15468, new_AGEMA_signal_15467, mcs1_mcs_mat1_6_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_17947, new_AGEMA_signal_17946, new_AGEMA_signal_17945, mcs1_mcs_mat1_6_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_18589, new_AGEMA_signal_18588, new_AGEMA_signal_18587, mcs1_mcs_mat1_6_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .c ({new_AGEMA_signal_19252, new_AGEMA_signal_19251, new_AGEMA_signal_19250, mcs1_mcs_mat1_6_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_17953, new_AGEMA_signal_17952, new_AGEMA_signal_17951, mcs1_mcs_mat1_6_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_15469, new_AGEMA_signal_15468, new_AGEMA_signal_15467, mcs1_mcs_mat1_6_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_18589, new_AGEMA_signal_18588, new_AGEMA_signal_18587, mcs1_mcs_mat1_6_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_19255, new_AGEMA_signal_19254, new_AGEMA_signal_19253, mcs1_mcs_mat1_6_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_11392, new_AGEMA_signal_11391, new_AGEMA_signal_11390, mcs1_mcs_mat1_6_mcs_out[86]}), .c ({new_AGEMA_signal_19966, new_AGEMA_signal_19965, new_AGEMA_signal_19964, mcs1_mcs_mat1_6_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_17953, new_AGEMA_signal_17952, new_AGEMA_signal_17951, mcs1_mcs_mat1_6_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_18592, new_AGEMA_signal_18591, new_AGEMA_signal_18590, mcs1_mcs_mat1_6_mcs_out[20]}), .c ({new_AGEMA_signal_19255, new_AGEMA_signal_19254, new_AGEMA_signal_19253, mcs1_mcs_mat1_6_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_17950, new_AGEMA_signal_17949, new_AGEMA_signal_17948, mcs1_mcs_mat1_6_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .c ({new_AGEMA_signal_18592, new_AGEMA_signal_18591, new_AGEMA_signal_18590, mcs1_mcs_mat1_6_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_17275, new_AGEMA_signal_17274, new_AGEMA_signal_17273, mcs1_mcs_mat1_6_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_14044, new_AGEMA_signal_14043, new_AGEMA_signal_14042, mcs1_mcs_mat1_6_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_17950, new_AGEMA_signal_17949, new_AGEMA_signal_17948, mcs1_mcs_mat1_6_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6113], Fresh[6112], Fresh[6111], Fresh[6110], Fresh[6109], Fresh[6108]}), .c ({new_AGEMA_signal_17953, new_AGEMA_signal_17952, new_AGEMA_signal_17951, mcs1_mcs_mat1_6_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6119], Fresh[6118], Fresh[6117], Fresh[6116], Fresh[6115], Fresh[6114]}), .c ({new_AGEMA_signal_15469, new_AGEMA_signal_15468, new_AGEMA_signal_15467, mcs1_mcs_mat1_6_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6125], Fresh[6124], Fresh[6123], Fresh[6122], Fresh[6121], Fresh[6120]}), .c ({new_AGEMA_signal_17275, new_AGEMA_signal_17274, new_AGEMA_signal_17273, mcs1_mcs_mat1_6_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_12595, new_AGEMA_signal_12594, new_AGEMA_signal_12593, mcs1_mcs_mat1_6_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_12604, new_AGEMA_signal_12603, new_AGEMA_signal_12602, mcs1_mcs_mat1_6_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_14047, new_AGEMA_signal_14046, new_AGEMA_signal_14045, mcs1_mcs_mat1_6_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_14050, new_AGEMA_signal_14049, new_AGEMA_signal_14048, mcs1_mcs_mat1_6_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_9067, new_AGEMA_signal_9066, new_AGEMA_signal_9065, mcs1_mcs_mat1_6_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_15472, new_AGEMA_signal_15471, new_AGEMA_signal_15470, mcs1_mcs_mat1_6_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_15475, new_AGEMA_signal_15474, new_AGEMA_signal_15473, mcs1_mcs_mat1_6_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_9970, new_AGEMA_signal_9969, new_AGEMA_signal_9968, mcs1_mcs_mat1_6_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_16480, new_AGEMA_signal_16479, new_AGEMA_signal_16478, mcs1_mcs_mat1_6_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_8419, new_AGEMA_signal_8418, new_AGEMA_signal_8417, mcs1_mcs_mat1_6_mcs_out[50]}), .b ({new_AGEMA_signal_14050, new_AGEMA_signal_14049, new_AGEMA_signal_14048, mcs1_mcs_mat1_6_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_15475, new_AGEMA_signal_15474, new_AGEMA_signal_15473, mcs1_mcs_mat1_6_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_12598, new_AGEMA_signal_12597, new_AGEMA_signal_12596, mcs1_mcs_mat1_6_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .c ({new_AGEMA_signal_14050, new_AGEMA_signal_14049, new_AGEMA_signal_14048, mcs1_mcs_mat1_6_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_11227, new_AGEMA_signal_11226, new_AGEMA_signal_11225, mcs1_mcs_mat1_6_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_11230, new_AGEMA_signal_11229, new_AGEMA_signal_11228, mcs1_mcs_mat1_6_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_12598, new_AGEMA_signal_12597, new_AGEMA_signal_12596, mcs1_mcs_mat1_6_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_12601, new_AGEMA_signal_12600, new_AGEMA_signal_12599, mcs1_mcs_mat1_6_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_9970, new_AGEMA_signal_9969, new_AGEMA_signal_9968, mcs1_mcs_mat1_6_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_14053, new_AGEMA_signal_14052, new_AGEMA_signal_14051, mcs1_mcs_mat1_6_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6131], Fresh[6130], Fresh[6129], Fresh[6128], Fresh[6127], Fresh[6126]}), .c ({new_AGEMA_signal_12604, new_AGEMA_signal_12603, new_AGEMA_signal_12602, mcs1_mcs_mat1_6_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6137], Fresh[6136], Fresh[6135], Fresh[6134], Fresh[6133], Fresh[6132]}), .c ({new_AGEMA_signal_9970, new_AGEMA_signal_9969, new_AGEMA_signal_9968, mcs1_mcs_mat1_6_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6143], Fresh[6142], Fresh[6141], Fresh[6140], Fresh[6139], Fresh[6138]}), .c ({new_AGEMA_signal_11230, new_AGEMA_signal_11229, new_AGEMA_signal_11228, mcs1_mcs_mat1_6_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_15484, new_AGEMA_signal_15483, new_AGEMA_signal_15482, mcs1_mcs_mat1_6_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_10351, new_AGEMA_signal_10350, new_AGEMA_signal_10349, mcs1_mcs_mat1_6_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_16483, new_AGEMA_signal_16482, new_AGEMA_signal_16481, mcs1_mcs_mat1_6_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_14062, new_AGEMA_signal_14061, new_AGEMA_signal_14060, mcs1_mcs_mat1_6_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_14056, new_AGEMA_signal_14055, new_AGEMA_signal_14054, mcs1_mcs_mat1_6_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_15478, new_AGEMA_signal_15477, new_AGEMA_signal_15476, mcs1_mcs_mat1_6_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_12610, new_AGEMA_signal_12609, new_AGEMA_signal_12608, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_9973, new_AGEMA_signal_9972, new_AGEMA_signal_9971, mcs1_mcs_mat1_6_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_14056, new_AGEMA_signal_14055, new_AGEMA_signal_14054, mcs1_mcs_mat1_6_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_10351, new_AGEMA_signal_10350, new_AGEMA_signal_10349, mcs1_mcs_mat1_6_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_14059, new_AGEMA_signal_14058, new_AGEMA_signal_14057, mcs1_mcs_mat1_6_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_15481, new_AGEMA_signal_15480, new_AGEMA_signal_15479, mcs1_mcs_mat1_6_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_12607, new_AGEMA_signal_12606, new_AGEMA_signal_12605, mcs1_mcs_mat1_6_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_12610, new_AGEMA_signal_12609, new_AGEMA_signal_12608, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_14059, new_AGEMA_signal_14058, new_AGEMA_signal_14057, mcs1_mcs_mat1_6_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_9070, new_AGEMA_signal_9069, new_AGEMA_signal_9068, mcs1_mcs_mat1_6_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_9973, new_AGEMA_signal_9972, new_AGEMA_signal_9971, mcs1_mcs_mat1_6_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_10351, new_AGEMA_signal_10350, new_AGEMA_signal_10349, mcs1_mcs_mat1_6_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_16486, new_AGEMA_signal_16485, new_AGEMA_signal_16484, mcs1_mcs_mat1_6_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .c ({new_AGEMA_signal_17278, new_AGEMA_signal_17277, new_AGEMA_signal_17276, mcs1_mcs_mat1_6_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_15484, new_AGEMA_signal_15483, new_AGEMA_signal_15482, mcs1_mcs_mat1_6_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_12610, new_AGEMA_signal_12609, new_AGEMA_signal_12608, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_16486, new_AGEMA_signal_16485, new_AGEMA_signal_16484, mcs1_mcs_mat1_6_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({new_AGEMA_signal_14062, new_AGEMA_signal_14061, new_AGEMA_signal_14060, mcs1_mcs_mat1_6_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_15484, new_AGEMA_signal_15483, new_AGEMA_signal_15482, mcs1_mcs_mat1_6_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({new_AGEMA_signal_12607, new_AGEMA_signal_12606, new_AGEMA_signal_12605, mcs1_mcs_mat1_6_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_14062, new_AGEMA_signal_14061, new_AGEMA_signal_14060, mcs1_mcs_mat1_6_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_8365, new_AGEMA_signal_8364, new_AGEMA_signal_8363, shiftr_out[100]}), .b ({new_AGEMA_signal_11233, new_AGEMA_signal_11232, new_AGEMA_signal_11231, mcs1_mcs_mat1_6_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_12607, new_AGEMA_signal_12606, new_AGEMA_signal_12605, mcs1_mcs_mat1_6_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10404, new_AGEMA_signal_10403, mcs1_mcs_mat1_6_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6149], Fresh[6148], Fresh[6147], Fresh[6146], Fresh[6145], Fresh[6144]}), .c ({new_AGEMA_signal_12610, new_AGEMA_signal_12609, new_AGEMA_signal_12608, mcs1_mcs_mat1_6_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8568, new_AGEMA_signal_8567, mcs1_mcs_mat1_6_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6155], Fresh[6154], Fresh[6153], Fresh[6152], Fresh[6151], Fresh[6150]}), .c ({new_AGEMA_signal_9973, new_AGEMA_signal_9972, new_AGEMA_signal_9971, mcs1_mcs_mat1_6_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10207, new_AGEMA_signal_10206, new_AGEMA_signal_10205, mcs1_mcs_mat1_6_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6161], Fresh[6160], Fresh[6159], Fresh[6158], Fresh[6157], Fresh[6156]}), .c ({new_AGEMA_signal_11233, new_AGEMA_signal_11232, new_AGEMA_signal_11231, mcs1_mcs_mat1_6_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, new_AGEMA_signal_10352, mcs1_mcs_mat1_6_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .c ({new_AGEMA_signal_11236, new_AGEMA_signal_11235, new_AGEMA_signal_11234, mcs1_mcs_mat1_6_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_14068, new_AGEMA_signal_14067, new_AGEMA_signal_14066, mcs1_mcs_mat1_6_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .c ({new_AGEMA_signal_15487, new_AGEMA_signal_15486, new_AGEMA_signal_15485, mcs1_mcs_mat1_6_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_12613, new_AGEMA_signal_12612, new_AGEMA_signal_12611, mcs1_mcs_mat1_6_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .c ({new_AGEMA_signal_14065, new_AGEMA_signal_14064, new_AGEMA_signal_14063, mcs1_mcs_mat1_6_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_11239, new_AGEMA_signal_11238, new_AGEMA_signal_11237, mcs1_mcs_mat1_6_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, new_AGEMA_signal_10352, mcs1_mcs_mat1_6_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_12613, new_AGEMA_signal_12612, new_AGEMA_signal_12611, mcs1_mcs_mat1_6_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_9073, new_AGEMA_signal_9072, new_AGEMA_signal_9071, mcs1_mcs_mat1_6_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_9976, new_AGEMA_signal_9975, new_AGEMA_signal_9974, mcs1_mcs_mat1_6_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_10354, new_AGEMA_signal_10353, new_AGEMA_signal_10352, mcs1_mcs_mat1_6_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_15490, new_AGEMA_signal_15489, new_AGEMA_signal_15488, mcs1_mcs_mat1_6_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_8380, new_AGEMA_signal_8379, new_AGEMA_signal_8378, shiftr_out[68]}), .c ({new_AGEMA_signal_16489, new_AGEMA_signal_16488, new_AGEMA_signal_16487, mcs1_mcs_mat1_6_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_9073, new_AGEMA_signal_9072, new_AGEMA_signal_9071, mcs1_mcs_mat1_6_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_14068, new_AGEMA_signal_14067, new_AGEMA_signal_14066, mcs1_mcs_mat1_6_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_15490, new_AGEMA_signal_15489, new_AGEMA_signal_15488, mcs1_mcs_mat1_6_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_12616, new_AGEMA_signal_12615, new_AGEMA_signal_12614, mcs1_mcs_mat1_6_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_11239, new_AGEMA_signal_11238, new_AGEMA_signal_11237, mcs1_mcs_mat1_6_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_14068, new_AGEMA_signal_14067, new_AGEMA_signal_14066, mcs1_mcs_mat1_6_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10420, new_AGEMA_signal_10419, new_AGEMA_signal_10418, mcs1_mcs_mat1_6_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6167], Fresh[6166], Fresh[6165], Fresh[6164], Fresh[6163], Fresh[6162]}), .c ({new_AGEMA_signal_12616, new_AGEMA_signal_12615, new_AGEMA_signal_12614, mcs1_mcs_mat1_6_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8584, new_AGEMA_signal_8583, new_AGEMA_signal_8582, mcs1_mcs_mat1_6_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6173], Fresh[6172], Fresh[6171], Fresh[6170], Fresh[6169], Fresh[6168]}), .c ({new_AGEMA_signal_9976, new_AGEMA_signal_9975, new_AGEMA_signal_9974, mcs1_mcs_mat1_6_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10222, new_AGEMA_signal_10221, new_AGEMA_signal_10220, shiftr_out[71]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6179], Fresh[6178], Fresh[6177], Fresh[6176], Fresh[6175], Fresh[6174]}), .c ({new_AGEMA_signal_11239, new_AGEMA_signal_11238, new_AGEMA_signal_11237, mcs1_mcs_mat1_6_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_20722, new_AGEMA_signal_20721, new_AGEMA_signal_20720, mcs1_mcs_mat1_6_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_17284, new_AGEMA_signal_17283, new_AGEMA_signal_17282, mcs1_mcs_mat1_6_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_21328, new_AGEMA_signal_21327, new_AGEMA_signal_21326, mcs1_mcs_mat1_6_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_19969, new_AGEMA_signal_19968, new_AGEMA_signal_19967, mcs1_mcs_mat1_6_mcs_out[7]}), .b ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .c ({new_AGEMA_signal_20722, new_AGEMA_signal_20721, new_AGEMA_signal_20720, mcs1_mcs_mat1_6_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_19258, new_AGEMA_signal_19257, new_AGEMA_signal_19256, mcs1_mcs_mat1_6_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .c ({new_AGEMA_signal_19969, new_AGEMA_signal_19968, new_AGEMA_signal_19967, mcs1_mcs_mat1_6_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_18595, new_AGEMA_signal_18594, new_AGEMA_signal_18593, mcs1_mcs_mat1_6_mcs_out[6]}), .b ({new_AGEMA_signal_15496, new_AGEMA_signal_15495, new_AGEMA_signal_15494, mcs1_mcs_mat1_6_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_19258, new_AGEMA_signal_19257, new_AGEMA_signal_19256, mcs1_mcs_mat1_6_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_15493, new_AGEMA_signal_15492, new_AGEMA_signal_15491, mcs1_mcs_mat1_6_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_17956, new_AGEMA_signal_17955, new_AGEMA_signal_17954, mcs1_mcs_mat1_6_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_18595, new_AGEMA_signal_18594, new_AGEMA_signal_18593, mcs1_mcs_mat1_6_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16618, new_AGEMA_signal_16617, new_AGEMA_signal_16616, shiftr_out[37]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6185], Fresh[6184], Fresh[6183], Fresh[6182], Fresh[6181], Fresh[6180]}), .c ({new_AGEMA_signal_17956, new_AGEMA_signal_17955, new_AGEMA_signal_17954, mcs1_mcs_mat1_6_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12832, new_AGEMA_signal_12831, new_AGEMA_signal_12830, shiftr_out[38]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6191], Fresh[6190], Fresh[6189], Fresh[6188], Fresh[6187], Fresh[6186]}), .c ({new_AGEMA_signal_15496, new_AGEMA_signal_15495, new_AGEMA_signal_15494, mcs1_mcs_mat1_6_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15706, new_AGEMA_signal_15705, new_AGEMA_signal_15704, mcs1_mcs_mat1_6_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6197], Fresh[6196], Fresh[6195], Fresh[6194], Fresh[6193], Fresh[6192]}), .c ({new_AGEMA_signal_17284, new_AGEMA_signal_17283, new_AGEMA_signal_17282, mcs1_mcs_mat1_6_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_11242, new_AGEMA_signal_11241, new_AGEMA_signal_11240, mcs1_mcs_mat1_6_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_12619, new_AGEMA_signal_12618, new_AGEMA_signal_12617, mcs1_mcs_mat1_6_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_14077, new_AGEMA_signal_14076, new_AGEMA_signal_14075, mcs1_mcs_mat1_6_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .b ({new_AGEMA_signal_11245, new_AGEMA_signal_11244, new_AGEMA_signal_11243, mcs1_mcs_mat1_6_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_12619, new_AGEMA_signal_12618, new_AGEMA_signal_12617, mcs1_mcs_mat1_6_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_14080, new_AGEMA_signal_14079, new_AGEMA_signal_14078, mcs1_mcs_mat1_6_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_9979, new_AGEMA_signal_9978, new_AGEMA_signal_9977, mcs1_mcs_mat1_6_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_15499, new_AGEMA_signal_15498, new_AGEMA_signal_15497, mcs1_mcs_mat1_6_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_14083, new_AGEMA_signal_14082, new_AGEMA_signal_14081, mcs1_mcs_mat1_6_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_12625, new_AGEMA_signal_12624, new_AGEMA_signal_12623, mcs1_mcs_mat1_6_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_15502, new_AGEMA_signal_15501, new_AGEMA_signal_15500, mcs1_mcs_mat1_6_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_12628, new_AGEMA_signal_12627, new_AGEMA_signal_12626, mcs1_mcs_mat1_6_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_9076, new_AGEMA_signal_9075, new_AGEMA_signal_9074, mcs1_mcs_mat1_6_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_14083, new_AGEMA_signal_14082, new_AGEMA_signal_14081, mcs1_mcs_mat1_6_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10459, new_AGEMA_signal_10458, new_AGEMA_signal_10457, shiftr_out[5]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6203], Fresh[6202], Fresh[6201], Fresh[6200], Fresh[6199], Fresh[6198]}), .c ({new_AGEMA_signal_12628, new_AGEMA_signal_12627, new_AGEMA_signal_12626, mcs1_mcs_mat1_6_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8623, new_AGEMA_signal_8622, new_AGEMA_signal_8621, shiftr_out[6]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6209], Fresh[6208], Fresh[6207], Fresh[6206], Fresh[6205], Fresh[6204]}), .c ({new_AGEMA_signal_9979, new_AGEMA_signal_9978, new_AGEMA_signal_9977, mcs1_mcs_mat1_6_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_6_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10260, new_AGEMA_signal_10259, mcs1_mcs_mat1_6_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6215], Fresh[6214], Fresh[6213], Fresh[6212], Fresh[6211], Fresh[6210]}), .c ({new_AGEMA_signal_11245, new_AGEMA_signal_11244, new_AGEMA_signal_11243, mcs1_mcs_mat1_6_mcs_rom0_31_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U96 ( .a ({new_AGEMA_signal_17287, new_AGEMA_signal_17286, new_AGEMA_signal_17285, mcs1_mcs_mat1_7_n128}), .b ({new_AGEMA_signal_19972, new_AGEMA_signal_19971, new_AGEMA_signal_19970, mcs1_mcs_mat1_7_n127}), .c ({temp_next_s3[65], temp_next_s2[65], temp_next_s1[65], temp_next_s0[65]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U95 ( .a ({new_AGEMA_signal_19327, new_AGEMA_signal_19326, new_AGEMA_signal_19325, mcs1_mcs_mat1_7_mcs_out[41]}), .b ({new_AGEMA_signal_12736, new_AGEMA_signal_12735, new_AGEMA_signal_12734, mcs1_mcs_mat1_7_mcs_out[45]}), .c ({new_AGEMA_signal_19972, new_AGEMA_signal_19971, new_AGEMA_signal_19970, mcs1_mcs_mat1_7_n127}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U94 ( .a ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, new_AGEMA_signal_10358, mcs1_mcs_mat1_7_mcs_out[33]}), .b ({new_AGEMA_signal_16570, new_AGEMA_signal_16569, new_AGEMA_signal_16568, mcs1_mcs_mat1_7_mcs_out[37]}), .c ({new_AGEMA_signal_17287, new_AGEMA_signal_17286, new_AGEMA_signal_17285, mcs1_mcs_mat1_7_n128}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U93 ( .a ({new_AGEMA_signal_17959, new_AGEMA_signal_17958, new_AGEMA_signal_17957, mcs1_mcs_mat1_7_n126}), .b ({new_AGEMA_signal_19261, new_AGEMA_signal_19260, new_AGEMA_signal_19259, mcs1_mcs_mat1_7_n125}), .c ({temp_next_s3[64], temp_next_s2[64], temp_next_s1[64], temp_next_s0[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U92 ( .a ({new_AGEMA_signal_18658, new_AGEMA_signal_18657, new_AGEMA_signal_18656, mcs1_mcs_mat1_7_mcs_out[40]}), .b ({new_AGEMA_signal_17365, new_AGEMA_signal_17364, new_AGEMA_signal_17363, mcs1_mcs_mat1_7_mcs_out[44]}), .c ({new_AGEMA_signal_19261, new_AGEMA_signal_19260, new_AGEMA_signal_19259, mcs1_mcs_mat1_7_n125}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U91 ( .a ({new_AGEMA_signal_17374, new_AGEMA_signal_17373, new_AGEMA_signal_17372, mcs1_mcs_mat1_7_mcs_out[32]}), .b ({new_AGEMA_signal_14188, new_AGEMA_signal_14187, new_AGEMA_signal_14186, mcs1_mcs_mat1_7_mcs_out[36]}), .c ({new_AGEMA_signal_17959, new_AGEMA_signal_17958, new_AGEMA_signal_17957, mcs1_mcs_mat1_7_n126}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U90 ( .a ({new_AGEMA_signal_15505, new_AGEMA_signal_15504, new_AGEMA_signal_15503, mcs1_mcs_mat1_7_n124}), .b ({new_AGEMA_signal_19264, new_AGEMA_signal_19263, new_AGEMA_signal_19262, mcs1_mcs_mat1_7_n123}), .c ({temp_next_s3[35], temp_next_s2[35], temp_next_s1[35], temp_next_s0[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U89 ( .a ({new_AGEMA_signal_18661, new_AGEMA_signal_18660, new_AGEMA_signal_18659, mcs1_mcs_mat1_7_mcs_out[27]}), .b ({new_AGEMA_signal_16576, new_AGEMA_signal_16575, new_AGEMA_signal_16574, mcs1_mcs_mat1_7_mcs_out[31]}), .c ({new_AGEMA_signal_19264, new_AGEMA_signal_19263, new_AGEMA_signal_19262, mcs1_mcs_mat1_7_n123}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U88 ( .a ({new_AGEMA_signal_14218, new_AGEMA_signal_14217, new_AGEMA_signal_14216, mcs1_mcs_mat1_7_mcs_out[19]}), .b ({new_AGEMA_signal_14209, new_AGEMA_signal_14208, new_AGEMA_signal_14207, mcs1_mcs_mat1_7_mcs_out[23]}), .c ({new_AGEMA_signal_15505, new_AGEMA_signal_15504, new_AGEMA_signal_15503, mcs1_mcs_mat1_7_n124}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U87 ( .a ({new_AGEMA_signal_16492, new_AGEMA_signal_16491, new_AGEMA_signal_16490, mcs1_mcs_mat1_7_n122}), .b ({new_AGEMA_signal_19981, new_AGEMA_signal_19980, new_AGEMA_signal_19979, mcs1_mcs_mat1_7_n121}), .c ({temp_next_s3[34], temp_next_s2[34], temp_next_s1[34], temp_next_s0[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U86 ( .a ({new_AGEMA_signal_19330, new_AGEMA_signal_19329, new_AGEMA_signal_19328, mcs1_mcs_mat1_7_mcs_out[26]}), .b ({new_AGEMA_signal_15640, new_AGEMA_signal_15639, new_AGEMA_signal_15638, mcs1_mcs_mat1_7_mcs_out[30]}), .c ({new_AGEMA_signal_19981, new_AGEMA_signal_19980, new_AGEMA_signal_19979, mcs1_mcs_mat1_7_n121}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U85 ( .a ({new_AGEMA_signal_15655, new_AGEMA_signal_15654, new_AGEMA_signal_15653, mcs1_mcs_mat1_7_mcs_out[18]}), .b ({new_AGEMA_signal_15649, new_AGEMA_signal_15648, new_AGEMA_signal_15647, mcs1_mcs_mat1_7_mcs_out[22]}), .c ({new_AGEMA_signal_16492, new_AGEMA_signal_16491, new_AGEMA_signal_16490, mcs1_mcs_mat1_7_n122}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U84 ( .a ({new_AGEMA_signal_17290, new_AGEMA_signal_17289, new_AGEMA_signal_17288, mcs1_mcs_mat1_7_n120}), .b ({new_AGEMA_signal_20731, new_AGEMA_signal_20730, new_AGEMA_signal_20729, mcs1_mcs_mat1_7_n119}), .c ({temp_next_s3[33], temp_next_s2[33], temp_next_s1[33], temp_next_s0[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U83 ( .a ({new_AGEMA_signal_20038, new_AGEMA_signal_20037, new_AGEMA_signal_20036, mcs1_mcs_mat1_7_mcs_out[25]}), .b ({new_AGEMA_signal_14200, new_AGEMA_signal_14199, new_AGEMA_signal_14198, mcs1_mcs_mat1_7_mcs_out[29]}), .c ({new_AGEMA_signal_20731, new_AGEMA_signal_20730, new_AGEMA_signal_20729, mcs1_mcs_mat1_7_n119}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U82 ( .a ({new_AGEMA_signal_16585, new_AGEMA_signal_16584, new_AGEMA_signal_16583, mcs1_mcs_mat1_7_mcs_out[17]}), .b ({new_AGEMA_signal_16582, new_AGEMA_signal_16581, new_AGEMA_signal_16580, mcs1_mcs_mat1_7_mcs_out[21]}), .c ({new_AGEMA_signal_17290, new_AGEMA_signal_17289, new_AGEMA_signal_17288, mcs1_mcs_mat1_7_n120}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U81 ( .a ({new_AGEMA_signal_15508, new_AGEMA_signal_15507, new_AGEMA_signal_15506, mcs1_mcs_mat1_7_n118}), .b ({new_AGEMA_signal_19267, new_AGEMA_signal_19266, new_AGEMA_signal_19265, mcs1_mcs_mat1_7_n117}), .c ({temp_next_s3[32], temp_next_s2[32], temp_next_s1[32], temp_next_s0[32]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U80 ( .a ({new_AGEMA_signal_18667, new_AGEMA_signal_18666, new_AGEMA_signal_18665, mcs1_mcs_mat1_7_mcs_out[24]}), .b ({new_AGEMA_signal_16579, new_AGEMA_signal_16578, new_AGEMA_signal_16577, mcs1_mcs_mat1_7_mcs_out[28]}), .c ({new_AGEMA_signal_19267, new_AGEMA_signal_19266, new_AGEMA_signal_19265, mcs1_mcs_mat1_7_n117}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U79 ( .a ({new_AGEMA_signal_14224, new_AGEMA_signal_14223, new_AGEMA_signal_14222, mcs1_mcs_mat1_7_mcs_out[16]}), .b ({new_AGEMA_signal_14215, new_AGEMA_signal_14214, new_AGEMA_signal_14213, mcs1_mcs_mat1_7_mcs_out[20]}), .c ({new_AGEMA_signal_15508, new_AGEMA_signal_15507, new_AGEMA_signal_15506, mcs1_mcs_mat1_7_n118}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U78 ( .a ({new_AGEMA_signal_17962, new_AGEMA_signal_17961, new_AGEMA_signal_17960, mcs1_mcs_mat1_7_n116}), .b ({new_AGEMA_signal_17293, new_AGEMA_signal_17292, new_AGEMA_signal_17291, mcs1_mcs_mat1_7_n115}), .c ({temp_next_s3[3], temp_next_s2[3], temp_next_s1[3], temp_next_s0[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U77 ( .a ({new_AGEMA_signal_14242, new_AGEMA_signal_14241, new_AGEMA_signal_14240, mcs1_mcs_mat1_7_mcs_out[3]}), .b ({new_AGEMA_signal_16597, new_AGEMA_signal_16596, new_AGEMA_signal_16595, mcs1_mcs_mat1_7_mcs_out[7]}), .c ({new_AGEMA_signal_17293, new_AGEMA_signal_17292, new_AGEMA_signal_17291, mcs1_mcs_mat1_7_n115}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U76 ( .a ({new_AGEMA_signal_17383, new_AGEMA_signal_17382, new_AGEMA_signal_17381, mcs1_mcs_mat1_7_mcs_out[11]}), .b ({new_AGEMA_signal_16588, new_AGEMA_signal_16587, new_AGEMA_signal_16586, mcs1_mcs_mat1_7_mcs_out[15]}), .c ({new_AGEMA_signal_17962, new_AGEMA_signal_17961, new_AGEMA_signal_17960, mcs1_mcs_mat1_7_n116}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U75 ( .a ({new_AGEMA_signal_17296, new_AGEMA_signal_17295, new_AGEMA_signal_17294, mcs1_mcs_mat1_7_n114}), .b ({new_AGEMA_signal_20734, new_AGEMA_signal_20733, new_AGEMA_signal_20732, mcs1_mcs_mat1_7_n113}), .c ({new_AGEMA_signal_21334, new_AGEMA_signal_21333, new_AGEMA_signal_21332, mcs_out[227]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U74 ( .a ({new_AGEMA_signal_20023, new_AGEMA_signal_20022, new_AGEMA_signal_20021, mcs1_mcs_mat1_7_mcs_out[123]}), .b ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_20734, new_AGEMA_signal_20733, new_AGEMA_signal_20732, mcs1_mcs_mat1_7_n113}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U73 ( .a ({new_AGEMA_signal_15541, new_AGEMA_signal_15540, new_AGEMA_signal_15539, mcs1_mcs_mat1_7_mcs_out[115]}), .b ({new_AGEMA_signal_16510, new_AGEMA_signal_16509, new_AGEMA_signal_16508, mcs1_mcs_mat1_7_mcs_out[119]}), .c ({new_AGEMA_signal_17296, new_AGEMA_signal_17295, new_AGEMA_signal_17294, mcs1_mcs_mat1_7_n114}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U72 ( .a ({new_AGEMA_signal_17299, new_AGEMA_signal_17298, new_AGEMA_signal_17297, mcs1_mcs_mat1_7_n112}), .b ({new_AGEMA_signal_18601, new_AGEMA_signal_18600, new_AGEMA_signal_18599, mcs1_mcs_mat1_7_n111}), .c ({new_AGEMA_signal_19270, new_AGEMA_signal_19269, new_AGEMA_signal_19268, mcs_out[226]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U71 ( .a ({new_AGEMA_signal_17983, new_AGEMA_signal_17982, new_AGEMA_signal_17981, mcs1_mcs_mat1_7_mcs_out[122]}), .b ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_18601, new_AGEMA_signal_18600, new_AGEMA_signal_18599, mcs1_mcs_mat1_7_n111}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U70 ( .a ({new_AGEMA_signal_14095, new_AGEMA_signal_14094, new_AGEMA_signal_14093, mcs1_mcs_mat1_7_mcs_out[114]}), .b ({new_AGEMA_signal_16513, new_AGEMA_signal_16512, new_AGEMA_signal_16511, mcs1_mcs_mat1_7_mcs_out[118]}), .c ({new_AGEMA_signal_17299, new_AGEMA_signal_17298, new_AGEMA_signal_17297, mcs1_mcs_mat1_7_n112}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U69 ( .a ({new_AGEMA_signal_19987, new_AGEMA_signal_19986, new_AGEMA_signal_19985, mcs1_mcs_mat1_7_n110}), .b ({new_AGEMA_signal_15511, new_AGEMA_signal_15510, new_AGEMA_signal_15509, mcs1_mcs_mat1_7_n109}), .c ({temp_next_s3[2], temp_next_s2[2], temp_next_s1[2], temp_next_s0[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U68 ( .a ({new_AGEMA_signal_14245, new_AGEMA_signal_14244, new_AGEMA_signal_14243, mcs1_mcs_mat1_7_mcs_out[2]}), .b ({new_AGEMA_signal_14239, new_AGEMA_signal_14238, new_AGEMA_signal_14237, mcs1_mcs_mat1_7_mcs_out[6]}), .c ({new_AGEMA_signal_15511, new_AGEMA_signal_15510, new_AGEMA_signal_15509, mcs1_mcs_mat1_7_n109}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U67 ( .a ({new_AGEMA_signal_19336, new_AGEMA_signal_19335, new_AGEMA_signal_19334, mcs1_mcs_mat1_7_mcs_out[10]}), .b ({new_AGEMA_signal_15661, new_AGEMA_signal_15660, new_AGEMA_signal_15659, mcs1_mcs_mat1_7_mcs_out[14]}), .c ({new_AGEMA_signal_19987, new_AGEMA_signal_19986, new_AGEMA_signal_19985, mcs1_mcs_mat1_7_n110}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U66 ( .a ({new_AGEMA_signal_16495, new_AGEMA_signal_16494, new_AGEMA_signal_16493, mcs1_mcs_mat1_7_n108}), .b ({new_AGEMA_signal_20740, new_AGEMA_signal_20739, new_AGEMA_signal_20738, mcs1_mcs_mat1_7_n107}), .c ({new_AGEMA_signal_21337, new_AGEMA_signal_21336, new_AGEMA_signal_21335, mcs_out[225]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U65 ( .a ({new_AGEMA_signal_20026, new_AGEMA_signal_20025, new_AGEMA_signal_20024, mcs1_mcs_mat1_7_mcs_out[121]}), .b ({new_AGEMA_signal_11248, new_AGEMA_signal_11247, new_AGEMA_signal_11246, mcs1_mcs_mat1_7_mcs_out[125]}), .c ({new_AGEMA_signal_20740, new_AGEMA_signal_20739, new_AGEMA_signal_20738, mcs1_mcs_mat1_7_n107}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U64 ( .a ({new_AGEMA_signal_12640, new_AGEMA_signal_12639, new_AGEMA_signal_12638, mcs1_mcs_mat1_7_mcs_out[113]}), .b ({new_AGEMA_signal_15538, new_AGEMA_signal_15537, new_AGEMA_signal_15536, mcs1_mcs_mat1_7_mcs_out[117]}), .c ({new_AGEMA_signal_16495, new_AGEMA_signal_16494, new_AGEMA_signal_16493, mcs1_mcs_mat1_7_n108}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U63 ( .a ({new_AGEMA_signal_17302, new_AGEMA_signal_17301, new_AGEMA_signal_17300, mcs1_mcs_mat1_7_n106}), .b ({new_AGEMA_signal_19990, new_AGEMA_signal_19989, new_AGEMA_signal_19988, mcs1_mcs_mat1_7_n105}), .c ({new_AGEMA_signal_20743, new_AGEMA_signal_20742, new_AGEMA_signal_20741, mcs_out[224]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U62 ( .a ({new_AGEMA_signal_19297, new_AGEMA_signal_19296, new_AGEMA_signal_19295, mcs1_mcs_mat1_7_mcs_out[120]}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_19990, new_AGEMA_signal_19989, new_AGEMA_signal_19988, mcs1_mcs_mat1_7_n105}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U61 ( .a ({new_AGEMA_signal_16516, new_AGEMA_signal_16515, new_AGEMA_signal_16514, mcs1_mcs_mat1_7_mcs_out[112]}), .b ({new_AGEMA_signal_14092, new_AGEMA_signal_14091, new_AGEMA_signal_14090, mcs1_mcs_mat1_7_mcs_out[116]}), .c ({new_AGEMA_signal_17302, new_AGEMA_signal_17301, new_AGEMA_signal_17300, mcs1_mcs_mat1_7_n106}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U60 ( .a ({new_AGEMA_signal_19993, new_AGEMA_signal_19992, new_AGEMA_signal_19991, mcs1_mcs_mat1_7_n104}), .b ({new_AGEMA_signal_17305, new_AGEMA_signal_17304, new_AGEMA_signal_17303, mcs1_mcs_mat1_7_n103}), .c ({new_AGEMA_signal_20746, new_AGEMA_signal_20745, new_AGEMA_signal_20744, mcs_out[195]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U59 ( .a ({new_AGEMA_signal_16519, new_AGEMA_signal_16518, new_AGEMA_signal_16517, mcs1_mcs_mat1_7_mcs_out[111]}), .b ({new_AGEMA_signal_16531, new_AGEMA_signal_16530, new_AGEMA_signal_16529, mcs1_mcs_mat1_7_mcs_out[99]}), .c ({new_AGEMA_signal_17305, new_AGEMA_signal_17304, new_AGEMA_signal_17303, mcs1_mcs_mat1_7_n103}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U58 ( .a ({new_AGEMA_signal_15556, new_AGEMA_signal_15555, new_AGEMA_signal_15554, mcs1_mcs_mat1_7_mcs_out[103]}), .b ({new_AGEMA_signal_19300, new_AGEMA_signal_19299, new_AGEMA_signal_19298, mcs1_mcs_mat1_7_mcs_out[107]}), .c ({new_AGEMA_signal_19993, new_AGEMA_signal_19992, new_AGEMA_signal_19991, mcs1_mcs_mat1_7_n104}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U57 ( .a ({new_AGEMA_signal_19996, new_AGEMA_signal_19995, new_AGEMA_signal_19994, mcs1_mcs_mat1_7_n102}), .b ({new_AGEMA_signal_17308, new_AGEMA_signal_17307, new_AGEMA_signal_17306, mcs1_mcs_mat1_7_n101}), .c ({new_AGEMA_signal_20749, new_AGEMA_signal_20748, new_AGEMA_signal_20747, mcs_out[194]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U56 ( .a ({new_AGEMA_signal_16522, new_AGEMA_signal_16521, new_AGEMA_signal_16520, mcs1_mcs_mat1_7_mcs_out[110]}), .b ({new_AGEMA_signal_14122, new_AGEMA_signal_14121, new_AGEMA_signal_14120, mcs1_mcs_mat1_7_mcs_out[98]}), .c ({new_AGEMA_signal_17308, new_AGEMA_signal_17307, new_AGEMA_signal_17306, mcs1_mcs_mat1_7_n101}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U55 ( .a ({new_AGEMA_signal_12655, new_AGEMA_signal_12654, new_AGEMA_signal_12653, mcs1_mcs_mat1_7_mcs_out[102]}), .b ({new_AGEMA_signal_19303, new_AGEMA_signal_19302, new_AGEMA_signal_19301, mcs1_mcs_mat1_7_mcs_out[106]}), .c ({new_AGEMA_signal_19996, new_AGEMA_signal_19995, new_AGEMA_signal_19994, mcs1_mcs_mat1_7_n102}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U54 ( .a ({new_AGEMA_signal_19999, new_AGEMA_signal_19998, new_AGEMA_signal_19997, mcs1_mcs_mat1_7_n100}), .b ({new_AGEMA_signal_17311, new_AGEMA_signal_17310, new_AGEMA_signal_17309, mcs1_mcs_mat1_7_n99}), .c ({new_AGEMA_signal_20752, new_AGEMA_signal_20751, new_AGEMA_signal_20750, mcs_out[193]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U53 ( .a ({new_AGEMA_signal_16525, new_AGEMA_signal_16524, new_AGEMA_signal_16523, mcs1_mcs_mat1_7_mcs_out[109]}), .b ({new_AGEMA_signal_11275, new_AGEMA_signal_11274, new_AGEMA_signal_11273, mcs1_mcs_mat1_7_mcs_out[97]}), .c ({new_AGEMA_signal_17311, new_AGEMA_signal_17310, new_AGEMA_signal_17309, mcs1_mcs_mat1_7_n99}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U52 ( .a ({new_AGEMA_signal_14116, new_AGEMA_signal_14115, new_AGEMA_signal_14114, mcs1_mcs_mat1_7_mcs_out[101]}), .b ({new_AGEMA_signal_19306, new_AGEMA_signal_19305, new_AGEMA_signal_19304, mcs1_mcs_mat1_7_mcs_out[105]}), .c ({new_AGEMA_signal_19999, new_AGEMA_signal_19998, new_AGEMA_signal_19997, mcs1_mcs_mat1_7_n100}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U51 ( .a ({new_AGEMA_signal_20755, new_AGEMA_signal_20754, new_AGEMA_signal_20753, mcs1_mcs_mat1_7_n98}), .b ({new_AGEMA_signal_18604, new_AGEMA_signal_18603, new_AGEMA_signal_18602, mcs1_mcs_mat1_7_n97}), .c ({new_AGEMA_signal_21340, new_AGEMA_signal_21339, new_AGEMA_signal_21338, mcs_out[192]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U50 ( .a ({new_AGEMA_signal_16528, new_AGEMA_signal_16527, new_AGEMA_signal_16526, mcs1_mcs_mat1_7_mcs_out[108]}), .b ({new_AGEMA_signal_17995, new_AGEMA_signal_17994, new_AGEMA_signal_17993, mcs1_mcs_mat1_7_mcs_out[96]}), .c ({new_AGEMA_signal_18604, new_AGEMA_signal_18603, new_AGEMA_signal_18602, mcs1_mcs_mat1_7_n97}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U49 ( .a ({new_AGEMA_signal_15559, new_AGEMA_signal_15558, new_AGEMA_signal_15557, mcs1_mcs_mat1_7_mcs_out[100]}), .b ({new_AGEMA_signal_20029, new_AGEMA_signal_20028, new_AGEMA_signal_20027, mcs1_mcs_mat1_7_mcs_out[104]}), .c ({new_AGEMA_signal_20755, new_AGEMA_signal_20754, new_AGEMA_signal_20753, mcs1_mcs_mat1_7_n98}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U48 ( .a ({new_AGEMA_signal_15514, new_AGEMA_signal_15513, new_AGEMA_signal_15512, mcs1_mcs_mat1_7_n96}), .b ({new_AGEMA_signal_17965, new_AGEMA_signal_17964, new_AGEMA_signal_17963, mcs1_mcs_mat1_7_n95}), .c ({new_AGEMA_signal_18607, new_AGEMA_signal_18606, new_AGEMA_signal_18605, mcs_out[163]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U47 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_15565, new_AGEMA_signal_15564, new_AGEMA_signal_15563, mcs1_mcs_mat1_7_mcs_out[95]}), .c ({new_AGEMA_signal_17965, new_AGEMA_signal_17964, new_AGEMA_signal_17963, mcs1_mcs_mat1_7_n95}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U46 ( .a ({new_AGEMA_signal_14131, new_AGEMA_signal_14130, new_AGEMA_signal_14129, mcs1_mcs_mat1_7_mcs_out[83]}), .b ({new_AGEMA_signal_12679, new_AGEMA_signal_12678, new_AGEMA_signal_12677, mcs1_mcs_mat1_7_mcs_out[87]}), .c ({new_AGEMA_signal_15514, new_AGEMA_signal_15513, new_AGEMA_signal_15512, mcs1_mcs_mat1_7_n96}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U45 ( .a ({new_AGEMA_signal_15517, new_AGEMA_signal_15516, new_AGEMA_signal_15515, mcs1_mcs_mat1_7_n94}), .b ({new_AGEMA_signal_17968, new_AGEMA_signal_17967, new_AGEMA_signal_17966, mcs1_mcs_mat1_7_n93}), .c ({new_AGEMA_signal_18610, new_AGEMA_signal_18609, new_AGEMA_signal_18608, mcs_out[162]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U43 ( .a ({new_AGEMA_signal_14134, new_AGEMA_signal_14133, new_AGEMA_signal_14132, mcs1_mcs_mat1_7_mcs_out[82]}), .b ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_15517, new_AGEMA_signal_15516, new_AGEMA_signal_15515, mcs1_mcs_mat1_7_n94}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U42 ( .a ({new_AGEMA_signal_15520, new_AGEMA_signal_15519, new_AGEMA_signal_15518, mcs1_mcs_mat1_7_n92}), .b ({new_AGEMA_signal_17971, new_AGEMA_signal_17970, new_AGEMA_signal_17969, mcs1_mcs_mat1_7_n91}), .c ({new_AGEMA_signal_18613, new_AGEMA_signal_18612, new_AGEMA_signal_18611, mcs_out[161]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U41 ( .a ({new_AGEMA_signal_17353, new_AGEMA_signal_17352, new_AGEMA_signal_17351, mcs1_mcs_mat1_7_mcs_out[89]}), .b ({new_AGEMA_signal_12673, new_AGEMA_signal_12672, new_AGEMA_signal_12671, mcs1_mcs_mat1_7_mcs_out[93]}), .c ({new_AGEMA_signal_17971, new_AGEMA_signal_17970, new_AGEMA_signal_17969, mcs1_mcs_mat1_7_n91}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U40 ( .a ({new_AGEMA_signal_14137, new_AGEMA_signal_14136, new_AGEMA_signal_14135, mcs1_mcs_mat1_7_mcs_out[81]}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_15520, new_AGEMA_signal_15519, new_AGEMA_signal_15518, mcs1_mcs_mat1_7_n92}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U39 ( .a ({new_AGEMA_signal_16498, new_AGEMA_signal_16497, new_AGEMA_signal_16496, mcs1_mcs_mat1_7_n90}), .b ({new_AGEMA_signal_17314, new_AGEMA_signal_17313, new_AGEMA_signal_17312, mcs1_mcs_mat1_7_n89}), .c ({new_AGEMA_signal_17974, new_AGEMA_signal_17973, new_AGEMA_signal_17972, mcs_out[160]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U38 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_16534, new_AGEMA_signal_16533, new_AGEMA_signal_16532, mcs1_mcs_mat1_7_mcs_out[92]}), .c ({new_AGEMA_signal_17314, new_AGEMA_signal_17313, new_AGEMA_signal_17312, mcs1_mcs_mat1_7_n89}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U37 ( .a ({new_AGEMA_signal_15571, new_AGEMA_signal_15570, new_AGEMA_signal_15569, mcs1_mcs_mat1_7_mcs_out[80]}), .b ({new_AGEMA_signal_14128, new_AGEMA_signal_14127, new_AGEMA_signal_14126, mcs1_mcs_mat1_7_mcs_out[84]}), .c ({new_AGEMA_signal_16498, new_AGEMA_signal_16497, new_AGEMA_signal_16496, mcs1_mcs_mat1_7_n90}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U36 ( .a ({new_AGEMA_signal_16501, new_AGEMA_signal_16500, new_AGEMA_signal_16499, mcs1_mcs_mat1_7_n88}), .b ({new_AGEMA_signal_19273, new_AGEMA_signal_19272, new_AGEMA_signal_19271, mcs1_mcs_mat1_7_n87}), .c ({temp_next_s3[1], temp_next_s2[1], temp_next_s1[1], temp_next_s0[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U35 ( .a ({new_AGEMA_signal_11344, new_AGEMA_signal_11343, new_AGEMA_signal_11342, mcs1_mcs_mat1_7_mcs_out[5]}), .b ({new_AGEMA_signal_18670, new_AGEMA_signal_18669, new_AGEMA_signal_18668, mcs1_mcs_mat1_7_mcs_out[9]}), .c ({new_AGEMA_signal_19273, new_AGEMA_signal_19272, new_AGEMA_signal_19271, mcs1_mcs_mat1_7_n87}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U34 ( .a ({new_AGEMA_signal_15664, new_AGEMA_signal_15663, new_AGEMA_signal_15662, mcs1_mcs_mat1_7_mcs_out[13]}), .b ({new_AGEMA_signal_15676, new_AGEMA_signal_15675, new_AGEMA_signal_15674, mcs1_mcs_mat1_7_mcs_out[1]}), .c ({new_AGEMA_signal_16501, new_AGEMA_signal_16500, new_AGEMA_signal_16499, mcs1_mcs_mat1_7_n88}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U33 ( .a ({new_AGEMA_signal_17317, new_AGEMA_signal_17316, new_AGEMA_signal_17315, mcs1_mcs_mat1_7_n86}), .b ({new_AGEMA_signal_18616, new_AGEMA_signal_18615, new_AGEMA_signal_18614, mcs1_mcs_mat1_7_n85}), .c ({new_AGEMA_signal_19276, new_AGEMA_signal_19275, new_AGEMA_signal_19274, mcs_out[131]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U32 ( .a ({new_AGEMA_signal_17998, new_AGEMA_signal_17997, new_AGEMA_signal_17996, mcs1_mcs_mat1_7_mcs_out[75]}), .b ({new_AGEMA_signal_15574, new_AGEMA_signal_15573, new_AGEMA_signal_15572, mcs1_mcs_mat1_7_mcs_out[79]}), .c ({new_AGEMA_signal_18616, new_AGEMA_signal_18615, new_AGEMA_signal_18614, mcs1_mcs_mat1_7_n85}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U31 ( .a ({new_AGEMA_signal_16549, new_AGEMA_signal_16548, new_AGEMA_signal_16547, mcs1_mcs_mat1_7_mcs_out[67]}), .b ({new_AGEMA_signal_15586, new_AGEMA_signal_15585, new_AGEMA_signal_15584, mcs1_mcs_mat1_7_mcs_out[71]}), .c ({new_AGEMA_signal_17317, new_AGEMA_signal_17316, new_AGEMA_signal_17315, mcs1_mcs_mat1_7_n86}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U30 ( .a ({new_AGEMA_signal_17320, new_AGEMA_signal_17319, new_AGEMA_signal_17318, mcs1_mcs_mat1_7_n84}), .b ({new_AGEMA_signal_20758, new_AGEMA_signal_20757, new_AGEMA_signal_20756, mcs1_mcs_mat1_7_n83}), .c ({new_AGEMA_signal_21343, new_AGEMA_signal_21342, new_AGEMA_signal_21341, mcs_out[130]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U29 ( .a ({new_AGEMA_signal_20032, new_AGEMA_signal_20031, new_AGEMA_signal_20030, mcs1_mcs_mat1_7_mcs_out[74]}), .b ({new_AGEMA_signal_10009, new_AGEMA_signal_10008, new_AGEMA_signal_10007, mcs1_mcs_mat1_7_mcs_out[78]}), .c ({new_AGEMA_signal_20758, new_AGEMA_signal_20757, new_AGEMA_signal_20756, mcs1_mcs_mat1_7_n83}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U28 ( .a ({new_AGEMA_signal_15595, new_AGEMA_signal_15594, new_AGEMA_signal_15593, mcs1_mcs_mat1_7_mcs_out[66]}), .b ({new_AGEMA_signal_16543, new_AGEMA_signal_16542, new_AGEMA_signal_16541, mcs1_mcs_mat1_7_mcs_out[70]}), .c ({new_AGEMA_signal_17320, new_AGEMA_signal_17319, new_AGEMA_signal_17318, mcs1_mcs_mat1_7_n84}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U27 ( .a ({new_AGEMA_signal_17323, new_AGEMA_signal_17322, new_AGEMA_signal_17321, mcs1_mcs_mat1_7_n82}), .b ({new_AGEMA_signal_19279, new_AGEMA_signal_19278, new_AGEMA_signal_19277, mcs1_mcs_mat1_7_n81}), .c ({new_AGEMA_signal_20005, new_AGEMA_signal_20004, new_AGEMA_signal_20003, mcs_out[129]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U26 ( .a ({new_AGEMA_signal_18634, new_AGEMA_signal_18633, new_AGEMA_signal_18632, mcs1_mcs_mat1_7_mcs_out[73]}), .b ({new_AGEMA_signal_12694, new_AGEMA_signal_12693, new_AGEMA_signal_12692, mcs1_mcs_mat1_7_mcs_out[77]}), .c ({new_AGEMA_signal_19279, new_AGEMA_signal_19278, new_AGEMA_signal_19277, mcs1_mcs_mat1_7_n81}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U25 ( .a ({new_AGEMA_signal_12709, new_AGEMA_signal_12708, new_AGEMA_signal_12707, mcs1_mcs_mat1_7_mcs_out[65]}), .b ({new_AGEMA_signal_16546, new_AGEMA_signal_16545, new_AGEMA_signal_16544, mcs1_mcs_mat1_7_mcs_out[69]}), .c ({new_AGEMA_signal_17323, new_AGEMA_signal_17322, new_AGEMA_signal_17321, mcs1_mcs_mat1_7_n82}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U24 ( .a ({new_AGEMA_signal_17977, new_AGEMA_signal_17976, new_AGEMA_signal_17975, mcs1_mcs_mat1_7_n80}), .b ({new_AGEMA_signal_20761, new_AGEMA_signal_20760, new_AGEMA_signal_20759, mcs1_mcs_mat1_7_n79}), .c ({new_AGEMA_signal_21346, new_AGEMA_signal_21345, new_AGEMA_signal_21344, mcs_out[128]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U23 ( .a ({new_AGEMA_signal_20035, new_AGEMA_signal_20034, new_AGEMA_signal_20033, mcs1_mcs_mat1_7_mcs_out[72]}), .b ({new_AGEMA_signal_16537, new_AGEMA_signal_16536, new_AGEMA_signal_16535, mcs1_mcs_mat1_7_mcs_out[76]}), .c ({new_AGEMA_signal_20761, new_AGEMA_signal_20760, new_AGEMA_signal_20759, mcs1_mcs_mat1_7_n79}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U22 ( .a ({new_AGEMA_signal_17359, new_AGEMA_signal_17358, new_AGEMA_signal_17357, mcs1_mcs_mat1_7_mcs_out[64]}), .b ({new_AGEMA_signal_15592, new_AGEMA_signal_15591, new_AGEMA_signal_15590, mcs1_mcs_mat1_7_mcs_out[68]}), .c ({new_AGEMA_signal_17977, new_AGEMA_signal_17976, new_AGEMA_signal_17975, mcs1_mcs_mat1_7_n80}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U21 ( .a ({new_AGEMA_signal_16504, new_AGEMA_signal_16503, new_AGEMA_signal_16502, mcs1_mcs_mat1_7_n78}), .b ({new_AGEMA_signal_19282, new_AGEMA_signal_19281, new_AGEMA_signal_19280, mcs1_mcs_mat1_7_n77}), .c ({temp_next_s3[99], temp_next_s2[99], temp_next_s1[99], temp_next_s0[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U20 ( .a ({new_AGEMA_signal_18640, new_AGEMA_signal_18639, new_AGEMA_signal_18638, mcs1_mcs_mat1_7_mcs_out[59]}), .b ({new_AGEMA_signal_15601, new_AGEMA_signal_15600, new_AGEMA_signal_15599, mcs1_mcs_mat1_7_mcs_out[63]}), .c ({new_AGEMA_signal_19282, new_AGEMA_signal_19281, new_AGEMA_signal_19280, mcs1_mcs_mat1_7_n77}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U19 ( .a ({new_AGEMA_signal_12733, new_AGEMA_signal_12732, new_AGEMA_signal_12731, mcs1_mcs_mat1_7_mcs_out[51]}), .b ({new_AGEMA_signal_15616, new_AGEMA_signal_15615, new_AGEMA_signal_15614, mcs1_mcs_mat1_7_mcs_out[55]}), .c ({new_AGEMA_signal_16504, new_AGEMA_signal_16503, new_AGEMA_signal_16502, mcs1_mcs_mat1_7_n78}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U18 ( .a ({new_AGEMA_signal_17326, new_AGEMA_signal_17325, new_AGEMA_signal_17324, mcs1_mcs_mat1_7_n76}), .b ({new_AGEMA_signal_18619, new_AGEMA_signal_18618, new_AGEMA_signal_18617, mcs1_mcs_mat1_7_n75}), .c ({temp_next_s3[98], temp_next_s2[98], temp_next_s1[98], temp_next_s0[98]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U17 ( .a ({new_AGEMA_signal_18007, new_AGEMA_signal_18006, new_AGEMA_signal_18005, mcs1_mcs_mat1_7_mcs_out[58]}), .b ({new_AGEMA_signal_14158, new_AGEMA_signal_14157, new_AGEMA_signal_14156, mcs1_mcs_mat1_7_mcs_out[62]}), .c ({new_AGEMA_signal_18619, new_AGEMA_signal_18618, new_AGEMA_signal_18617, mcs1_mcs_mat1_7_n75}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U16 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_16558, new_AGEMA_signal_16557, new_AGEMA_signal_16556, mcs1_mcs_mat1_7_mcs_out[54]}), .c ({new_AGEMA_signal_17326, new_AGEMA_signal_17325, new_AGEMA_signal_17324, mcs1_mcs_mat1_7_n76}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U15 ( .a ({new_AGEMA_signal_17329, new_AGEMA_signal_17328, new_AGEMA_signal_17327, mcs1_mcs_mat1_7_n74}), .b ({new_AGEMA_signal_19288, new_AGEMA_signal_19287, new_AGEMA_signal_19286, mcs1_mcs_mat1_7_n73}), .c ({temp_next_s3[97], temp_next_s2[97], temp_next_s1[97], temp_next_s0[97]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U14 ( .a ({new_AGEMA_signal_18643, new_AGEMA_signal_18642, new_AGEMA_signal_18641, mcs1_mcs_mat1_7_mcs_out[57]}), .b ({new_AGEMA_signal_14161, new_AGEMA_signal_14160, new_AGEMA_signal_14159, mcs1_mcs_mat1_7_mcs_out[61]}), .c ({new_AGEMA_signal_19288, new_AGEMA_signal_19287, new_AGEMA_signal_19286, mcs1_mcs_mat1_7_n73}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U13 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({new_AGEMA_signal_16561, new_AGEMA_signal_16560, new_AGEMA_signal_16559, mcs1_mcs_mat1_7_mcs_out[53]}), .c ({new_AGEMA_signal_17329, new_AGEMA_signal_17328, new_AGEMA_signal_17327, mcs1_mcs_mat1_7_n74}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U12 ( .a ({new_AGEMA_signal_16507, new_AGEMA_signal_16506, new_AGEMA_signal_16505, mcs1_mcs_mat1_7_n72}), .b ({new_AGEMA_signal_20014, new_AGEMA_signal_20013, new_AGEMA_signal_20012, mcs1_mcs_mat1_7_n71}), .c ({temp_next_s3[96], temp_next_s2[96], temp_next_s1[96], temp_next_s0[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U11 ( .a ({new_AGEMA_signal_19318, new_AGEMA_signal_19317, new_AGEMA_signal_19316, mcs1_mcs_mat1_7_mcs_out[56]}), .b ({new_AGEMA_signal_16555, new_AGEMA_signal_16554, new_AGEMA_signal_16553, mcs1_mcs_mat1_7_mcs_out[60]}), .c ({new_AGEMA_signal_20014, new_AGEMA_signal_20013, new_AGEMA_signal_20012, mcs1_mcs_mat1_7_n71}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U10 ( .a ({new_AGEMA_signal_14176, new_AGEMA_signal_14175, new_AGEMA_signal_14174, mcs1_mcs_mat1_7_mcs_out[48]}), .b ({new_AGEMA_signal_15622, new_AGEMA_signal_15621, new_AGEMA_signal_15620, mcs1_mcs_mat1_7_mcs_out[52]}), .c ({new_AGEMA_signal_16507, new_AGEMA_signal_16506, new_AGEMA_signal_16505, mcs1_mcs_mat1_7_n72}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U9 ( .a ({new_AGEMA_signal_17332, new_AGEMA_signal_17331, new_AGEMA_signal_17330, mcs1_mcs_mat1_7_n70}), .b ({new_AGEMA_signal_20017, new_AGEMA_signal_20016, new_AGEMA_signal_20015, mcs1_mcs_mat1_7_n69}), .c ({temp_next_s3[67], temp_next_s2[67], temp_next_s1[67], temp_next_s0[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U8 ( .a ({new_AGEMA_signal_19321, new_AGEMA_signal_19320, new_AGEMA_signal_19319, mcs1_mcs_mat1_7_mcs_out[43]}), .b ({new_AGEMA_signal_15625, new_AGEMA_signal_15624, new_AGEMA_signal_15623, mcs1_mcs_mat1_7_mcs_out[47]}), .c ({new_AGEMA_signal_20017, new_AGEMA_signal_20016, new_AGEMA_signal_20015, mcs1_mcs_mat1_7_n69}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U7 ( .a ({new_AGEMA_signal_15634, new_AGEMA_signal_15633, new_AGEMA_signal_15632, mcs1_mcs_mat1_7_mcs_out[35]}), .b ({new_AGEMA_signal_16567, new_AGEMA_signal_16566, new_AGEMA_signal_16565, mcs1_mcs_mat1_7_mcs_out[39]}), .c ({new_AGEMA_signal_17332, new_AGEMA_signal_17331, new_AGEMA_signal_17330, mcs1_mcs_mat1_7_n70}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U6 ( .a ({new_AGEMA_signal_15523, new_AGEMA_signal_15522, new_AGEMA_signal_15521, mcs1_mcs_mat1_7_n68}), .b ({new_AGEMA_signal_20020, new_AGEMA_signal_20019, new_AGEMA_signal_20018, mcs1_mcs_mat1_7_n67}), .c ({temp_next_s3[66], temp_next_s2[66], temp_next_s1[66], temp_next_s0[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U5 ( .a ({new_AGEMA_signal_19324, new_AGEMA_signal_19323, new_AGEMA_signal_19322, mcs1_mcs_mat1_7_mcs_out[42]}), .b ({new_AGEMA_signal_11311, new_AGEMA_signal_11310, new_AGEMA_signal_11309, mcs1_mcs_mat1_7_mcs_out[46]}), .c ({new_AGEMA_signal_20020, new_AGEMA_signal_20019, new_AGEMA_signal_20018, mcs1_mcs_mat1_7_n67}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U4 ( .a ({new_AGEMA_signal_14191, new_AGEMA_signal_14190, new_AGEMA_signal_14189, mcs1_mcs_mat1_7_mcs_out[34]}), .b ({new_AGEMA_signal_12742, new_AGEMA_signal_12741, new_AGEMA_signal_12740, mcs1_mcs_mat1_7_mcs_out[38]}), .c ({new_AGEMA_signal_15523, new_AGEMA_signal_15522, new_AGEMA_signal_15521, mcs1_mcs_mat1_7_n68}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U3 ( .a ({new_AGEMA_signal_17980, new_AGEMA_signal_17979, new_AGEMA_signal_17978, mcs1_mcs_mat1_7_n66}), .b ({new_AGEMA_signal_20773, new_AGEMA_signal_20772, new_AGEMA_signal_20771, mcs1_mcs_mat1_7_n65}), .c ({temp_next_s3[0], temp_next_s2[0], temp_next_s1[0], temp_next_s0[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U2 ( .a ({new_AGEMA_signal_18043, new_AGEMA_signal_18042, new_AGEMA_signal_18041, mcs1_mcs_mat1_7_mcs_out[4]}), .b ({new_AGEMA_signal_20041, new_AGEMA_signal_20040, new_AGEMA_signal_20039, mcs1_mcs_mat1_7_mcs_out[8]}), .c ({new_AGEMA_signal_20773, new_AGEMA_signal_20772, new_AGEMA_signal_20771, mcs1_mcs_mat1_7_n65}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_U1 ( .a ({new_AGEMA_signal_15679, new_AGEMA_signal_15678, new_AGEMA_signal_15677, mcs1_mcs_mat1_7_mcs_out[0]}), .b ({new_AGEMA_signal_17380, new_AGEMA_signal_17379, new_AGEMA_signal_17378, mcs1_mcs_mat1_7_mcs_out[12]}), .c ({new_AGEMA_signal_17980, new_AGEMA_signal_17979, new_AGEMA_signal_17978, mcs1_mcs_mat1_7_n66}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U10 ( .a ({new_AGEMA_signal_19291, new_AGEMA_signal_19290, new_AGEMA_signal_19289, mcs1_mcs_mat1_7_mcs_rom0_1_n12}), .b ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_20023, new_AGEMA_signal_20022, new_AGEMA_signal_20021, mcs1_mcs_mat1_7_mcs_out[123]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U9 ( .a ({new_AGEMA_signal_18622, new_AGEMA_signal_18621, new_AGEMA_signal_18620, mcs1_mcs_mat1_7_mcs_rom0_1_n11}), .b ({new_AGEMA_signal_14086, new_AGEMA_signal_14085, new_AGEMA_signal_14084, mcs1_mcs_mat1_7_mcs_rom0_1_x0x4}), .c ({new_AGEMA_signal_19291, new_AGEMA_signal_19290, new_AGEMA_signal_19289, mcs1_mcs_mat1_7_mcs_rom0_1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U8 ( .a ({new_AGEMA_signal_15526, new_AGEMA_signal_15525, new_AGEMA_signal_15524, mcs1_mcs_mat1_7_mcs_rom0_1_n10}), .b ({new_AGEMA_signal_17335, new_AGEMA_signal_17334, new_AGEMA_signal_17333, mcs1_mcs_mat1_7_mcs_rom0_1_n9}), .c ({new_AGEMA_signal_17983, new_AGEMA_signal_17982, new_AGEMA_signal_17981, mcs1_mcs_mat1_7_mcs_out[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U7 ( .a ({new_AGEMA_signal_15529, new_AGEMA_signal_15528, new_AGEMA_signal_15527, mcs1_mcs_mat1_7_mcs_rom0_1_x2x4}), .b ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .c ({new_AGEMA_signal_17335, new_AGEMA_signal_17334, new_AGEMA_signal_17333, mcs1_mcs_mat1_7_mcs_rom0_1_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U5 ( .a ({new_AGEMA_signal_19294, new_AGEMA_signal_19293, new_AGEMA_signal_19292, mcs1_mcs_mat1_7_mcs_rom0_1_n8}), .b ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .c ({new_AGEMA_signal_20026, new_AGEMA_signal_20025, new_AGEMA_signal_20024, mcs1_mcs_mat1_7_mcs_out[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U4 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_18622, new_AGEMA_signal_18621, new_AGEMA_signal_18620, mcs1_mcs_mat1_7_mcs_rom0_1_n11}), .c ({new_AGEMA_signal_19294, new_AGEMA_signal_19293, new_AGEMA_signal_19292, mcs1_mcs_mat1_7_mcs_rom0_1_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U3 ( .a ({new_AGEMA_signal_17986, new_AGEMA_signal_17985, new_AGEMA_signal_17984, mcs1_mcs_mat1_7_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_17338, new_AGEMA_signal_17337, new_AGEMA_signal_17336, mcs1_mcs_mat1_7_mcs_rom0_1_x3x4}), .c ({new_AGEMA_signal_18622, new_AGEMA_signal_18621, new_AGEMA_signal_18620, mcs1_mcs_mat1_7_mcs_rom0_1_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U2 ( .a ({new_AGEMA_signal_18625, new_AGEMA_signal_18624, new_AGEMA_signal_18623, mcs1_mcs_mat1_7_mcs_rom0_1_n7}), .b ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_19297, new_AGEMA_signal_19296, new_AGEMA_signal_19295, mcs1_mcs_mat1_7_mcs_out[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_U1 ( .a ({new_AGEMA_signal_17986, new_AGEMA_signal_17985, new_AGEMA_signal_17984, mcs1_mcs_mat1_7_mcs_rom0_1_x1x4}), .b ({new_AGEMA_signal_15529, new_AGEMA_signal_15528, new_AGEMA_signal_15527, mcs1_mcs_mat1_7_mcs_rom0_1_x2x4}), .c ({new_AGEMA_signal_18625, new_AGEMA_signal_18624, new_AGEMA_signal_18623, mcs1_mcs_mat1_7_mcs_rom0_1_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6221], Fresh[6220], Fresh[6219], Fresh[6218], Fresh[6217], Fresh[6216]}), .c ({new_AGEMA_signal_17986, new_AGEMA_signal_17985, new_AGEMA_signal_17984, mcs1_mcs_mat1_7_mcs_rom0_1_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6227], Fresh[6226], Fresh[6225], Fresh[6224], Fresh[6223], Fresh[6222]}), .c ({new_AGEMA_signal_15529, new_AGEMA_signal_15528, new_AGEMA_signal_15527, mcs1_mcs_mat1_7_mcs_rom0_1_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_1_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6233], Fresh[6232], Fresh[6231], Fresh[6230], Fresh[6229], Fresh[6228]}), .c ({new_AGEMA_signal_17338, new_AGEMA_signal_17337, new_AGEMA_signal_17336, mcs1_mcs_mat1_7_mcs_rom0_1_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U11 ( .a ({new_AGEMA_signal_15532, new_AGEMA_signal_15531, new_AGEMA_signal_15530, mcs1_mcs_mat1_7_mcs_rom0_2_n14}), .b ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .c ({new_AGEMA_signal_16510, new_AGEMA_signal_16509, new_AGEMA_signal_16508, mcs1_mcs_mat1_7_mcs_out[119]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U10 ( .a ({new_AGEMA_signal_14089, new_AGEMA_signal_14088, new_AGEMA_signal_14087, mcs1_mcs_mat1_7_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_11257, new_AGEMA_signal_11256, new_AGEMA_signal_11255, mcs1_mcs_mat1_7_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_15532, new_AGEMA_signal_15531, new_AGEMA_signal_15530, mcs1_mcs_mat1_7_mcs_rom0_2_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U9 ( .a ({new_AGEMA_signal_15535, new_AGEMA_signal_15534, new_AGEMA_signal_15533, mcs1_mcs_mat1_7_mcs_rom0_2_n12}), .b ({new_AGEMA_signal_12634, new_AGEMA_signal_12633, new_AGEMA_signal_12632, mcs1_mcs_mat1_7_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_16513, new_AGEMA_signal_16512, new_AGEMA_signal_16511, mcs1_mcs_mat1_7_mcs_out[118]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U8 ( .a ({new_AGEMA_signal_14089, new_AGEMA_signal_14088, new_AGEMA_signal_14087, mcs1_mcs_mat1_7_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .c ({new_AGEMA_signal_15535, new_AGEMA_signal_15534, new_AGEMA_signal_15533, mcs1_mcs_mat1_7_mcs_rom0_2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U7 ( .a ({new_AGEMA_signal_14089, new_AGEMA_signal_14088, new_AGEMA_signal_14087, mcs1_mcs_mat1_7_mcs_rom0_2_n13}), .b ({new_AGEMA_signal_12631, new_AGEMA_signal_12630, new_AGEMA_signal_12629, mcs1_mcs_mat1_7_mcs_rom0_2_n10}), .c ({new_AGEMA_signal_15538, new_AGEMA_signal_15537, new_AGEMA_signal_15536, mcs1_mcs_mat1_7_mcs_out[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U4 ( .a ({new_AGEMA_signal_12637, new_AGEMA_signal_12636, new_AGEMA_signal_12635, mcs1_mcs_mat1_7_mcs_rom0_2_x1x4}), .b ({new_AGEMA_signal_9982, new_AGEMA_signal_9981, new_AGEMA_signal_9980, mcs1_mcs_mat1_7_mcs_rom0_2_x2x4}), .c ({new_AGEMA_signal_14089, new_AGEMA_signal_14088, new_AGEMA_signal_14087, mcs1_mcs_mat1_7_mcs_rom0_2_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U3 ( .a ({new_AGEMA_signal_11254, new_AGEMA_signal_11253, new_AGEMA_signal_11252, mcs1_mcs_mat1_7_mcs_rom0_2_n8}), .b ({new_AGEMA_signal_12634, new_AGEMA_signal_12633, new_AGEMA_signal_12632, mcs1_mcs_mat1_7_mcs_rom0_2_n11}), .c ({new_AGEMA_signal_14092, new_AGEMA_signal_14091, new_AGEMA_signal_14090, mcs1_mcs_mat1_7_mcs_out[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U2 ( .a ({new_AGEMA_signal_9079, new_AGEMA_signal_9078, new_AGEMA_signal_9077, mcs1_mcs_mat1_7_mcs_rom0_2_x0x4}), .b ({new_AGEMA_signal_11257, new_AGEMA_signal_11256, new_AGEMA_signal_11255, mcs1_mcs_mat1_7_mcs_rom0_2_x3x4}), .c ({new_AGEMA_signal_12634, new_AGEMA_signal_12633, new_AGEMA_signal_12632, mcs1_mcs_mat1_7_mcs_rom0_2_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_U1 ( .a ({new_AGEMA_signal_9982, new_AGEMA_signal_9981, new_AGEMA_signal_9980, mcs1_mcs_mat1_7_mcs_rom0_2_x2x4}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_11254, new_AGEMA_signal_11253, new_AGEMA_signal_11252, mcs1_mcs_mat1_7_mcs_rom0_2_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6239], Fresh[6238], Fresh[6237], Fresh[6236], Fresh[6235], Fresh[6234]}), .c ({new_AGEMA_signal_12637, new_AGEMA_signal_12636, new_AGEMA_signal_12635, mcs1_mcs_mat1_7_mcs_rom0_2_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6245], Fresh[6244], Fresh[6243], Fresh[6242], Fresh[6241], Fresh[6240]}), .c ({new_AGEMA_signal_9982, new_AGEMA_signal_9981, new_AGEMA_signal_9980, mcs1_mcs_mat1_7_mcs_rom0_2_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_2_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6251], Fresh[6250], Fresh[6249], Fresh[6248], Fresh[6247], Fresh[6246]}), .c ({new_AGEMA_signal_11257, new_AGEMA_signal_11256, new_AGEMA_signal_11255, mcs1_mcs_mat1_7_mcs_rom0_2_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U10 ( .a ({new_AGEMA_signal_14098, new_AGEMA_signal_14097, new_AGEMA_signal_14096, mcs1_mcs_mat1_7_mcs_rom0_3_n12}), .b ({new_AGEMA_signal_9985, new_AGEMA_signal_9984, new_AGEMA_signal_9983, mcs1_mcs_mat1_7_mcs_rom0_3_n11}), .c ({new_AGEMA_signal_15541, new_AGEMA_signal_15540, new_AGEMA_signal_15539, mcs1_mcs_mat1_7_mcs_out[115]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U8 ( .a ({new_AGEMA_signal_11260, new_AGEMA_signal_11259, new_AGEMA_signal_11258, mcs1_mcs_mat1_7_mcs_rom0_3_n9}), .b ({new_AGEMA_signal_11263, new_AGEMA_signal_11262, new_AGEMA_signal_11261, mcs1_mcs_mat1_7_mcs_rom0_3_x3x4}), .c ({new_AGEMA_signal_12640, new_AGEMA_signal_12639, new_AGEMA_signal_12638, mcs1_mcs_mat1_7_mcs_out[113]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U5 ( .a ({new_AGEMA_signal_14101, new_AGEMA_signal_14100, new_AGEMA_signal_14099, mcs1_mcs_mat1_7_mcs_rom0_3_n8}), .b ({new_AGEMA_signal_15544, new_AGEMA_signal_15543, new_AGEMA_signal_15542, mcs1_mcs_mat1_7_mcs_rom0_3_n7}), .c ({new_AGEMA_signal_16516, new_AGEMA_signal_16515, new_AGEMA_signal_16514, mcs1_mcs_mat1_7_mcs_out[112]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U4 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_14098, new_AGEMA_signal_14097, new_AGEMA_signal_14096, mcs1_mcs_mat1_7_mcs_rom0_3_n12}), .c ({new_AGEMA_signal_15544, new_AGEMA_signal_15543, new_AGEMA_signal_15542, mcs1_mcs_mat1_7_mcs_rom0_3_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U3 ( .a ({new_AGEMA_signal_9082, new_AGEMA_signal_9081, new_AGEMA_signal_9080, mcs1_mcs_mat1_7_mcs_rom0_3_x0x4}), .b ({new_AGEMA_signal_12646, new_AGEMA_signal_12645, new_AGEMA_signal_12644, mcs1_mcs_mat1_7_mcs_rom0_3_x1x4}), .c ({new_AGEMA_signal_14098, new_AGEMA_signal_14097, new_AGEMA_signal_14096, mcs1_mcs_mat1_7_mcs_rom0_3_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_U2 ( .a ({new_AGEMA_signal_9988, new_AGEMA_signal_9987, new_AGEMA_signal_9986, mcs1_mcs_mat1_7_mcs_rom0_3_x2x4}), .b ({new_AGEMA_signal_12643, new_AGEMA_signal_12642, new_AGEMA_signal_12641, mcs1_mcs_mat1_7_mcs_rom0_3_n10}), .c ({new_AGEMA_signal_14101, new_AGEMA_signal_14100, new_AGEMA_signal_14099, mcs1_mcs_mat1_7_mcs_rom0_3_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6257], Fresh[6256], Fresh[6255], Fresh[6254], Fresh[6253], Fresh[6252]}), .c ({new_AGEMA_signal_12646, new_AGEMA_signal_12645, new_AGEMA_signal_12644, mcs1_mcs_mat1_7_mcs_rom0_3_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6263], Fresh[6262], Fresh[6261], Fresh[6260], Fresh[6259], Fresh[6258]}), .c ({new_AGEMA_signal_9988, new_AGEMA_signal_9987, new_AGEMA_signal_9986, mcs1_mcs_mat1_7_mcs_rom0_3_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_3_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6269], Fresh[6268], Fresh[6267], Fresh[6266], Fresh[6265], Fresh[6264]}), .c ({new_AGEMA_signal_11263, new_AGEMA_signal_11262, new_AGEMA_signal_11261, mcs1_mcs_mat1_7_mcs_rom0_3_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U9 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({new_AGEMA_signal_15547, new_AGEMA_signal_15546, new_AGEMA_signal_15545, mcs1_mcs_mat1_7_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_16519, new_AGEMA_signal_16518, new_AGEMA_signal_16517, mcs1_mcs_mat1_7_mcs_out[111]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U8 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({new_AGEMA_signal_15550, new_AGEMA_signal_15549, new_AGEMA_signal_15548, mcs1_mcs_mat1_7_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_16522, new_AGEMA_signal_16521, new_AGEMA_signal_16520, mcs1_mcs_mat1_7_mcs_out[110]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U7 ( .a ({new_AGEMA_signal_11266, new_AGEMA_signal_11265, new_AGEMA_signal_11264, mcs1_mcs_mat1_7_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_15547, new_AGEMA_signal_15546, new_AGEMA_signal_15545, mcs1_mcs_mat1_7_mcs_rom0_4_n10}), .c ({new_AGEMA_signal_16525, new_AGEMA_signal_16524, new_AGEMA_signal_16523, mcs1_mcs_mat1_7_mcs_out[109]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U6 ( .a ({new_AGEMA_signal_9991, new_AGEMA_signal_9990, new_AGEMA_signal_9989, mcs1_mcs_mat1_7_mcs_rom0_4_x2x4}), .b ({new_AGEMA_signal_14104, new_AGEMA_signal_14103, new_AGEMA_signal_14102, mcs1_mcs_mat1_7_mcs_rom0_4_n8}), .c ({new_AGEMA_signal_15547, new_AGEMA_signal_15546, new_AGEMA_signal_15545, mcs1_mcs_mat1_7_mcs_rom0_4_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U4 ( .a ({new_AGEMA_signal_12649, new_AGEMA_signal_12648, new_AGEMA_signal_12647, mcs1_mcs_mat1_7_mcs_rom0_4_n7}), .b ({new_AGEMA_signal_15550, new_AGEMA_signal_15549, new_AGEMA_signal_15548, mcs1_mcs_mat1_7_mcs_rom0_4_n9}), .c ({new_AGEMA_signal_16528, new_AGEMA_signal_16527, new_AGEMA_signal_16526, mcs1_mcs_mat1_7_mcs_out[108]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U3 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_14107, new_AGEMA_signal_14106, new_AGEMA_signal_14105, mcs1_mcs_mat1_7_mcs_rom0_4_n6}), .c ({new_AGEMA_signal_15550, new_AGEMA_signal_15549, new_AGEMA_signal_15548, mcs1_mcs_mat1_7_mcs_rom0_4_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_U2 ( .a ({new_AGEMA_signal_11266, new_AGEMA_signal_11265, new_AGEMA_signal_11264, mcs1_mcs_mat1_7_mcs_rom0_4_x3x4}), .b ({new_AGEMA_signal_12652, new_AGEMA_signal_12651, new_AGEMA_signal_12650, mcs1_mcs_mat1_7_mcs_rom0_4_x1x4}), .c ({new_AGEMA_signal_14107, new_AGEMA_signal_14106, new_AGEMA_signal_14105, mcs1_mcs_mat1_7_mcs_rom0_4_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6275], Fresh[6274], Fresh[6273], Fresh[6272], Fresh[6271], Fresh[6270]}), .c ({new_AGEMA_signal_12652, new_AGEMA_signal_12651, new_AGEMA_signal_12650, mcs1_mcs_mat1_7_mcs_rom0_4_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6281], Fresh[6280], Fresh[6279], Fresh[6278], Fresh[6277], Fresh[6276]}), .c ({new_AGEMA_signal_9991, new_AGEMA_signal_9990, new_AGEMA_signal_9989, mcs1_mcs_mat1_7_mcs_rom0_4_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_4_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6287], Fresh[6286], Fresh[6285], Fresh[6284], Fresh[6283], Fresh[6282]}), .c ({new_AGEMA_signal_11266, new_AGEMA_signal_11265, new_AGEMA_signal_11264, mcs1_mcs_mat1_7_mcs_rom0_4_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U9 ( .a ({new_AGEMA_signal_18631, new_AGEMA_signal_18630, new_AGEMA_signal_18629, mcs1_mcs_mat1_7_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_18628, new_AGEMA_signal_18627, new_AGEMA_signal_18626, mcs1_mcs_mat1_7_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_19300, new_AGEMA_signal_19299, new_AGEMA_signal_19298, mcs1_mcs_mat1_7_mcs_out[107]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U8 ( .a ({new_AGEMA_signal_18628, new_AGEMA_signal_18627, new_AGEMA_signal_18626, mcs1_mcs_mat1_7_mcs_rom0_5_n10}), .b ({new_AGEMA_signal_17341, new_AGEMA_signal_17340, new_AGEMA_signal_17339, mcs1_mcs_mat1_7_mcs_rom0_5_n9}), .c ({new_AGEMA_signal_19303, new_AGEMA_signal_19302, new_AGEMA_signal_19301, mcs1_mcs_mat1_7_mcs_out[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U7 ( .a ({new_AGEMA_signal_15553, new_AGEMA_signal_15552, new_AGEMA_signal_15551, mcs1_mcs_mat1_7_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .c ({new_AGEMA_signal_17341, new_AGEMA_signal_17340, new_AGEMA_signal_17339, mcs1_mcs_mat1_7_mcs_rom0_5_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U6 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({new_AGEMA_signal_18628, new_AGEMA_signal_18627, new_AGEMA_signal_18626, mcs1_mcs_mat1_7_mcs_rom0_5_n10}), .c ({new_AGEMA_signal_19306, new_AGEMA_signal_19305, new_AGEMA_signal_19304, mcs1_mcs_mat1_7_mcs_out[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U5 ( .a ({new_AGEMA_signal_17992, new_AGEMA_signal_17991, new_AGEMA_signal_17990, mcs1_mcs_mat1_7_mcs_rom0_5_x1x4}), .b ({new_AGEMA_signal_14110, new_AGEMA_signal_14109, new_AGEMA_signal_14108, mcs1_mcs_mat1_7_mcs_rom0_5_x0x4}), .c ({new_AGEMA_signal_18628, new_AGEMA_signal_18627, new_AGEMA_signal_18626, mcs1_mcs_mat1_7_mcs_rom0_5_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U4 ( .a ({new_AGEMA_signal_19309, new_AGEMA_signal_19308, new_AGEMA_signal_19307, mcs1_mcs_mat1_7_mcs_rom0_5_n8}), .b ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_20029, new_AGEMA_signal_20028, new_AGEMA_signal_20027, mcs1_mcs_mat1_7_mcs_out[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U3 ( .a ({new_AGEMA_signal_18631, new_AGEMA_signal_18630, new_AGEMA_signal_18629, mcs1_mcs_mat1_7_mcs_rom0_5_n11}), .b ({new_AGEMA_signal_17992, new_AGEMA_signal_17991, new_AGEMA_signal_17990, mcs1_mcs_mat1_7_mcs_rom0_5_x1x4}), .c ({new_AGEMA_signal_19309, new_AGEMA_signal_19308, new_AGEMA_signal_19307, mcs1_mcs_mat1_7_mcs_rom0_5_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U2 ( .a ({new_AGEMA_signal_17989, new_AGEMA_signal_17988, new_AGEMA_signal_17987, mcs1_mcs_mat1_7_mcs_rom0_5_n7}), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .c ({new_AGEMA_signal_18631, new_AGEMA_signal_18630, new_AGEMA_signal_18629, mcs1_mcs_mat1_7_mcs_rom0_5_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_U1 ( .a ({new_AGEMA_signal_15553, new_AGEMA_signal_15552, new_AGEMA_signal_15551, mcs1_mcs_mat1_7_mcs_rom0_5_x2x4}), .b ({new_AGEMA_signal_17344, new_AGEMA_signal_17343, new_AGEMA_signal_17342, mcs1_mcs_mat1_7_mcs_rom0_5_x3x4}), .c ({new_AGEMA_signal_17989, new_AGEMA_signal_17988, new_AGEMA_signal_17987, mcs1_mcs_mat1_7_mcs_rom0_5_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6293], Fresh[6292], Fresh[6291], Fresh[6290], Fresh[6289], Fresh[6288]}), .c ({new_AGEMA_signal_17992, new_AGEMA_signal_17991, new_AGEMA_signal_17990, mcs1_mcs_mat1_7_mcs_rom0_5_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6299], Fresh[6298], Fresh[6297], Fresh[6296], Fresh[6295], Fresh[6294]}), .c ({new_AGEMA_signal_15553, new_AGEMA_signal_15552, new_AGEMA_signal_15551, mcs1_mcs_mat1_7_mcs_rom0_5_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_5_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6305], Fresh[6304], Fresh[6303], Fresh[6302], Fresh[6301], Fresh[6300]}), .c ({new_AGEMA_signal_17344, new_AGEMA_signal_17343, new_AGEMA_signal_17342, mcs1_mcs_mat1_7_mcs_rom0_5_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U9 ( .a ({new_AGEMA_signal_11269, new_AGEMA_signal_11268, new_AGEMA_signal_11267, mcs1_mcs_mat1_7_mcs_rom0_6_n10}), .b ({new_AGEMA_signal_14113, new_AGEMA_signal_14112, new_AGEMA_signal_14111, mcs1_mcs_mat1_7_mcs_rom0_6_n9}), .c ({new_AGEMA_signal_15556, new_AGEMA_signal_15555, new_AGEMA_signal_15554, mcs1_mcs_mat1_7_mcs_out[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U8 ( .a ({new_AGEMA_signal_12664, new_AGEMA_signal_12663, new_AGEMA_signal_12662, mcs1_mcs_mat1_7_mcs_rom0_6_x1x4}), .b ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_14113, new_AGEMA_signal_14112, new_AGEMA_signal_14111, mcs1_mcs_mat1_7_mcs_rom0_6_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U5 ( .a ({new_AGEMA_signal_12658, new_AGEMA_signal_12657, new_AGEMA_signal_12656, mcs1_mcs_mat1_7_mcs_rom0_6_n8}), .b ({new_AGEMA_signal_11272, new_AGEMA_signal_11271, new_AGEMA_signal_11270, mcs1_mcs_mat1_7_mcs_rom0_6_x3x4}), .c ({new_AGEMA_signal_14116, new_AGEMA_signal_14115, new_AGEMA_signal_14114, mcs1_mcs_mat1_7_mcs_out[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U3 ( .a ({new_AGEMA_signal_12661, new_AGEMA_signal_12660, new_AGEMA_signal_12659, mcs1_mcs_mat1_7_mcs_rom0_6_n7}), .b ({new_AGEMA_signal_14119, new_AGEMA_signal_14118, new_AGEMA_signal_14117, mcs1_mcs_mat1_7_mcs_rom0_6_n6}), .c ({new_AGEMA_signal_15559, new_AGEMA_signal_15558, new_AGEMA_signal_15557, mcs1_mcs_mat1_7_mcs_out[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U2 ( .a ({new_AGEMA_signal_9088, new_AGEMA_signal_9087, new_AGEMA_signal_9086, mcs1_mcs_mat1_7_mcs_rom0_6_x0x4}), .b ({new_AGEMA_signal_12664, new_AGEMA_signal_12663, new_AGEMA_signal_12662, mcs1_mcs_mat1_7_mcs_rom0_6_x1x4}), .c ({new_AGEMA_signal_14119, new_AGEMA_signal_14118, new_AGEMA_signal_14117, mcs1_mcs_mat1_7_mcs_rom0_6_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_U1 ( .a ({new_AGEMA_signal_9994, new_AGEMA_signal_9993, new_AGEMA_signal_9992, mcs1_mcs_mat1_7_mcs_rom0_6_x2x4}), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .c ({new_AGEMA_signal_12661, new_AGEMA_signal_12660, new_AGEMA_signal_12659, mcs1_mcs_mat1_7_mcs_rom0_6_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6311], Fresh[6310], Fresh[6309], Fresh[6308], Fresh[6307], Fresh[6306]}), .c ({new_AGEMA_signal_12664, new_AGEMA_signal_12663, new_AGEMA_signal_12662, mcs1_mcs_mat1_7_mcs_rom0_6_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6317], Fresh[6316], Fresh[6315], Fresh[6314], Fresh[6313], Fresh[6312]}), .c ({new_AGEMA_signal_9994, new_AGEMA_signal_9993, new_AGEMA_signal_9992, mcs1_mcs_mat1_7_mcs_rom0_6_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_6_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6323], Fresh[6322], Fresh[6321], Fresh[6320], Fresh[6319], Fresh[6318]}), .c ({new_AGEMA_signal_11272, new_AGEMA_signal_11271, new_AGEMA_signal_11270, mcs1_mcs_mat1_7_mcs_rom0_6_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U6 ( .a ({new_AGEMA_signal_17347, new_AGEMA_signal_17346, new_AGEMA_signal_17345, mcs1_mcs_mat1_7_mcs_rom0_7_n7}), .b ({new_AGEMA_signal_11278, new_AGEMA_signal_11277, new_AGEMA_signal_11276, mcs1_mcs_mat1_7_mcs_rom0_7_x3x4}), .c ({new_AGEMA_signal_17995, new_AGEMA_signal_17994, new_AGEMA_signal_17993, mcs1_mcs_mat1_7_mcs_out[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U5 ( .a ({new_AGEMA_signal_16531, new_AGEMA_signal_16530, new_AGEMA_signal_16529, mcs1_mcs_mat1_7_mcs_out[99]}), .b ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .c ({new_AGEMA_signal_17347, new_AGEMA_signal_17346, new_AGEMA_signal_17345, mcs1_mcs_mat1_7_mcs_rom0_7_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U4 ( .a ({new_AGEMA_signal_15562, new_AGEMA_signal_15561, new_AGEMA_signal_15560, mcs1_mcs_mat1_7_mcs_rom0_7_n6}), .b ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .c ({new_AGEMA_signal_16531, new_AGEMA_signal_16530, new_AGEMA_signal_16529, mcs1_mcs_mat1_7_mcs_out[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U3 ( .a ({new_AGEMA_signal_14122, new_AGEMA_signal_14121, new_AGEMA_signal_14120, mcs1_mcs_mat1_7_mcs_out[98]}), .b ({new_AGEMA_signal_10000, new_AGEMA_signal_9999, new_AGEMA_signal_9998, mcs1_mcs_mat1_7_mcs_rom0_7_x2x4}), .c ({new_AGEMA_signal_15562, new_AGEMA_signal_15561, new_AGEMA_signal_15560, mcs1_mcs_mat1_7_mcs_rom0_7_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_U2 ( .a ({new_AGEMA_signal_9997, new_AGEMA_signal_9996, new_AGEMA_signal_9995, mcs1_mcs_mat1_7_mcs_rom0_7_n5}), .b ({new_AGEMA_signal_12667, new_AGEMA_signal_12666, new_AGEMA_signal_12665, mcs1_mcs_mat1_7_mcs_rom0_7_x1x4}), .c ({new_AGEMA_signal_14122, new_AGEMA_signal_14121, new_AGEMA_signal_14120, mcs1_mcs_mat1_7_mcs_out[98]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6329], Fresh[6328], Fresh[6327], Fresh[6326], Fresh[6325], Fresh[6324]}), .c ({new_AGEMA_signal_12667, new_AGEMA_signal_12666, new_AGEMA_signal_12665, mcs1_mcs_mat1_7_mcs_rom0_7_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6335], Fresh[6334], Fresh[6333], Fresh[6332], Fresh[6331], Fresh[6330]}), .c ({new_AGEMA_signal_10000, new_AGEMA_signal_9999, new_AGEMA_signal_9998, mcs1_mcs_mat1_7_mcs_rom0_7_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_7_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6341], Fresh[6340], Fresh[6339], Fresh[6338], Fresh[6337], Fresh[6336]}), .c ({new_AGEMA_signal_11278, new_AGEMA_signal_11277, new_AGEMA_signal_11276, mcs1_mcs_mat1_7_mcs_rom0_7_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U8 ( .a ({new_AGEMA_signal_14125, new_AGEMA_signal_14124, new_AGEMA_signal_14123, mcs1_mcs_mat1_7_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_15565, new_AGEMA_signal_15564, new_AGEMA_signal_15563, mcs1_mcs_mat1_7_mcs_out[95]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U5 ( .a ({new_AGEMA_signal_11284, new_AGEMA_signal_11283, new_AGEMA_signal_11282, mcs1_mcs_mat1_7_mcs_rom0_8_n6}), .b ({new_AGEMA_signal_11287, new_AGEMA_signal_11286, new_AGEMA_signal_11285, mcs1_mcs_mat1_7_mcs_rom0_8_x3x4}), .c ({new_AGEMA_signal_12673, new_AGEMA_signal_12672, new_AGEMA_signal_12671, mcs1_mcs_mat1_7_mcs_out[93]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U3 ( .a ({new_AGEMA_signal_15568, new_AGEMA_signal_15567, new_AGEMA_signal_15566, mcs1_mcs_mat1_7_mcs_rom0_8_n5}), .b ({new_AGEMA_signal_10003, new_AGEMA_signal_10002, new_AGEMA_signal_10001, mcs1_mcs_mat1_7_mcs_rom0_8_x2x4}), .c ({new_AGEMA_signal_16534, new_AGEMA_signal_16533, new_AGEMA_signal_16532, mcs1_mcs_mat1_7_mcs_out[92]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U2 ( .a ({new_AGEMA_signal_14125, new_AGEMA_signal_14124, new_AGEMA_signal_14123, mcs1_mcs_mat1_7_mcs_rom0_8_n8}), .b ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .c ({new_AGEMA_signal_15568, new_AGEMA_signal_15567, new_AGEMA_signal_15566, mcs1_mcs_mat1_7_mcs_rom0_8_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_U1 ( .a ({new_AGEMA_signal_9094, new_AGEMA_signal_9093, new_AGEMA_signal_9092, mcs1_mcs_mat1_7_mcs_rom0_8_x0x4}), .b ({new_AGEMA_signal_12676, new_AGEMA_signal_12675, new_AGEMA_signal_12674, mcs1_mcs_mat1_7_mcs_rom0_8_x1x4}), .c ({new_AGEMA_signal_14125, new_AGEMA_signal_14124, new_AGEMA_signal_14123, mcs1_mcs_mat1_7_mcs_rom0_8_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6347], Fresh[6346], Fresh[6345], Fresh[6344], Fresh[6343], Fresh[6342]}), .c ({new_AGEMA_signal_12676, new_AGEMA_signal_12675, new_AGEMA_signal_12674, mcs1_mcs_mat1_7_mcs_rom0_8_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6353], Fresh[6352], Fresh[6351], Fresh[6350], Fresh[6349], Fresh[6348]}), .c ({new_AGEMA_signal_10003, new_AGEMA_signal_10002, new_AGEMA_signal_10001, mcs1_mcs_mat1_7_mcs_rom0_8_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_8_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6359], Fresh[6358], Fresh[6357], Fresh[6356], Fresh[6355], Fresh[6354]}), .c ({new_AGEMA_signal_11287, new_AGEMA_signal_11286, new_AGEMA_signal_11285, mcs1_mcs_mat1_7_mcs_rom0_8_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U8 ( .a ({new_AGEMA_signal_12688, new_AGEMA_signal_12687, new_AGEMA_signal_12686, mcs1_mcs_mat1_7_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_12691, new_AGEMA_signal_12690, new_AGEMA_signal_12689, mcs1_mcs_mat1_7_mcs_rom0_11_x1x4}), .c ({new_AGEMA_signal_14131, new_AGEMA_signal_14130, new_AGEMA_signal_14129, mcs1_mcs_mat1_7_mcs_out[83]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U7 ( .a ({new_AGEMA_signal_12682, new_AGEMA_signal_12681, new_AGEMA_signal_12680, mcs1_mcs_mat1_7_mcs_rom0_11_n7}), .b ({new_AGEMA_signal_9097, new_AGEMA_signal_9096, new_AGEMA_signal_9095, mcs1_mcs_mat1_7_mcs_rom0_11_x0x4}), .c ({new_AGEMA_signal_14134, new_AGEMA_signal_14133, new_AGEMA_signal_14132, mcs1_mcs_mat1_7_mcs_out[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U6 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_11290, new_AGEMA_signal_11289, new_AGEMA_signal_11288, mcs1_mcs_mat1_7_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_12682, new_AGEMA_signal_12681, new_AGEMA_signal_12680, mcs1_mcs_mat1_7_mcs_rom0_11_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U5 ( .a ({new_AGEMA_signal_12685, new_AGEMA_signal_12684, new_AGEMA_signal_12683, mcs1_mcs_mat1_7_mcs_rom0_11_n6}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_14137, new_AGEMA_signal_14136, new_AGEMA_signal_14135, mcs1_mcs_mat1_7_mcs_out[81]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U4 ( .a ({new_AGEMA_signal_10006, new_AGEMA_signal_10005, new_AGEMA_signal_10004, mcs1_mcs_mat1_7_mcs_rom0_11_x2x4}), .b ({new_AGEMA_signal_11290, new_AGEMA_signal_11289, new_AGEMA_signal_11288, mcs1_mcs_mat1_7_mcs_rom0_11_x3x4}), .c ({new_AGEMA_signal_12685, new_AGEMA_signal_12684, new_AGEMA_signal_12683, mcs1_mcs_mat1_7_mcs_rom0_11_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U3 ( .a ({new_AGEMA_signal_14140, new_AGEMA_signal_14139, new_AGEMA_signal_14138, mcs1_mcs_mat1_7_mcs_rom0_11_n5}), .b ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .c ({new_AGEMA_signal_15571, new_AGEMA_signal_15570, new_AGEMA_signal_15569, mcs1_mcs_mat1_7_mcs_out[80]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_U2 ( .a ({new_AGEMA_signal_12688, new_AGEMA_signal_12687, new_AGEMA_signal_12686, mcs1_mcs_mat1_7_mcs_rom0_11_n8}), .b ({new_AGEMA_signal_10006, new_AGEMA_signal_10005, new_AGEMA_signal_10004, mcs1_mcs_mat1_7_mcs_rom0_11_x2x4}), .c ({new_AGEMA_signal_14140, new_AGEMA_signal_14139, new_AGEMA_signal_14138, mcs1_mcs_mat1_7_mcs_rom0_11_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6365], Fresh[6364], Fresh[6363], Fresh[6362], Fresh[6361], Fresh[6360]}), .c ({new_AGEMA_signal_12691, new_AGEMA_signal_12690, new_AGEMA_signal_12689, mcs1_mcs_mat1_7_mcs_rom0_11_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6371], Fresh[6370], Fresh[6369], Fresh[6368], Fresh[6367], Fresh[6366]}), .c ({new_AGEMA_signal_10006, new_AGEMA_signal_10005, new_AGEMA_signal_10004, mcs1_mcs_mat1_7_mcs_rom0_11_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_11_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6377], Fresh[6376], Fresh[6375], Fresh[6374], Fresh[6373], Fresh[6372]}), .c ({new_AGEMA_signal_11290, new_AGEMA_signal_11289, new_AGEMA_signal_11288, mcs1_mcs_mat1_7_mcs_rom0_11_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U6 ( .a ({new_AGEMA_signal_14143, new_AGEMA_signal_14142, new_AGEMA_signal_14141, mcs1_mcs_mat1_7_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_15574, new_AGEMA_signal_15573, new_AGEMA_signal_15572, mcs1_mcs_mat1_7_mcs_out[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U4 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_11293, new_AGEMA_signal_11292, new_AGEMA_signal_11291, mcs1_mcs_mat1_7_mcs_rom0_12_x3x4}), .c ({new_AGEMA_signal_12694, new_AGEMA_signal_12693, new_AGEMA_signal_12692, mcs1_mcs_mat1_7_mcs_out[77]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U3 ( .a ({new_AGEMA_signal_15577, new_AGEMA_signal_15576, new_AGEMA_signal_15575, mcs1_mcs_mat1_7_mcs_rom0_12_n3}), .b ({new_AGEMA_signal_10012, new_AGEMA_signal_10011, new_AGEMA_signal_10010, mcs1_mcs_mat1_7_mcs_rom0_12_x2x4}), .c ({new_AGEMA_signal_16537, new_AGEMA_signal_16536, new_AGEMA_signal_16535, mcs1_mcs_mat1_7_mcs_out[76]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U2 ( .a ({new_AGEMA_signal_14143, new_AGEMA_signal_14142, new_AGEMA_signal_14141, mcs1_mcs_mat1_7_mcs_rom0_12_n4}), .b ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .c ({new_AGEMA_signal_15577, new_AGEMA_signal_15576, new_AGEMA_signal_15575, mcs1_mcs_mat1_7_mcs_rom0_12_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_U1 ( .a ({new_AGEMA_signal_9100, new_AGEMA_signal_9099, new_AGEMA_signal_9098, mcs1_mcs_mat1_7_mcs_rom0_12_x0x4}), .b ({new_AGEMA_signal_12697, new_AGEMA_signal_12696, new_AGEMA_signal_12695, mcs1_mcs_mat1_7_mcs_rom0_12_x1x4}), .c ({new_AGEMA_signal_14143, new_AGEMA_signal_14142, new_AGEMA_signal_14141, mcs1_mcs_mat1_7_mcs_rom0_12_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6383], Fresh[6382], Fresh[6381], Fresh[6380], Fresh[6379], Fresh[6378]}), .c ({new_AGEMA_signal_12697, new_AGEMA_signal_12696, new_AGEMA_signal_12695, mcs1_mcs_mat1_7_mcs_rom0_12_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6389], Fresh[6388], Fresh[6387], Fresh[6386], Fresh[6385], Fresh[6384]}), .c ({new_AGEMA_signal_10012, new_AGEMA_signal_10011, new_AGEMA_signal_10010, mcs1_mcs_mat1_7_mcs_rom0_12_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_12_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6395], Fresh[6394], Fresh[6393], Fresh[6392], Fresh[6391], Fresh[6390]}), .c ({new_AGEMA_signal_11293, new_AGEMA_signal_11292, new_AGEMA_signal_11291, mcs1_mcs_mat1_7_mcs_rom0_12_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U10 ( .a ({new_AGEMA_signal_19312, new_AGEMA_signal_19311, new_AGEMA_signal_19310, mcs1_mcs_mat1_7_mcs_rom0_13_n14}), .b ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_20032, new_AGEMA_signal_20031, new_AGEMA_signal_20030, mcs1_mcs_mat1_7_mcs_out[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U9 ( .a ({new_AGEMA_signal_18637, new_AGEMA_signal_18636, new_AGEMA_signal_18635, mcs1_mcs_mat1_7_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_18001, new_AGEMA_signal_18000, new_AGEMA_signal_17999, mcs1_mcs_mat1_7_mcs_rom0_13_n12}), .c ({new_AGEMA_signal_19312, new_AGEMA_signal_19311, new_AGEMA_signal_19310, mcs1_mcs_mat1_7_mcs_rom0_13_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U8 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({new_AGEMA_signal_16540, new_AGEMA_signal_16539, new_AGEMA_signal_16538, mcs1_mcs_mat1_7_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_17998, new_AGEMA_signal_17997, new_AGEMA_signal_17996, mcs1_mcs_mat1_7_mcs_out[75]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U7 ( .a ({new_AGEMA_signal_18001, new_AGEMA_signal_18000, new_AGEMA_signal_17999, mcs1_mcs_mat1_7_mcs_rom0_13_n12}), .b ({new_AGEMA_signal_16540, new_AGEMA_signal_16539, new_AGEMA_signal_16538, mcs1_mcs_mat1_7_mcs_rom0_13_n11}), .c ({new_AGEMA_signal_18634, new_AGEMA_signal_18633, new_AGEMA_signal_18632, mcs1_mcs_mat1_7_mcs_out[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U6 ( .a ({new_AGEMA_signal_15580, new_AGEMA_signal_15579, new_AGEMA_signal_15578, mcs1_mcs_mat1_7_mcs_rom0_13_n10}), .b ({new_AGEMA_signal_15583, new_AGEMA_signal_15582, new_AGEMA_signal_15581, mcs1_mcs_mat1_7_mcs_rom0_13_x2x4}), .c ({new_AGEMA_signal_16540, new_AGEMA_signal_16539, new_AGEMA_signal_16538, mcs1_mcs_mat1_7_mcs_rom0_13_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U5 ( .a ({new_AGEMA_signal_17356, new_AGEMA_signal_17355, new_AGEMA_signal_17354, mcs1_mcs_mat1_7_mcs_rom0_13_x3x4}), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .c ({new_AGEMA_signal_18001, new_AGEMA_signal_18000, new_AGEMA_signal_17999, mcs1_mcs_mat1_7_mcs_rom0_13_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U4 ( .a ({new_AGEMA_signal_19315, new_AGEMA_signal_19314, new_AGEMA_signal_19313, mcs1_mcs_mat1_7_mcs_rom0_13_n9}), .b ({new_AGEMA_signal_15580, new_AGEMA_signal_15579, new_AGEMA_signal_15578, mcs1_mcs_mat1_7_mcs_rom0_13_n10}), .c ({new_AGEMA_signal_20035, new_AGEMA_signal_20034, new_AGEMA_signal_20033, mcs1_mcs_mat1_7_mcs_out[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U2 ( .a ({new_AGEMA_signal_18637, new_AGEMA_signal_18636, new_AGEMA_signal_18635, mcs1_mcs_mat1_7_mcs_rom0_13_n13}), .b ({new_AGEMA_signal_17356, new_AGEMA_signal_17355, new_AGEMA_signal_17354, mcs1_mcs_mat1_7_mcs_rom0_13_x3x4}), .c ({new_AGEMA_signal_19315, new_AGEMA_signal_19314, new_AGEMA_signal_19313, mcs1_mcs_mat1_7_mcs_rom0_13_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_U1 ( .a ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .b ({new_AGEMA_signal_18004, new_AGEMA_signal_18003, new_AGEMA_signal_18002, mcs1_mcs_mat1_7_mcs_rom0_13_x1x4}), .c ({new_AGEMA_signal_18637, new_AGEMA_signal_18636, new_AGEMA_signal_18635, mcs1_mcs_mat1_7_mcs_rom0_13_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6401], Fresh[6400], Fresh[6399], Fresh[6398], Fresh[6397], Fresh[6396]}), .c ({new_AGEMA_signal_18004, new_AGEMA_signal_18003, new_AGEMA_signal_18002, mcs1_mcs_mat1_7_mcs_rom0_13_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6407], Fresh[6406], Fresh[6405], Fresh[6404], Fresh[6403], Fresh[6402]}), .c ({new_AGEMA_signal_15583, new_AGEMA_signal_15582, new_AGEMA_signal_15581, mcs1_mcs_mat1_7_mcs_rom0_13_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_13_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6413], Fresh[6412], Fresh[6411], Fresh[6410], Fresh[6409], Fresh[6408]}), .c ({new_AGEMA_signal_17356, new_AGEMA_signal_17355, new_AGEMA_signal_17354, mcs1_mcs_mat1_7_mcs_rom0_13_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U10 ( .a ({new_AGEMA_signal_14149, new_AGEMA_signal_14148, new_AGEMA_signal_14147, mcs1_mcs_mat1_7_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_11296, new_AGEMA_signal_11295, new_AGEMA_signal_11294, mcs1_mcs_mat1_7_mcs_rom0_14_n11}), .c ({new_AGEMA_signal_15586, new_AGEMA_signal_15585, new_AGEMA_signal_15584, mcs1_mcs_mat1_7_mcs_out[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U9 ( .a ({new_AGEMA_signal_12703, new_AGEMA_signal_12702, new_AGEMA_signal_12701, mcs1_mcs_mat1_7_mcs_rom0_14_n10}), .b ({new_AGEMA_signal_15589, new_AGEMA_signal_15588, new_AGEMA_signal_15587, mcs1_mcs_mat1_7_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_16543, new_AGEMA_signal_16542, new_AGEMA_signal_16541, mcs1_mcs_mat1_7_mcs_out[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U8 ( .a ({new_AGEMA_signal_14149, new_AGEMA_signal_14148, new_AGEMA_signal_14147, mcs1_mcs_mat1_7_mcs_rom0_14_n12}), .b ({new_AGEMA_signal_15589, new_AGEMA_signal_15588, new_AGEMA_signal_15587, mcs1_mcs_mat1_7_mcs_rom0_14_n9}), .c ({new_AGEMA_signal_16546, new_AGEMA_signal_16545, new_AGEMA_signal_16544, mcs1_mcs_mat1_7_mcs_out[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U7 ( .a ({new_AGEMA_signal_11296, new_AGEMA_signal_11295, new_AGEMA_signal_11294, mcs1_mcs_mat1_7_mcs_rom0_14_n11}), .b ({new_AGEMA_signal_14152, new_AGEMA_signal_14151, new_AGEMA_signal_14150, mcs1_mcs_mat1_7_mcs_rom0_14_n8}), .c ({new_AGEMA_signal_15589, new_AGEMA_signal_15588, new_AGEMA_signal_15587, mcs1_mcs_mat1_7_mcs_rom0_14_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U6 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({new_AGEMA_signal_10015, new_AGEMA_signal_10014, new_AGEMA_signal_10013, mcs1_mcs_mat1_7_mcs_rom0_14_x2x4}), .c ({new_AGEMA_signal_11296, new_AGEMA_signal_11295, new_AGEMA_signal_11294, mcs1_mcs_mat1_7_mcs_rom0_14_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U5 ( .a ({new_AGEMA_signal_12700, new_AGEMA_signal_12699, new_AGEMA_signal_12698, mcs1_mcs_mat1_7_mcs_rom0_14_n7}), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .c ({new_AGEMA_signal_14149, new_AGEMA_signal_14148, new_AGEMA_signal_14147, mcs1_mcs_mat1_7_mcs_rom0_14_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U4 ( .a ({new_AGEMA_signal_11299, new_AGEMA_signal_11298, new_AGEMA_signal_11297, mcs1_mcs_mat1_7_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_9103, new_AGEMA_signal_9102, new_AGEMA_signal_9101, mcs1_mcs_mat1_7_mcs_rom0_14_x0x4}), .c ({new_AGEMA_signal_12700, new_AGEMA_signal_12699, new_AGEMA_signal_12698, mcs1_mcs_mat1_7_mcs_rom0_14_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U3 ( .a ({new_AGEMA_signal_14152, new_AGEMA_signal_14151, new_AGEMA_signal_14150, mcs1_mcs_mat1_7_mcs_rom0_14_n8}), .b ({new_AGEMA_signal_12703, new_AGEMA_signal_12702, new_AGEMA_signal_12701, mcs1_mcs_mat1_7_mcs_rom0_14_n10}), .c ({new_AGEMA_signal_15592, new_AGEMA_signal_15591, new_AGEMA_signal_15590, mcs1_mcs_mat1_7_mcs_out[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U2 ( .a ({new_AGEMA_signal_11299, new_AGEMA_signal_11298, new_AGEMA_signal_11297, mcs1_mcs_mat1_7_mcs_rom0_14_x3x4}), .b ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_12703, new_AGEMA_signal_12702, new_AGEMA_signal_12701, mcs1_mcs_mat1_7_mcs_rom0_14_n10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({new_AGEMA_signal_12706, new_AGEMA_signal_12705, new_AGEMA_signal_12704, mcs1_mcs_mat1_7_mcs_rom0_14_x1x4}), .c ({new_AGEMA_signal_14152, new_AGEMA_signal_14151, new_AGEMA_signal_14150, mcs1_mcs_mat1_7_mcs_rom0_14_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6419], Fresh[6418], Fresh[6417], Fresh[6416], Fresh[6415], Fresh[6414]}), .c ({new_AGEMA_signal_12706, new_AGEMA_signal_12705, new_AGEMA_signal_12704, mcs1_mcs_mat1_7_mcs_rom0_14_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6425], Fresh[6424], Fresh[6423], Fresh[6422], Fresh[6421], Fresh[6420]}), .c ({new_AGEMA_signal_10015, new_AGEMA_signal_10014, new_AGEMA_signal_10013, mcs1_mcs_mat1_7_mcs_rom0_14_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_14_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6431], Fresh[6430], Fresh[6429], Fresh[6428], Fresh[6427], Fresh[6426]}), .c ({new_AGEMA_signal_11299, new_AGEMA_signal_11298, new_AGEMA_signal_11297, mcs1_mcs_mat1_7_mcs_rom0_14_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U7 ( .a ({new_AGEMA_signal_15598, new_AGEMA_signal_15597, new_AGEMA_signal_15596, mcs1_mcs_mat1_7_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .c ({new_AGEMA_signal_16549, new_AGEMA_signal_16548, new_AGEMA_signal_16547, mcs1_mcs_mat1_7_mcs_out[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U6 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({new_AGEMA_signal_14155, new_AGEMA_signal_14154, new_AGEMA_signal_14153, mcs1_mcs_mat1_7_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_15595, new_AGEMA_signal_15594, new_AGEMA_signal_15593, mcs1_mcs_mat1_7_mcs_out[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U4 ( .a ({new_AGEMA_signal_16552, new_AGEMA_signal_16551, new_AGEMA_signal_16550, mcs1_mcs_mat1_7_mcs_rom0_15_n5}), .b ({new_AGEMA_signal_11302, new_AGEMA_signal_11301, new_AGEMA_signal_11300, mcs1_mcs_mat1_7_mcs_rom0_15_x3x4}), .c ({new_AGEMA_signal_17359, new_AGEMA_signal_17358, new_AGEMA_signal_17357, mcs1_mcs_mat1_7_mcs_out[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U3 ( .a ({new_AGEMA_signal_15598, new_AGEMA_signal_15597, new_AGEMA_signal_15596, mcs1_mcs_mat1_7_mcs_rom0_15_n7}), .b ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .c ({new_AGEMA_signal_16552, new_AGEMA_signal_16551, new_AGEMA_signal_16550, mcs1_mcs_mat1_7_mcs_rom0_15_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U2 ( .a ({new_AGEMA_signal_10018, new_AGEMA_signal_10017, new_AGEMA_signal_10016, mcs1_mcs_mat1_7_mcs_rom0_15_x2x4}), .b ({new_AGEMA_signal_14155, new_AGEMA_signal_14154, new_AGEMA_signal_14153, mcs1_mcs_mat1_7_mcs_rom0_15_n6}), .c ({new_AGEMA_signal_15598, new_AGEMA_signal_15597, new_AGEMA_signal_15596, mcs1_mcs_mat1_7_mcs_rom0_15_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_U1 ( .a ({new_AGEMA_signal_9106, new_AGEMA_signal_9105, new_AGEMA_signal_9104, mcs1_mcs_mat1_7_mcs_rom0_15_x0x4}), .b ({new_AGEMA_signal_12712, new_AGEMA_signal_12711, new_AGEMA_signal_12710, mcs1_mcs_mat1_7_mcs_rom0_15_x1x4}), .c ({new_AGEMA_signal_14155, new_AGEMA_signal_14154, new_AGEMA_signal_14153, mcs1_mcs_mat1_7_mcs_rom0_15_n6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6437], Fresh[6436], Fresh[6435], Fresh[6434], Fresh[6433], Fresh[6432]}), .c ({new_AGEMA_signal_12712, new_AGEMA_signal_12711, new_AGEMA_signal_12710, mcs1_mcs_mat1_7_mcs_rom0_15_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6443], Fresh[6442], Fresh[6441], Fresh[6440], Fresh[6439], Fresh[6438]}), .c ({new_AGEMA_signal_10018, new_AGEMA_signal_10017, new_AGEMA_signal_10016, mcs1_mcs_mat1_7_mcs_rom0_15_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_15_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6449], Fresh[6448], Fresh[6447], Fresh[6446], Fresh[6445], Fresh[6444]}), .c ({new_AGEMA_signal_11302, new_AGEMA_signal_11301, new_AGEMA_signal_11300, mcs1_mcs_mat1_7_mcs_rom0_15_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U7 ( .a ({new_AGEMA_signal_14164, new_AGEMA_signal_14163, new_AGEMA_signal_14162, mcs1_mcs_mat1_7_mcs_rom0_16_n6}), .b ({new_AGEMA_signal_11305, new_AGEMA_signal_11304, new_AGEMA_signal_11303, mcs1_mcs_mat1_7_mcs_rom0_16_x3x4}), .c ({new_AGEMA_signal_15601, new_AGEMA_signal_15600, new_AGEMA_signal_15599, mcs1_mcs_mat1_7_mcs_out[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U6 ( .a ({new_AGEMA_signal_10021, new_AGEMA_signal_10020, new_AGEMA_signal_10019, mcs1_mcs_mat1_7_mcs_rom0_16_x2x4}), .b ({new_AGEMA_signal_12715, new_AGEMA_signal_12714, new_AGEMA_signal_12713, mcs1_mcs_mat1_7_mcs_rom0_16_n5}), .c ({new_AGEMA_signal_14158, new_AGEMA_signal_14157, new_AGEMA_signal_14156, mcs1_mcs_mat1_7_mcs_out[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_U5 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({new_AGEMA_signal_12718, new_AGEMA_signal_12717, new_AGEMA_signal_12716, mcs1_mcs_mat1_7_mcs_rom0_16_x1x4}), .c ({new_AGEMA_signal_14161, new_AGEMA_signal_14160, new_AGEMA_signal_14159, mcs1_mcs_mat1_7_mcs_out[61]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6455], Fresh[6454], Fresh[6453], Fresh[6452], Fresh[6451], Fresh[6450]}), .c ({new_AGEMA_signal_12718, new_AGEMA_signal_12717, new_AGEMA_signal_12716, mcs1_mcs_mat1_7_mcs_rom0_16_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6461], Fresh[6460], Fresh[6459], Fresh[6458], Fresh[6457], Fresh[6456]}), .c ({new_AGEMA_signal_10021, new_AGEMA_signal_10020, new_AGEMA_signal_10019, mcs1_mcs_mat1_7_mcs_rom0_16_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_16_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6467], Fresh[6466], Fresh[6465], Fresh[6464], Fresh[6463], Fresh[6462]}), .c ({new_AGEMA_signal_11305, new_AGEMA_signal_11304, new_AGEMA_signal_11303, mcs1_mcs_mat1_7_mcs_rom0_16_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U7 ( .a ({new_AGEMA_signal_15610, new_AGEMA_signal_15609, new_AGEMA_signal_15608, mcs1_mcs_mat1_7_mcs_rom0_17_n8}), .b ({new_AGEMA_signal_17362, new_AGEMA_signal_17361, new_AGEMA_signal_17360, mcs1_mcs_mat1_7_mcs_rom0_17_x3x4}), .c ({new_AGEMA_signal_18007, new_AGEMA_signal_18006, new_AGEMA_signal_18005, mcs1_mcs_mat1_7_mcs_out[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U5 ( .a ({new_AGEMA_signal_15613, new_AGEMA_signal_15612, new_AGEMA_signal_15611, mcs1_mcs_mat1_7_mcs_rom0_17_x2x4}), .b ({new_AGEMA_signal_18010, new_AGEMA_signal_18009, new_AGEMA_signal_18008, mcs1_mcs_mat1_7_mcs_rom0_17_n10}), .c ({new_AGEMA_signal_18643, new_AGEMA_signal_18642, new_AGEMA_signal_18641, mcs1_mcs_mat1_7_mcs_out[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U3 ( .a ({new_AGEMA_signal_18646, new_AGEMA_signal_18645, new_AGEMA_signal_18644, mcs1_mcs_mat1_7_mcs_rom0_17_n7}), .b ({new_AGEMA_signal_18013, new_AGEMA_signal_18012, new_AGEMA_signal_18011, mcs1_mcs_mat1_7_mcs_rom0_17_n6}), .c ({new_AGEMA_signal_19318, new_AGEMA_signal_19317, new_AGEMA_signal_19316, mcs1_mcs_mat1_7_mcs_out[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_U1 ( .a ({new_AGEMA_signal_18016, new_AGEMA_signal_18015, new_AGEMA_signal_18014, mcs1_mcs_mat1_7_mcs_rom0_17_x1x4}), .b ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_18646, new_AGEMA_signal_18645, new_AGEMA_signal_18644, mcs1_mcs_mat1_7_mcs_rom0_17_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6473], Fresh[6472], Fresh[6471], Fresh[6470], Fresh[6469], Fresh[6468]}), .c ({new_AGEMA_signal_18016, new_AGEMA_signal_18015, new_AGEMA_signal_18014, mcs1_mcs_mat1_7_mcs_rom0_17_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6479], Fresh[6478], Fresh[6477], Fresh[6476], Fresh[6475], Fresh[6474]}), .c ({new_AGEMA_signal_15613, new_AGEMA_signal_15612, new_AGEMA_signal_15611, mcs1_mcs_mat1_7_mcs_rom0_17_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_17_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6485], Fresh[6484], Fresh[6483], Fresh[6482], Fresh[6481], Fresh[6480]}), .c ({new_AGEMA_signal_17362, new_AGEMA_signal_17361, new_AGEMA_signal_17360, mcs1_mcs_mat1_7_mcs_rom0_17_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U10 ( .a ({new_AGEMA_signal_12724, new_AGEMA_signal_12723, new_AGEMA_signal_12722, mcs1_mcs_mat1_7_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_14170, new_AGEMA_signal_14169, new_AGEMA_signal_14168, mcs1_mcs_mat1_7_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_15616, new_AGEMA_signal_15615, new_AGEMA_signal_15614, mcs1_mcs_mat1_7_mcs_out[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U9 ( .a ({new_AGEMA_signal_15619, new_AGEMA_signal_15618, new_AGEMA_signal_15617, mcs1_mcs_mat1_7_mcs_rom0_18_n11}), .b ({new_AGEMA_signal_12721, new_AGEMA_signal_12720, new_AGEMA_signal_12719, mcs1_mcs_mat1_7_mcs_rom0_18_n10}), .c ({new_AGEMA_signal_16558, new_AGEMA_signal_16557, new_AGEMA_signal_16556, mcs1_mcs_mat1_7_mcs_out[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U8 ( .a ({new_AGEMA_signal_11308, new_AGEMA_signal_11307, new_AGEMA_signal_11306, mcs1_mcs_mat1_7_mcs_rom0_18_x3x4}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_12721, new_AGEMA_signal_12720, new_AGEMA_signal_12719, mcs1_mcs_mat1_7_mcs_rom0_18_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U7 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({new_AGEMA_signal_15619, new_AGEMA_signal_15618, new_AGEMA_signal_15617, mcs1_mcs_mat1_7_mcs_rom0_18_n11}), .c ({new_AGEMA_signal_16561, new_AGEMA_signal_16560, new_AGEMA_signal_16559, mcs1_mcs_mat1_7_mcs_out[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U6 ( .a ({new_AGEMA_signal_9112, new_AGEMA_signal_9111, new_AGEMA_signal_9110, mcs1_mcs_mat1_7_mcs_rom0_18_x0x4}), .b ({new_AGEMA_signal_14170, new_AGEMA_signal_14169, new_AGEMA_signal_14168, mcs1_mcs_mat1_7_mcs_rom0_18_n12}), .c ({new_AGEMA_signal_15619, new_AGEMA_signal_15618, new_AGEMA_signal_15617, mcs1_mcs_mat1_7_mcs_rom0_18_n11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U5 ( .a ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, new_AGEMA_signal_10022, mcs1_mcs_mat1_7_mcs_rom0_18_x2x4}), .b ({new_AGEMA_signal_12730, new_AGEMA_signal_12729, new_AGEMA_signal_12728, mcs1_mcs_mat1_7_mcs_rom0_18_x1x4}), .c ({new_AGEMA_signal_14170, new_AGEMA_signal_14169, new_AGEMA_signal_14168, mcs1_mcs_mat1_7_mcs_rom0_18_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U4 ( .a ({new_AGEMA_signal_12727, new_AGEMA_signal_12726, new_AGEMA_signal_12725, mcs1_mcs_mat1_7_mcs_rom0_18_n9}), .b ({new_AGEMA_signal_14173, new_AGEMA_signal_14172, new_AGEMA_signal_14171, mcs1_mcs_mat1_7_mcs_rom0_18_n8}), .c ({new_AGEMA_signal_15622, new_AGEMA_signal_15621, new_AGEMA_signal_15620, mcs1_mcs_mat1_7_mcs_out[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U3 ( .a ({new_AGEMA_signal_12724, new_AGEMA_signal_12723, new_AGEMA_signal_12722, mcs1_mcs_mat1_7_mcs_rom0_18_n13}), .b ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, new_AGEMA_signal_10022, mcs1_mcs_mat1_7_mcs_rom0_18_x2x4}), .c ({new_AGEMA_signal_14173, new_AGEMA_signal_14172, new_AGEMA_signal_14171, mcs1_mcs_mat1_7_mcs_rom0_18_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_U2 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_11308, new_AGEMA_signal_11307, new_AGEMA_signal_11306, mcs1_mcs_mat1_7_mcs_rom0_18_x3x4}), .c ({new_AGEMA_signal_12724, new_AGEMA_signal_12723, new_AGEMA_signal_12722, mcs1_mcs_mat1_7_mcs_rom0_18_n13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6491], Fresh[6490], Fresh[6489], Fresh[6488], Fresh[6487], Fresh[6486]}), .c ({new_AGEMA_signal_12730, new_AGEMA_signal_12729, new_AGEMA_signal_12728, mcs1_mcs_mat1_7_mcs_rom0_18_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6497], Fresh[6496], Fresh[6495], Fresh[6494], Fresh[6493], Fresh[6492]}), .c ({new_AGEMA_signal_10024, new_AGEMA_signal_10023, new_AGEMA_signal_10022, mcs1_mcs_mat1_7_mcs_rom0_18_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_18_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6503], Fresh[6502], Fresh[6501], Fresh[6500], Fresh[6499], Fresh[6498]}), .c ({new_AGEMA_signal_11308, new_AGEMA_signal_11307, new_AGEMA_signal_11306, mcs1_mcs_mat1_7_mcs_rom0_18_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U5 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_11314, new_AGEMA_signal_11313, new_AGEMA_signal_11312, mcs1_mcs_mat1_7_mcs_rom0_20_x3x4}), .c ({new_AGEMA_signal_12736, new_AGEMA_signal_12735, new_AGEMA_signal_12734, mcs1_mcs_mat1_7_mcs_out[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U4 ( .a ({new_AGEMA_signal_16564, new_AGEMA_signal_16563, new_AGEMA_signal_16562, mcs1_mcs_mat1_7_mcs_rom0_20_n5}), .b ({new_AGEMA_signal_10027, new_AGEMA_signal_10026, new_AGEMA_signal_10025, mcs1_mcs_mat1_7_mcs_rom0_20_x2x4}), .c ({new_AGEMA_signal_17365, new_AGEMA_signal_17364, new_AGEMA_signal_17363, mcs1_mcs_mat1_7_mcs_out[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U3 ( .a ({new_AGEMA_signal_15625, new_AGEMA_signal_15624, new_AGEMA_signal_15623, mcs1_mcs_mat1_7_mcs_out[47]}), .b ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .c ({new_AGEMA_signal_16564, new_AGEMA_signal_16563, new_AGEMA_signal_16562, mcs1_mcs_mat1_7_mcs_rom0_20_n5}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U2 ( .a ({new_AGEMA_signal_14179, new_AGEMA_signal_14178, new_AGEMA_signal_14177, mcs1_mcs_mat1_7_mcs_rom0_20_n4}), .b ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .c ({new_AGEMA_signal_15625, new_AGEMA_signal_15624, new_AGEMA_signal_15623, mcs1_mcs_mat1_7_mcs_out[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_U1 ( .a ({new_AGEMA_signal_9115, new_AGEMA_signal_9114, new_AGEMA_signal_9113, mcs1_mcs_mat1_7_mcs_rom0_20_x0x4}), .b ({new_AGEMA_signal_12739, new_AGEMA_signal_12738, new_AGEMA_signal_12737, mcs1_mcs_mat1_7_mcs_rom0_20_x1x4}), .c ({new_AGEMA_signal_14179, new_AGEMA_signal_14178, new_AGEMA_signal_14177, mcs1_mcs_mat1_7_mcs_rom0_20_n4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6509], Fresh[6508], Fresh[6507], Fresh[6506], Fresh[6505], Fresh[6504]}), .c ({new_AGEMA_signal_12739, new_AGEMA_signal_12738, new_AGEMA_signal_12737, mcs1_mcs_mat1_7_mcs_rom0_20_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6515], Fresh[6514], Fresh[6513], Fresh[6512], Fresh[6511], Fresh[6510]}), .c ({new_AGEMA_signal_10027, new_AGEMA_signal_10026, new_AGEMA_signal_10025, mcs1_mcs_mat1_7_mcs_rom0_20_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_20_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6521], Fresh[6520], Fresh[6519], Fresh[6518], Fresh[6517], Fresh[6516]}), .c ({new_AGEMA_signal_11314, new_AGEMA_signal_11313, new_AGEMA_signal_11312, mcs1_mcs_mat1_7_mcs_rom0_20_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U10 ( .a ({new_AGEMA_signal_18649, new_AGEMA_signal_18648, new_AGEMA_signal_18647, mcs1_mcs_mat1_7_mcs_rom0_21_n12}), .b ({new_AGEMA_signal_17368, new_AGEMA_signal_17367, new_AGEMA_signal_17366, mcs1_mcs_mat1_7_mcs_rom0_21_n11}), .c ({new_AGEMA_signal_19321, new_AGEMA_signal_19320, new_AGEMA_signal_19319, mcs1_mcs_mat1_7_mcs_out[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U9 ( .a ({new_AGEMA_signal_18019, new_AGEMA_signal_18018, new_AGEMA_signal_18017, mcs1_mcs_mat1_7_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_15628, new_AGEMA_signal_15627, new_AGEMA_signal_15626, mcs1_mcs_mat1_7_mcs_rom0_21_x2x4}), .c ({new_AGEMA_signal_18649, new_AGEMA_signal_18648, new_AGEMA_signal_18647, mcs1_mcs_mat1_7_mcs_rom0_21_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U8 ( .a ({new_AGEMA_signal_18652, new_AGEMA_signal_18651, new_AGEMA_signal_18650, mcs1_mcs_mat1_7_mcs_rom0_21_n9}), .b ({new_AGEMA_signal_18025, new_AGEMA_signal_18024, new_AGEMA_signal_18023, mcs1_mcs_mat1_7_mcs_rom0_21_x1x4}), .c ({new_AGEMA_signal_19324, new_AGEMA_signal_19323, new_AGEMA_signal_19322, mcs1_mcs_mat1_7_mcs_out[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U6 ( .a ({new_AGEMA_signal_18655, new_AGEMA_signal_18654, new_AGEMA_signal_18653, mcs1_mcs_mat1_7_mcs_rom0_21_n8}), .b ({new_AGEMA_signal_14182, new_AGEMA_signal_14181, new_AGEMA_signal_14180, mcs1_mcs_mat1_7_mcs_rom0_21_x0x4}), .c ({new_AGEMA_signal_19327, new_AGEMA_signal_19326, new_AGEMA_signal_19325, mcs1_mcs_mat1_7_mcs_out[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U5 ( .a ({new_AGEMA_signal_18019, new_AGEMA_signal_18018, new_AGEMA_signal_18017, mcs1_mcs_mat1_7_mcs_rom0_21_n10}), .b ({new_AGEMA_signal_17371, new_AGEMA_signal_17370, new_AGEMA_signal_17369, mcs1_mcs_mat1_7_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_18655, new_AGEMA_signal_18654, new_AGEMA_signal_18653, mcs1_mcs_mat1_7_mcs_rom0_21_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_U3 ( .a ({new_AGEMA_signal_18022, new_AGEMA_signal_18021, new_AGEMA_signal_18020, mcs1_mcs_mat1_7_mcs_rom0_21_n7}), .b ({new_AGEMA_signal_17371, new_AGEMA_signal_17370, new_AGEMA_signal_17369, mcs1_mcs_mat1_7_mcs_rom0_21_x3x4}), .c ({new_AGEMA_signal_18658, new_AGEMA_signal_18657, new_AGEMA_signal_18656, mcs1_mcs_mat1_7_mcs_out[40]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6527], Fresh[6526], Fresh[6525], Fresh[6524], Fresh[6523], Fresh[6522]}), .c ({new_AGEMA_signal_18025, new_AGEMA_signal_18024, new_AGEMA_signal_18023, mcs1_mcs_mat1_7_mcs_rom0_21_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6533], Fresh[6532], Fresh[6531], Fresh[6530], Fresh[6529], Fresh[6528]}), .c ({new_AGEMA_signal_15628, new_AGEMA_signal_15627, new_AGEMA_signal_15626, mcs1_mcs_mat1_7_mcs_rom0_21_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_21_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6539], Fresh[6538], Fresh[6537], Fresh[6536], Fresh[6535], Fresh[6534]}), .c ({new_AGEMA_signal_17371, new_AGEMA_signal_17370, new_AGEMA_signal_17369, mcs1_mcs_mat1_7_mcs_rom0_21_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U10 ( .a ({new_AGEMA_signal_15631, new_AGEMA_signal_15630, new_AGEMA_signal_15629, mcs1_mcs_mat1_7_mcs_rom0_22_n13}), .b ({new_AGEMA_signal_9118, new_AGEMA_signal_9117, new_AGEMA_signal_9116, mcs1_mcs_mat1_7_mcs_rom0_22_x0x4}), .c ({new_AGEMA_signal_16567, new_AGEMA_signal_16566, new_AGEMA_signal_16565, mcs1_mcs_mat1_7_mcs_out[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U9 ( .a ({new_AGEMA_signal_11320, new_AGEMA_signal_11319, new_AGEMA_signal_11318, mcs1_mcs_mat1_7_mcs_rom0_22_n12}), .b ({new_AGEMA_signal_11317, new_AGEMA_signal_11316, new_AGEMA_signal_11315, mcs1_mcs_mat1_7_mcs_rom0_22_n11}), .c ({new_AGEMA_signal_12742, new_AGEMA_signal_12741, new_AGEMA_signal_12740, mcs1_mcs_mat1_7_mcs_out[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U7 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({new_AGEMA_signal_15631, new_AGEMA_signal_15630, new_AGEMA_signal_15629, mcs1_mcs_mat1_7_mcs_rom0_22_n13}), .c ({new_AGEMA_signal_16570, new_AGEMA_signal_16569, new_AGEMA_signal_16568, mcs1_mcs_mat1_7_mcs_out[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U6 ( .a ({new_AGEMA_signal_12745, new_AGEMA_signal_12744, new_AGEMA_signal_12743, mcs1_mcs_mat1_7_mcs_rom0_22_n10}), .b ({new_AGEMA_signal_14185, new_AGEMA_signal_14184, new_AGEMA_signal_14183, mcs1_mcs_mat1_7_mcs_rom0_22_n9}), .c ({new_AGEMA_signal_15631, new_AGEMA_signal_15630, new_AGEMA_signal_15629, mcs1_mcs_mat1_7_mcs_rom0_22_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U5 ( .a ({new_AGEMA_signal_12748, new_AGEMA_signal_12747, new_AGEMA_signal_12746, mcs1_mcs_mat1_7_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_11323, new_AGEMA_signal_11322, new_AGEMA_signal_11321, mcs1_mcs_mat1_7_mcs_rom0_22_x3x4}), .c ({new_AGEMA_signal_14185, new_AGEMA_signal_14184, new_AGEMA_signal_14183, mcs1_mcs_mat1_7_mcs_rom0_22_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U3 ( .a ({new_AGEMA_signal_12748, new_AGEMA_signal_12747, new_AGEMA_signal_12746, mcs1_mcs_mat1_7_mcs_rom0_22_x1x4}), .b ({new_AGEMA_signal_11320, new_AGEMA_signal_11319, new_AGEMA_signal_11318, mcs1_mcs_mat1_7_mcs_rom0_22_n12}), .c ({new_AGEMA_signal_14188, new_AGEMA_signal_14187, new_AGEMA_signal_14186, mcs1_mcs_mat1_7_mcs_out[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U2 ( .a ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .b ({new_AGEMA_signal_10357, new_AGEMA_signal_10356, new_AGEMA_signal_10355, mcs1_mcs_mat1_7_mcs_rom0_22_n8}), .c ({new_AGEMA_signal_11320, new_AGEMA_signal_11319, new_AGEMA_signal_11318, mcs1_mcs_mat1_7_mcs_rom0_22_n12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({new_AGEMA_signal_10030, new_AGEMA_signal_10029, new_AGEMA_signal_10028, mcs1_mcs_mat1_7_mcs_rom0_22_x2x4}), .c ({new_AGEMA_signal_10357, new_AGEMA_signal_10356, new_AGEMA_signal_10355, mcs1_mcs_mat1_7_mcs_rom0_22_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6545], Fresh[6544], Fresh[6543], Fresh[6542], Fresh[6541], Fresh[6540]}), .c ({new_AGEMA_signal_12748, new_AGEMA_signal_12747, new_AGEMA_signal_12746, mcs1_mcs_mat1_7_mcs_rom0_22_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6551], Fresh[6550], Fresh[6549], Fresh[6548], Fresh[6547], Fresh[6546]}), .c ({new_AGEMA_signal_10030, new_AGEMA_signal_10029, new_AGEMA_signal_10028, mcs1_mcs_mat1_7_mcs_rom0_22_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_22_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6557], Fresh[6556], Fresh[6555], Fresh[6554], Fresh[6553], Fresh[6552]}), .c ({new_AGEMA_signal_11323, new_AGEMA_signal_11322, new_AGEMA_signal_11321, mcs1_mcs_mat1_7_mcs_rom0_22_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U7 ( .a ({new_AGEMA_signal_12751, new_AGEMA_signal_12750, new_AGEMA_signal_12749, mcs1_mcs_mat1_7_mcs_rom0_23_n6}), .b ({new_AGEMA_signal_11326, new_AGEMA_signal_11325, new_AGEMA_signal_11324, mcs1_mcs_mat1_7_mcs_rom0_23_x3x4}), .c ({new_AGEMA_signal_14191, new_AGEMA_signal_14190, new_AGEMA_signal_14189, mcs1_mcs_mat1_7_mcs_out[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U6 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_10033, new_AGEMA_signal_10032, new_AGEMA_signal_10031, mcs1_mcs_mat1_7_mcs_rom0_23_x2x4}), .c ({new_AGEMA_signal_10360, new_AGEMA_signal_10359, new_AGEMA_signal_10358, mcs1_mcs_mat1_7_mcs_out[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_U5 ( .a ({new_AGEMA_signal_16573, new_AGEMA_signal_16572, new_AGEMA_signal_16571, mcs1_mcs_mat1_7_mcs_rom0_23_n5}), .b ({new_AGEMA_signal_12754, new_AGEMA_signal_12753, new_AGEMA_signal_12752, mcs1_mcs_mat1_7_mcs_rom0_23_x1x4}), .c ({new_AGEMA_signal_17374, new_AGEMA_signal_17373, new_AGEMA_signal_17372, mcs1_mcs_mat1_7_mcs_out[32]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6563], Fresh[6562], Fresh[6561], Fresh[6560], Fresh[6559], Fresh[6558]}), .c ({new_AGEMA_signal_12754, new_AGEMA_signal_12753, new_AGEMA_signal_12752, mcs1_mcs_mat1_7_mcs_rom0_23_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6569], Fresh[6568], Fresh[6567], Fresh[6566], Fresh[6565], Fresh[6564]}), .c ({new_AGEMA_signal_10033, new_AGEMA_signal_10032, new_AGEMA_signal_10031, mcs1_mcs_mat1_7_mcs_rom0_23_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_23_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6575], Fresh[6574], Fresh[6573], Fresh[6572], Fresh[6571], Fresh[6570]}), .c ({new_AGEMA_signal_11326, new_AGEMA_signal_11325, new_AGEMA_signal_11324, mcs1_mcs_mat1_7_mcs_rom0_23_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U11 ( .a ({new_AGEMA_signal_15637, new_AGEMA_signal_15636, new_AGEMA_signal_15635, mcs1_mcs_mat1_7_mcs_rom0_24_n15}), .b ({new_AGEMA_signal_14197, new_AGEMA_signal_14196, new_AGEMA_signal_14195, mcs1_mcs_mat1_7_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_16576, new_AGEMA_signal_16575, new_AGEMA_signal_16574, mcs1_mcs_mat1_7_mcs_out[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U10 ( .a ({new_AGEMA_signal_10039, new_AGEMA_signal_10038, new_AGEMA_signal_10037, mcs1_mcs_mat1_7_mcs_rom0_24_x2x4}), .b ({new_AGEMA_signal_14200, new_AGEMA_signal_14199, new_AGEMA_signal_14198, mcs1_mcs_mat1_7_mcs_out[29]}), .c ({new_AGEMA_signal_15637, new_AGEMA_signal_15636, new_AGEMA_signal_15635, mcs1_mcs_mat1_7_mcs_rom0_24_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U9 ( .a ({new_AGEMA_signal_10036, new_AGEMA_signal_10035, new_AGEMA_signal_10034, mcs1_mcs_mat1_7_mcs_rom0_24_n13}), .b ({new_AGEMA_signal_14197, new_AGEMA_signal_14196, new_AGEMA_signal_14195, mcs1_mcs_mat1_7_mcs_rom0_24_n14}), .c ({new_AGEMA_signal_15640, new_AGEMA_signal_15639, new_AGEMA_signal_15638, mcs1_mcs_mat1_7_mcs_out[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U8 ( .a ({new_AGEMA_signal_12763, new_AGEMA_signal_12762, new_AGEMA_signal_12761, mcs1_mcs_mat1_7_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .c ({new_AGEMA_signal_14197, new_AGEMA_signal_14196, new_AGEMA_signal_14195, mcs1_mcs_mat1_7_mcs_rom0_24_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U5 ( .a ({new_AGEMA_signal_15643, new_AGEMA_signal_15642, new_AGEMA_signal_15641, mcs1_mcs_mat1_7_mcs_rom0_24_n11}), .b ({new_AGEMA_signal_12757, new_AGEMA_signal_12756, new_AGEMA_signal_12755, mcs1_mcs_mat1_7_mcs_rom0_24_n12}), .c ({new_AGEMA_signal_16579, new_AGEMA_signal_16578, new_AGEMA_signal_16577, mcs1_mcs_mat1_7_mcs_out[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U3 ( .a ({new_AGEMA_signal_14203, new_AGEMA_signal_14202, new_AGEMA_signal_14201, mcs1_mcs_mat1_7_mcs_rom0_24_n10}), .b ({new_AGEMA_signal_12760, new_AGEMA_signal_12759, new_AGEMA_signal_12758, mcs1_mcs_mat1_7_mcs_rom0_24_n9}), .c ({new_AGEMA_signal_15643, new_AGEMA_signal_15642, new_AGEMA_signal_15641, mcs1_mcs_mat1_7_mcs_rom0_24_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U2 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_11329, new_AGEMA_signal_11328, new_AGEMA_signal_11327, mcs1_mcs_mat1_7_mcs_rom0_24_x3x4}), .c ({new_AGEMA_signal_12760, new_AGEMA_signal_12759, new_AGEMA_signal_12758, mcs1_mcs_mat1_7_mcs_rom0_24_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_U1 ( .a ({new_AGEMA_signal_12763, new_AGEMA_signal_12762, new_AGEMA_signal_12761, mcs1_mcs_mat1_7_mcs_rom0_24_x1x4}), .b ({new_AGEMA_signal_10039, new_AGEMA_signal_10038, new_AGEMA_signal_10037, mcs1_mcs_mat1_7_mcs_rom0_24_x2x4}), .c ({new_AGEMA_signal_14203, new_AGEMA_signal_14202, new_AGEMA_signal_14201, mcs1_mcs_mat1_7_mcs_rom0_24_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6581], Fresh[6580], Fresh[6579], Fresh[6578], Fresh[6577], Fresh[6576]}), .c ({new_AGEMA_signal_12763, new_AGEMA_signal_12762, new_AGEMA_signal_12761, mcs1_mcs_mat1_7_mcs_rom0_24_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6587], Fresh[6586], Fresh[6585], Fresh[6584], Fresh[6583], Fresh[6582]}), .c ({new_AGEMA_signal_10039, new_AGEMA_signal_10038, new_AGEMA_signal_10037, mcs1_mcs_mat1_7_mcs_rom0_24_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_24_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6593], Fresh[6592], Fresh[6591], Fresh[6590], Fresh[6589], Fresh[6588]}), .c ({new_AGEMA_signal_11329, new_AGEMA_signal_11328, new_AGEMA_signal_11327, mcs1_mcs_mat1_7_mcs_rom0_24_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U8 ( .a ({new_AGEMA_signal_18028, new_AGEMA_signal_18027, new_AGEMA_signal_18026, mcs1_mcs_mat1_7_mcs_rom0_25_n8}), .b ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_18661, new_AGEMA_signal_18660, new_AGEMA_signal_18659, mcs1_mcs_mat1_7_mcs_out[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U7 ( .a ({new_AGEMA_signal_17377, new_AGEMA_signal_17376, new_AGEMA_signal_17375, mcs1_mcs_mat1_7_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_15646, new_AGEMA_signal_15645, new_AGEMA_signal_15644, mcs1_mcs_mat1_7_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_18028, new_AGEMA_signal_18027, new_AGEMA_signal_18026, mcs1_mcs_mat1_7_mcs_rom0_25_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U6 ( .a ({new_AGEMA_signal_18664, new_AGEMA_signal_18663, new_AGEMA_signal_18662, mcs1_mcs_mat1_7_mcs_rom0_25_n7}), .b ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_19330, new_AGEMA_signal_19329, new_AGEMA_signal_19328, mcs1_mcs_mat1_7_mcs_out[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U5 ( .a ({new_AGEMA_signal_18034, new_AGEMA_signal_18033, new_AGEMA_signal_18032, mcs1_mcs_mat1_7_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_15646, new_AGEMA_signal_15645, new_AGEMA_signal_15644, mcs1_mcs_mat1_7_mcs_rom0_25_x2x4}), .c ({new_AGEMA_signal_18664, new_AGEMA_signal_18663, new_AGEMA_signal_18662, mcs1_mcs_mat1_7_mcs_rom0_25_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U4 ( .a ({new_AGEMA_signal_19333, new_AGEMA_signal_19332, new_AGEMA_signal_19331, mcs1_mcs_mat1_7_mcs_rom0_25_n6}), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .c ({new_AGEMA_signal_20038, new_AGEMA_signal_20037, new_AGEMA_signal_20036, mcs1_mcs_mat1_7_mcs_out[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U3 ( .a ({new_AGEMA_signal_18034, new_AGEMA_signal_18033, new_AGEMA_signal_18032, mcs1_mcs_mat1_7_mcs_rom0_25_x1x4}), .b ({new_AGEMA_signal_18667, new_AGEMA_signal_18666, new_AGEMA_signal_18665, mcs1_mcs_mat1_7_mcs_out[24]}), .c ({new_AGEMA_signal_19333, new_AGEMA_signal_19332, new_AGEMA_signal_19331, mcs1_mcs_mat1_7_mcs_rom0_25_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U2 ( .a ({new_AGEMA_signal_18031, new_AGEMA_signal_18030, new_AGEMA_signal_18029, mcs1_mcs_mat1_7_mcs_rom0_25_n5}), .b ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .c ({new_AGEMA_signal_18667, new_AGEMA_signal_18666, new_AGEMA_signal_18665, mcs1_mcs_mat1_7_mcs_out[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_U1 ( .a ({new_AGEMA_signal_17377, new_AGEMA_signal_17376, new_AGEMA_signal_17375, mcs1_mcs_mat1_7_mcs_rom0_25_x3x4}), .b ({new_AGEMA_signal_14206, new_AGEMA_signal_14205, new_AGEMA_signal_14204, mcs1_mcs_mat1_7_mcs_rom0_25_x0x4}), .c ({new_AGEMA_signal_18031, new_AGEMA_signal_18030, new_AGEMA_signal_18029, mcs1_mcs_mat1_7_mcs_rom0_25_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6599], Fresh[6598], Fresh[6597], Fresh[6596], Fresh[6595], Fresh[6594]}), .c ({new_AGEMA_signal_18034, new_AGEMA_signal_18033, new_AGEMA_signal_18032, mcs1_mcs_mat1_7_mcs_rom0_25_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6605], Fresh[6604], Fresh[6603], Fresh[6602], Fresh[6601], Fresh[6600]}), .c ({new_AGEMA_signal_15646, new_AGEMA_signal_15645, new_AGEMA_signal_15644, mcs1_mcs_mat1_7_mcs_rom0_25_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_25_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6611], Fresh[6610], Fresh[6609], Fresh[6608], Fresh[6607], Fresh[6606]}), .c ({new_AGEMA_signal_17377, new_AGEMA_signal_17376, new_AGEMA_signal_17375, mcs1_mcs_mat1_7_mcs_rom0_25_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U8 ( .a ({new_AGEMA_signal_12766, new_AGEMA_signal_12765, new_AGEMA_signal_12764, mcs1_mcs_mat1_7_mcs_rom0_26_n8}), .b ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .c ({new_AGEMA_signal_14209, new_AGEMA_signal_14208, new_AGEMA_signal_14207, mcs1_mcs_mat1_7_mcs_out[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U7 ( .a ({new_AGEMA_signal_11332, new_AGEMA_signal_11331, new_AGEMA_signal_11330, mcs1_mcs_mat1_7_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_10042, new_AGEMA_signal_10041, new_AGEMA_signal_10040, mcs1_mcs_mat1_7_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_12766, new_AGEMA_signal_12765, new_AGEMA_signal_12764, mcs1_mcs_mat1_7_mcs_rom0_26_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U6 ( .a ({new_AGEMA_signal_14212, new_AGEMA_signal_14211, new_AGEMA_signal_14210, mcs1_mcs_mat1_7_mcs_rom0_26_n7}), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .c ({new_AGEMA_signal_15649, new_AGEMA_signal_15648, new_AGEMA_signal_15647, mcs1_mcs_mat1_7_mcs_out[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U5 ( .a ({new_AGEMA_signal_12772, new_AGEMA_signal_12771, new_AGEMA_signal_12770, mcs1_mcs_mat1_7_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_10042, new_AGEMA_signal_10041, new_AGEMA_signal_10040, mcs1_mcs_mat1_7_mcs_rom0_26_x2x4}), .c ({new_AGEMA_signal_14212, new_AGEMA_signal_14211, new_AGEMA_signal_14210, mcs1_mcs_mat1_7_mcs_rom0_26_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U4 ( .a ({new_AGEMA_signal_15652, new_AGEMA_signal_15651, new_AGEMA_signal_15650, mcs1_mcs_mat1_7_mcs_rom0_26_n6}), .b ({new_AGEMA_signal_8398, new_AGEMA_signal_8397, new_AGEMA_signal_8396, mcs1_mcs_mat1_7_mcs_out[86]}), .c ({new_AGEMA_signal_16582, new_AGEMA_signal_16581, new_AGEMA_signal_16580, mcs1_mcs_mat1_7_mcs_out[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U3 ( .a ({new_AGEMA_signal_12772, new_AGEMA_signal_12771, new_AGEMA_signal_12770, mcs1_mcs_mat1_7_mcs_rom0_26_x1x4}), .b ({new_AGEMA_signal_14215, new_AGEMA_signal_14214, new_AGEMA_signal_14213, mcs1_mcs_mat1_7_mcs_out[20]}), .c ({new_AGEMA_signal_15652, new_AGEMA_signal_15651, new_AGEMA_signal_15650, mcs1_mcs_mat1_7_mcs_rom0_26_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U2 ( .a ({new_AGEMA_signal_12769, new_AGEMA_signal_12768, new_AGEMA_signal_12767, mcs1_mcs_mat1_7_mcs_rom0_26_n5}), .b ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .c ({new_AGEMA_signal_14215, new_AGEMA_signal_14214, new_AGEMA_signal_14213, mcs1_mcs_mat1_7_mcs_out[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_U1 ( .a ({new_AGEMA_signal_11332, new_AGEMA_signal_11331, new_AGEMA_signal_11330, mcs1_mcs_mat1_7_mcs_rom0_26_x3x4}), .b ({new_AGEMA_signal_9127, new_AGEMA_signal_9126, new_AGEMA_signal_9125, mcs1_mcs_mat1_7_mcs_rom0_26_x0x4}), .c ({new_AGEMA_signal_12769, new_AGEMA_signal_12768, new_AGEMA_signal_12767, mcs1_mcs_mat1_7_mcs_rom0_26_n5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6617], Fresh[6616], Fresh[6615], Fresh[6614], Fresh[6613], Fresh[6612]}), .c ({new_AGEMA_signal_12772, new_AGEMA_signal_12771, new_AGEMA_signal_12770, mcs1_mcs_mat1_7_mcs_rom0_26_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6623], Fresh[6622], Fresh[6621], Fresh[6620], Fresh[6619], Fresh[6618]}), .c ({new_AGEMA_signal_10042, new_AGEMA_signal_10041, new_AGEMA_signal_10040, mcs1_mcs_mat1_7_mcs_rom0_26_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_26_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6629], Fresh[6628], Fresh[6627], Fresh[6626], Fresh[6625], Fresh[6624]}), .c ({new_AGEMA_signal_11332, new_AGEMA_signal_11331, new_AGEMA_signal_11330, mcs1_mcs_mat1_7_mcs_rom0_26_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U10 ( .a ({new_AGEMA_signal_12775, new_AGEMA_signal_12774, new_AGEMA_signal_12773, mcs1_mcs_mat1_7_mcs_rom0_27_n12}), .b ({new_AGEMA_signal_12784, new_AGEMA_signal_12783, new_AGEMA_signal_12782, mcs1_mcs_mat1_7_mcs_rom0_27_x1x4}), .c ({new_AGEMA_signal_14218, new_AGEMA_signal_14217, new_AGEMA_signal_14216, mcs1_mcs_mat1_7_mcs_out[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U8 ( .a ({new_AGEMA_signal_14221, new_AGEMA_signal_14220, new_AGEMA_signal_14219, mcs1_mcs_mat1_7_mcs_rom0_27_n10}), .b ({new_AGEMA_signal_9130, new_AGEMA_signal_9129, new_AGEMA_signal_9128, mcs1_mcs_mat1_7_mcs_rom0_27_x0x4}), .c ({new_AGEMA_signal_15655, new_AGEMA_signal_15654, new_AGEMA_signal_15653, mcs1_mcs_mat1_7_mcs_out[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U7 ( .a ({new_AGEMA_signal_15658, new_AGEMA_signal_15657, new_AGEMA_signal_15656, mcs1_mcs_mat1_7_mcs_rom0_27_n9}), .b ({new_AGEMA_signal_10045, new_AGEMA_signal_10044, new_AGEMA_signal_10043, mcs1_mcs_mat1_7_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_16585, new_AGEMA_signal_16584, new_AGEMA_signal_16583, mcs1_mcs_mat1_7_mcs_out[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U6 ( .a ({new_AGEMA_signal_8416, new_AGEMA_signal_8415, new_AGEMA_signal_8414, mcs1_mcs_mat1_7_mcs_out[50]}), .b ({new_AGEMA_signal_14221, new_AGEMA_signal_14220, new_AGEMA_signal_14219, mcs1_mcs_mat1_7_mcs_rom0_27_n10}), .c ({new_AGEMA_signal_15658, new_AGEMA_signal_15657, new_AGEMA_signal_15656, mcs1_mcs_mat1_7_mcs_rom0_27_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U5 ( .a ({new_AGEMA_signal_12778, new_AGEMA_signal_12777, new_AGEMA_signal_12776, mcs1_mcs_mat1_7_mcs_rom0_27_n8}), .b ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .c ({new_AGEMA_signal_14221, new_AGEMA_signal_14220, new_AGEMA_signal_14219, mcs1_mcs_mat1_7_mcs_rom0_27_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U4 ( .a ({new_AGEMA_signal_11335, new_AGEMA_signal_11334, new_AGEMA_signal_11333, mcs1_mcs_mat1_7_mcs_rom0_27_n11}), .b ({new_AGEMA_signal_11338, new_AGEMA_signal_11337, new_AGEMA_signal_11336, mcs1_mcs_mat1_7_mcs_rom0_27_x3x4}), .c ({new_AGEMA_signal_12778, new_AGEMA_signal_12777, new_AGEMA_signal_12776, mcs1_mcs_mat1_7_mcs_rom0_27_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_U2 ( .a ({new_AGEMA_signal_12781, new_AGEMA_signal_12780, new_AGEMA_signal_12779, mcs1_mcs_mat1_7_mcs_rom0_27_n7}), .b ({new_AGEMA_signal_10045, new_AGEMA_signal_10044, new_AGEMA_signal_10043, mcs1_mcs_mat1_7_mcs_rom0_27_x2x4}), .c ({new_AGEMA_signal_14224, new_AGEMA_signal_14223, new_AGEMA_signal_14222, mcs1_mcs_mat1_7_mcs_out[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6635], Fresh[6634], Fresh[6633], Fresh[6632], Fresh[6631], Fresh[6630]}), .c ({new_AGEMA_signal_12784, new_AGEMA_signal_12783, new_AGEMA_signal_12782, mcs1_mcs_mat1_7_mcs_rom0_27_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6641], Fresh[6640], Fresh[6639], Fresh[6638], Fresh[6637], Fresh[6636]}), .c ({new_AGEMA_signal_10045, new_AGEMA_signal_10044, new_AGEMA_signal_10043, mcs1_mcs_mat1_7_mcs_rom0_27_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_27_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6647], Fresh[6646], Fresh[6645], Fresh[6644], Fresh[6643], Fresh[6642]}), .c ({new_AGEMA_signal_11338, new_AGEMA_signal_11337, new_AGEMA_signal_11336, mcs1_mcs_mat1_7_mcs_rom0_27_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U11 ( .a ({new_AGEMA_signal_15667, new_AGEMA_signal_15666, new_AGEMA_signal_15665, mcs1_mcs_mat1_7_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_10363, new_AGEMA_signal_10362, new_AGEMA_signal_10361, mcs1_mcs_mat1_7_mcs_rom0_28_n14}), .c ({new_AGEMA_signal_16588, new_AGEMA_signal_16587, new_AGEMA_signal_16586, mcs1_mcs_mat1_7_mcs_out[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U10 ( .a ({new_AGEMA_signal_14233, new_AGEMA_signal_14232, new_AGEMA_signal_14231, mcs1_mcs_mat1_7_mcs_rom0_28_n13}), .b ({new_AGEMA_signal_14227, new_AGEMA_signal_14226, new_AGEMA_signal_14225, mcs1_mcs_mat1_7_mcs_rom0_28_n12}), .c ({new_AGEMA_signal_15661, new_AGEMA_signal_15660, new_AGEMA_signal_15659, mcs1_mcs_mat1_7_mcs_out[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U9 ( .a ({new_AGEMA_signal_12790, new_AGEMA_signal_12789, new_AGEMA_signal_12788, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}), .b ({new_AGEMA_signal_10048, new_AGEMA_signal_10047, new_AGEMA_signal_10046, mcs1_mcs_mat1_7_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_14227, new_AGEMA_signal_14226, new_AGEMA_signal_14225, mcs1_mcs_mat1_7_mcs_rom0_28_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U8 ( .a ({new_AGEMA_signal_10363, new_AGEMA_signal_10362, new_AGEMA_signal_10361, mcs1_mcs_mat1_7_mcs_rom0_28_n14}), .b ({new_AGEMA_signal_14230, new_AGEMA_signal_14229, new_AGEMA_signal_14228, mcs1_mcs_mat1_7_mcs_rom0_28_n11}), .c ({new_AGEMA_signal_15664, new_AGEMA_signal_15663, new_AGEMA_signal_15662, mcs1_mcs_mat1_7_mcs_out[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U7 ( .a ({new_AGEMA_signal_12787, new_AGEMA_signal_12786, new_AGEMA_signal_12785, mcs1_mcs_mat1_7_mcs_rom0_28_n10}), .b ({new_AGEMA_signal_12790, new_AGEMA_signal_12789, new_AGEMA_signal_12788, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_14230, new_AGEMA_signal_14229, new_AGEMA_signal_14228, mcs1_mcs_mat1_7_mcs_rom0_28_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U6 ( .a ({new_AGEMA_signal_9133, new_AGEMA_signal_9132, new_AGEMA_signal_9131, mcs1_mcs_mat1_7_mcs_rom0_28_x0x4}), .b ({new_AGEMA_signal_10048, new_AGEMA_signal_10047, new_AGEMA_signal_10046, mcs1_mcs_mat1_7_mcs_rom0_28_x2x4}), .c ({new_AGEMA_signal_10363, new_AGEMA_signal_10362, new_AGEMA_signal_10361, mcs1_mcs_mat1_7_mcs_rom0_28_n14}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U5 ( .a ({new_AGEMA_signal_16591, new_AGEMA_signal_16590, new_AGEMA_signal_16589, mcs1_mcs_mat1_7_mcs_rom0_28_n9}), .b ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .c ({new_AGEMA_signal_17380, new_AGEMA_signal_17379, new_AGEMA_signal_17378, mcs1_mcs_mat1_7_mcs_out[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U4 ( .a ({new_AGEMA_signal_15667, new_AGEMA_signal_15666, new_AGEMA_signal_15665, mcs1_mcs_mat1_7_mcs_rom0_28_n15}), .b ({new_AGEMA_signal_12790, new_AGEMA_signal_12789, new_AGEMA_signal_12788, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}), .c ({new_AGEMA_signal_16591, new_AGEMA_signal_16590, new_AGEMA_signal_16589, mcs1_mcs_mat1_7_mcs_rom0_28_n9}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U3 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({new_AGEMA_signal_14233, new_AGEMA_signal_14232, new_AGEMA_signal_14231, mcs1_mcs_mat1_7_mcs_rom0_28_n13}), .c ({new_AGEMA_signal_15667, new_AGEMA_signal_15666, new_AGEMA_signal_15665, mcs1_mcs_mat1_7_mcs_rom0_28_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U2 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({new_AGEMA_signal_12787, new_AGEMA_signal_12786, new_AGEMA_signal_12785, mcs1_mcs_mat1_7_mcs_rom0_28_n10}), .c ({new_AGEMA_signal_14233, new_AGEMA_signal_14232, new_AGEMA_signal_14231, mcs1_mcs_mat1_7_mcs_rom0_28_n13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_U1 ( .a ({new_AGEMA_signal_8362, new_AGEMA_signal_8361, new_AGEMA_signal_8360, shiftr_out[96]}), .b ({new_AGEMA_signal_11341, new_AGEMA_signal_11340, new_AGEMA_signal_11339, mcs1_mcs_mat1_7_mcs_rom0_28_x3x4}), .c ({new_AGEMA_signal_12787, new_AGEMA_signal_12786, new_AGEMA_signal_12785, mcs1_mcs_mat1_7_mcs_rom0_28_n10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10401, new_AGEMA_signal_10400, mcs1_mcs_mat1_7_mcs_out[126]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6653], Fresh[6652], Fresh[6651], Fresh[6650], Fresh[6649], Fresh[6648]}), .c ({new_AGEMA_signal_12790, new_AGEMA_signal_12789, new_AGEMA_signal_12788, mcs1_mcs_mat1_7_mcs_rom0_28_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8566, new_AGEMA_signal_8565, new_AGEMA_signal_8564, mcs1_mcs_mat1_7_mcs_out[127]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6659], Fresh[6658], Fresh[6657], Fresh[6656], Fresh[6655], Fresh[6654]}), .c ({new_AGEMA_signal_10048, new_AGEMA_signal_10047, new_AGEMA_signal_10046, mcs1_mcs_mat1_7_mcs_rom0_28_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_28_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10204, new_AGEMA_signal_10203, new_AGEMA_signal_10202, mcs1_mcs_mat1_7_mcs_out[124]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6665], Fresh[6664], Fresh[6663], Fresh[6662], Fresh[6661], Fresh[6660]}), .c ({new_AGEMA_signal_11341, new_AGEMA_signal_11340, new_AGEMA_signal_11339, mcs1_mcs_mat1_7_mcs_rom0_28_x3x4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U8 ( .a ({new_AGEMA_signal_16594, new_AGEMA_signal_16593, new_AGEMA_signal_16592, mcs1_mcs_mat1_7_mcs_rom0_29_n8}), .b ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .c ({new_AGEMA_signal_17383, new_AGEMA_signal_17382, new_AGEMA_signal_17381, mcs1_mcs_mat1_7_mcs_out[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U7 ( .a ({new_AGEMA_signal_18673, new_AGEMA_signal_18672, new_AGEMA_signal_18671, mcs1_mcs_mat1_7_mcs_rom0_29_n7}), .b ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .c ({new_AGEMA_signal_19336, new_AGEMA_signal_19335, new_AGEMA_signal_19334, mcs1_mcs_mat1_7_mcs_out[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U6 ( .a ({new_AGEMA_signal_18037, new_AGEMA_signal_18036, new_AGEMA_signal_18035, mcs1_mcs_mat1_7_mcs_rom0_29_n6}), .b ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .c ({new_AGEMA_signal_18670, new_AGEMA_signal_18669, new_AGEMA_signal_18668, mcs1_mcs_mat1_7_mcs_out[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U5 ( .a ({new_AGEMA_signal_17386, new_AGEMA_signal_17385, new_AGEMA_signal_17384, mcs1_mcs_mat1_7_mcs_rom0_29_x3x4}), .b ({new_AGEMA_signal_16594, new_AGEMA_signal_16593, new_AGEMA_signal_16592, mcs1_mcs_mat1_7_mcs_rom0_29_n8}), .c ({new_AGEMA_signal_18037, new_AGEMA_signal_18036, new_AGEMA_signal_18035, mcs1_mcs_mat1_7_mcs_rom0_29_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U4 ( .a ({new_AGEMA_signal_14236, new_AGEMA_signal_14235, new_AGEMA_signal_14234, mcs1_mcs_mat1_7_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_15670, new_AGEMA_signal_15669, new_AGEMA_signal_15668, mcs1_mcs_mat1_7_mcs_rom0_29_x2x4}), .c ({new_AGEMA_signal_16594, new_AGEMA_signal_16593, new_AGEMA_signal_16592, mcs1_mcs_mat1_7_mcs_rom0_29_n8}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U3 ( .a ({new_AGEMA_signal_19339, new_AGEMA_signal_19338, new_AGEMA_signal_19337, mcs1_mcs_mat1_7_mcs_rom0_29_n5}), .b ({new_AGEMA_signal_11386, new_AGEMA_signal_11385, new_AGEMA_signal_11384, shiftr_out[64]}), .c ({new_AGEMA_signal_20041, new_AGEMA_signal_20040, new_AGEMA_signal_20039, mcs1_mcs_mat1_7_mcs_out[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U2 ( .a ({new_AGEMA_signal_14236, new_AGEMA_signal_14235, new_AGEMA_signal_14234, mcs1_mcs_mat1_7_mcs_rom0_29_x0x4}), .b ({new_AGEMA_signal_18673, new_AGEMA_signal_18672, new_AGEMA_signal_18671, mcs1_mcs_mat1_7_mcs_rom0_29_n7}), .c ({new_AGEMA_signal_19339, new_AGEMA_signal_19338, new_AGEMA_signal_19337, mcs1_mcs_mat1_7_mcs_rom0_29_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_U1 ( .a ({new_AGEMA_signal_18040, new_AGEMA_signal_18039, new_AGEMA_signal_18038, mcs1_mcs_mat1_7_mcs_rom0_29_x1x4}), .b ({new_AGEMA_signal_17386, new_AGEMA_signal_17385, new_AGEMA_signal_17384, mcs1_mcs_mat1_7_mcs_rom0_29_x3x4}), .c ({new_AGEMA_signal_18673, new_AGEMA_signal_18672, new_AGEMA_signal_18671, mcs1_mcs_mat1_7_mcs_rom0_29_n7}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x1x4_AND_U1 ( .a ({new_AGEMA_signal_16612, new_AGEMA_signal_16611, new_AGEMA_signal_16610, mcs1_mcs_mat1_7_mcs_out[91]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6671], Fresh[6670], Fresh[6669], Fresh[6668], Fresh[6667], Fresh[6666]}), .c ({new_AGEMA_signal_18040, new_AGEMA_signal_18039, new_AGEMA_signal_18038, mcs1_mcs_mat1_7_mcs_rom0_29_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x2x4_AND_U1 ( .a ({new_AGEMA_signal_12826, new_AGEMA_signal_12825, new_AGEMA_signal_12824, mcs1_mcs_mat1_7_mcs_out[88]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6677], Fresh[6676], Fresh[6675], Fresh[6674], Fresh[6673], Fresh[6672]}), .c ({new_AGEMA_signal_15670, new_AGEMA_signal_15669, new_AGEMA_signal_15668, mcs1_mcs_mat1_7_mcs_rom0_29_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_29_x3x4_AND_U1 ( .a ({new_AGEMA_signal_15700, new_AGEMA_signal_15699, new_AGEMA_signal_15698, shiftr_out[67]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6683], Fresh[6682], Fresh[6681], Fresh[6680], Fresh[6679], Fresh[6678]}), .c ({new_AGEMA_signal_17386, new_AGEMA_signal_17385, new_AGEMA_signal_17384, mcs1_mcs_mat1_7_mcs_rom0_29_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U6 ( .a ({new_AGEMA_signal_17389, new_AGEMA_signal_17388, new_AGEMA_signal_17387, mcs1_mcs_mat1_7_mcs_rom0_30_n7}), .b ({new_AGEMA_signal_11347, new_AGEMA_signal_11346, new_AGEMA_signal_11345, mcs1_mcs_mat1_7_mcs_rom0_30_x3x4}), .c ({new_AGEMA_signal_18043, new_AGEMA_signal_18042, new_AGEMA_signal_18041, mcs1_mcs_mat1_7_mcs_out[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U5 ( .a ({new_AGEMA_signal_16597, new_AGEMA_signal_16596, new_AGEMA_signal_16595, mcs1_mcs_mat1_7_mcs_out[7]}), .b ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .c ({new_AGEMA_signal_17389, new_AGEMA_signal_17388, new_AGEMA_signal_17387, mcs1_mcs_mat1_7_mcs_rom0_30_n7}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U4 ( .a ({new_AGEMA_signal_15673, new_AGEMA_signal_15672, new_AGEMA_signal_15671, mcs1_mcs_mat1_7_mcs_rom0_30_n6}), .b ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .c ({new_AGEMA_signal_16597, new_AGEMA_signal_16596, new_AGEMA_signal_16595, mcs1_mcs_mat1_7_mcs_out[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U3 ( .a ({new_AGEMA_signal_14239, new_AGEMA_signal_14238, new_AGEMA_signal_14237, mcs1_mcs_mat1_7_mcs_out[6]}), .b ({new_AGEMA_signal_10054, new_AGEMA_signal_10053, new_AGEMA_signal_10052, mcs1_mcs_mat1_7_mcs_rom0_30_x2x4}), .c ({new_AGEMA_signal_15673, new_AGEMA_signal_15672, new_AGEMA_signal_15671, mcs1_mcs_mat1_7_mcs_rom0_30_n6}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_U2 ( .a ({new_AGEMA_signal_10051, new_AGEMA_signal_10050, new_AGEMA_signal_10049, mcs1_mcs_mat1_7_mcs_rom0_30_n5}), .b ({new_AGEMA_signal_12793, new_AGEMA_signal_12792, new_AGEMA_signal_12791, mcs1_mcs_mat1_7_mcs_rom0_30_x1x4}), .c ({new_AGEMA_signal_14239, new_AGEMA_signal_14238, new_AGEMA_signal_14237, mcs1_mcs_mat1_7_mcs_out[6]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10438, new_AGEMA_signal_10437, new_AGEMA_signal_10436, shiftr_out[33]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6689], Fresh[6688], Fresh[6687], Fresh[6686], Fresh[6685], Fresh[6684]}), .c ({new_AGEMA_signal_12793, new_AGEMA_signal_12792, new_AGEMA_signal_12791, mcs1_mcs_mat1_7_mcs_rom0_30_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8602, new_AGEMA_signal_8601, new_AGEMA_signal_8600, shiftr_out[34]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6695], Fresh[6694], Fresh[6693], Fresh[6692], Fresh[6691], Fresh[6690]}), .c ({new_AGEMA_signal_10054, new_AGEMA_signal_10053, new_AGEMA_signal_10052, mcs1_mcs_mat1_7_mcs_rom0_30_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_30_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10240, new_AGEMA_signal_10239, new_AGEMA_signal_10238, mcs1_mcs_mat1_7_mcs_out[85]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6701], Fresh[6700], Fresh[6699], Fresh[6698], Fresh[6697], Fresh[6696]}), .c ({new_AGEMA_signal_11347, new_AGEMA_signal_11346, new_AGEMA_signal_11345, mcs1_mcs_mat1_7_mcs_rom0_30_x3x4}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U9 ( .a ({new_AGEMA_signal_11350, new_AGEMA_signal_11349, new_AGEMA_signal_11348, mcs1_mcs_mat1_7_mcs_rom0_31_n11}), .b ({new_AGEMA_signal_12796, new_AGEMA_signal_12795, new_AGEMA_signal_12794, mcs1_mcs_mat1_7_mcs_rom0_31_n10}), .c ({new_AGEMA_signal_14245, new_AGEMA_signal_14244, new_AGEMA_signal_14243, mcs1_mcs_mat1_7_mcs_out[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U8 ( .a ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .b ({new_AGEMA_signal_11353, new_AGEMA_signal_11352, new_AGEMA_signal_11351, mcs1_mcs_mat1_7_mcs_rom0_31_x3x4}), .c ({new_AGEMA_signal_12796, new_AGEMA_signal_12795, new_AGEMA_signal_12794, mcs1_mcs_mat1_7_mcs_rom0_31_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U7 ( .a ({new_AGEMA_signal_14248, new_AGEMA_signal_14247, new_AGEMA_signal_14246, mcs1_mcs_mat1_7_mcs_rom0_31_n9}), .b ({new_AGEMA_signal_10057, new_AGEMA_signal_10056, new_AGEMA_signal_10055, mcs1_mcs_mat1_7_mcs_rom0_31_x2x4}), .c ({new_AGEMA_signal_15676, new_AGEMA_signal_15675, new_AGEMA_signal_15674, mcs1_mcs_mat1_7_mcs_out[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U3 ( .a ({new_AGEMA_signal_14251, new_AGEMA_signal_14250, new_AGEMA_signal_14249, mcs1_mcs_mat1_7_mcs_rom0_31_n8}), .b ({new_AGEMA_signal_12802, new_AGEMA_signal_12801, new_AGEMA_signal_12800, mcs1_mcs_mat1_7_mcs_rom0_31_n7}), .c ({new_AGEMA_signal_15679, new_AGEMA_signal_15678, new_AGEMA_signal_15677, mcs1_mcs_mat1_7_mcs_out[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_U1 ( .a ({new_AGEMA_signal_12805, new_AGEMA_signal_12804, new_AGEMA_signal_12803, mcs1_mcs_mat1_7_mcs_rom0_31_x1x4}), .b ({new_AGEMA_signal_9139, new_AGEMA_signal_9138, new_AGEMA_signal_9137, mcs1_mcs_mat1_7_mcs_rom0_31_x0x4}), .c ({new_AGEMA_signal_14251, new_AGEMA_signal_14250, new_AGEMA_signal_14249, mcs1_mcs_mat1_7_mcs_rom0_31_n8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x1x4_AND_U1 ( .a ({new_AGEMA_signal_10456, new_AGEMA_signal_10455, new_AGEMA_signal_10454, shiftr_out[1]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6707], Fresh[6706], Fresh[6705], Fresh[6704], Fresh[6703], Fresh[6702]}), .c ({new_AGEMA_signal_12805, new_AGEMA_signal_12804, new_AGEMA_signal_12803, mcs1_mcs_mat1_7_mcs_rom0_31_x1x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x2x4_AND_U1 ( .a ({new_AGEMA_signal_8620, new_AGEMA_signal_8619, new_AGEMA_signal_8618, shiftr_out[2]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6713], Fresh[6712], Fresh[6711], Fresh[6710], Fresh[6709], Fresh[6708]}), .c ({new_AGEMA_signal_10057, new_AGEMA_signal_10056, new_AGEMA_signal_10055, mcs1_mcs_mat1_7_mcs_rom0_31_x2x4}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) mcs1_mcs_mat1_7_mcs_rom0_31_x3x4_AND_U1 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10257, new_AGEMA_signal_10256, mcs1_mcs_mat1_7_mcs_out[49]}), .b ({1'b0, 1'b0, 1'b0, p256_sel}), .clk (clk), .r ({Fresh[6719], Fresh[6718], Fresh[6717], Fresh[6716], Fresh[6715], Fresh[6714]}), .c ({new_AGEMA_signal_11353, new_AGEMA_signal_11352, new_AGEMA_signal_11351, mcs1_mcs_mat1_7_mcs_rom0_31_x3x4}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_0_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21346, new_AGEMA_signal_21345, new_AGEMA_signal_21344, mcs_out[128]}), .a ({new_AGEMA_signal_21406, new_AGEMA_signal_21405, new_AGEMA_signal_21404, y0_1[0]}), .c ({y0_s3[0], y0_s2[0], y0_s1[0], y0_s0[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_1_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20005, new_AGEMA_signal_20004, new_AGEMA_signal_20003, mcs_out[129]}), .a ({new_AGEMA_signal_20095, new_AGEMA_signal_20094, new_AGEMA_signal_20093, y0_1[1]}), .c ({y0_s3[1], y0_s2[1], y0_s1[1], y0_s0[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_2_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21343, new_AGEMA_signal_21342, new_AGEMA_signal_21341, mcs_out[130]}), .a ({new_AGEMA_signal_21457, new_AGEMA_signal_21456, new_AGEMA_signal_21455, y0_1[2]}), .c ({y0_s3[2], y0_s2[2], y0_s1[2], y0_s0[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_3_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19276, new_AGEMA_signal_19275, new_AGEMA_signal_19274, mcs_out[131]}), .a ({new_AGEMA_signal_19396, new_AGEMA_signal_19395, new_AGEMA_signal_19394, y0_1[3]}), .c ({y0_s3[3], y0_s2[3], y0_s1[3], y0_s0[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_4_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20704, new_AGEMA_signal_20703, new_AGEMA_signal_20702, mcs_out[132]}), .a ({new_AGEMA_signal_20869, new_AGEMA_signal_20868, new_AGEMA_signal_20867, y0_1[4]}), .c ({y0_s3[4], y0_s2[4], y0_s1[4], y0_s0[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_5_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21316, new_AGEMA_signal_21315, new_AGEMA_signal_21314, mcs_out[133]}), .a ({new_AGEMA_signal_21463, new_AGEMA_signal_21462, new_AGEMA_signal_21461, y0_1[5]}), .c ({y0_s3[5], y0_s2[5], y0_s1[5], y0_s0[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_6_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21313, new_AGEMA_signal_21312, new_AGEMA_signal_21311, mcs_out[134]}), .a ({new_AGEMA_signal_21472, new_AGEMA_signal_21471, new_AGEMA_signal_21470, y0_1[6]}), .c ({y0_s3[6], y0_s2[6], y0_s1[6], y0_s0[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_7_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20695, new_AGEMA_signal_20694, new_AGEMA_signal_20693, mcs_out[135]}), .a ({new_AGEMA_signal_20893, new_AGEMA_signal_20892, new_AGEMA_signal_20891, y0_1[7]}), .c ({y0_s3[7], y0_s2[7], y0_s1[7], y0_s0[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_8_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21700, new_AGEMA_signal_21699, new_AGEMA_signal_21698, mcs_out[136]}), .a ({new_AGEMA_signal_21793, new_AGEMA_signal_21792, new_AGEMA_signal_21791, y0_1[8]}), .c ({y0_s3[8], y0_s2[8], y0_s1[8], y0_s0[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_9_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19141, new_AGEMA_signal_19140, new_AGEMA_signal_19139, mcs_out[137]}), .a ({new_AGEMA_signal_19423, new_AGEMA_signal_19422, new_AGEMA_signal_19421, y0_1[9]}), .c ({y0_s3[9], y0_s2[9], y0_s1[9], y0_s0[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_10_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20650, new_AGEMA_signal_20649, new_AGEMA_signal_20648, mcs_out[138]}), .a ({new_AGEMA_signal_20836, new_AGEMA_signal_20835, new_AGEMA_signal_20834, y0_1[10]}), .c ({y0_s3[10], y0_s2[10], y0_s1[10], y0_s0[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_11_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21289, new_AGEMA_signal_21288, new_AGEMA_signal_21287, mcs_out[139]}), .a ({new_AGEMA_signal_21430, new_AGEMA_signal_21429, new_AGEMA_signal_21428, y0_1[11]}), .c ({y0_s3[11], y0_s2[11], y0_s1[11], y0_s0[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_12_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21268, new_AGEMA_signal_21267, new_AGEMA_signal_21266, mcs_out[140]}), .a ({new_AGEMA_signal_21436, new_AGEMA_signal_21435, new_AGEMA_signal_21434, y0_1[12]}), .c ({y0_s3[12], y0_s2[12], y0_s1[12], y0_s0[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_13_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19057, new_AGEMA_signal_19056, new_AGEMA_signal_19055, mcs_out[141]}), .a ({new_AGEMA_signal_19381, new_AGEMA_signal_19380, new_AGEMA_signal_19379, y0_1[13]}), .c ({y0_s3[13], y0_s2[13], y0_s1[13], y0_s0[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_14_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_17734, new_AGEMA_signal_17733, new_AGEMA_signal_17732, mcs_out[142]}), .a ({new_AGEMA_signal_18064, new_AGEMA_signal_18063, new_AGEMA_signal_18062, y0_1[14]}), .c ({y0_s3[14], y0_s2[14], y0_s1[14], y0_s0[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_15_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20605, new_AGEMA_signal_20604, new_AGEMA_signal_20603, mcs_out[143]}), .a ({new_AGEMA_signal_20848, new_AGEMA_signal_20847, new_AGEMA_signal_20846, y0_1[15]}), .c ({y0_s3[15], y0_s2[15], y0_s1[15], y0_s0[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_16_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21235, new_AGEMA_signal_21234, new_AGEMA_signal_21233, mcs_out[144]}), .a ({new_AGEMA_signal_21439, new_AGEMA_signal_21438, new_AGEMA_signal_21437, y0_1[16]}), .c ({y0_s3[16], y0_s2[16], y0_s1[16], y0_s0[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_17_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19720, new_AGEMA_signal_19719, new_AGEMA_signal_19718, mcs_out[145]}), .a ({new_AGEMA_signal_20092, new_AGEMA_signal_20091, new_AGEMA_signal_20090, y0_1[17]}), .c ({y0_s3[17], y0_s2[17], y0_s1[17], y0_s0[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_18_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21232, new_AGEMA_signal_21231, new_AGEMA_signal_21230, mcs_out[146]}), .a ({new_AGEMA_signal_21442, new_AGEMA_signal_21441, new_AGEMA_signal_21440, y0_1[18]}), .c ({y0_s3[18], y0_s2[18], y0_s1[18], y0_s0[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_19_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18979, new_AGEMA_signal_18978, new_AGEMA_signal_18977, mcs_out[147]}), .a ({new_AGEMA_signal_19384, new_AGEMA_signal_19383, new_AGEMA_signal_19382, y0_1[19]}), .c ({y0_s3[19], y0_s2[19], y0_s1[19], y0_s0[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_20_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20497, new_AGEMA_signal_20496, new_AGEMA_signal_20495, mcs_out[148]}), .a ({new_AGEMA_signal_20851, new_AGEMA_signal_20850, new_AGEMA_signal_20849, y0_1[20]}), .c ({y0_s3[20], y0_s2[20], y0_s1[20], y0_s0[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_21_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21205, new_AGEMA_signal_21204, new_AGEMA_signal_21203, mcs_out[149]}), .a ({new_AGEMA_signal_21445, new_AGEMA_signal_21444, new_AGEMA_signal_21443, y0_1[21]}), .c ({y0_s3[21], y0_s2[21], y0_s1[21], y0_s0[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_22_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21202, new_AGEMA_signal_21201, new_AGEMA_signal_21200, mcs_out[150]}), .a ({new_AGEMA_signal_21448, new_AGEMA_signal_21447, new_AGEMA_signal_21446, y0_1[22]}), .c ({y0_s3[22], y0_s2[22], y0_s1[22], y0_s0[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_23_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20488, new_AGEMA_signal_20487, new_AGEMA_signal_20486, mcs_out[151]}), .a ({new_AGEMA_signal_20854, new_AGEMA_signal_20853, new_AGEMA_signal_20852, y0_1[23]}), .c ({y0_s3[23], y0_s2[23], y0_s1[23], y0_s0[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_24_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21682, new_AGEMA_signal_21681, new_AGEMA_signal_21680, mcs_out[152]}), .a ({new_AGEMA_signal_21790, new_AGEMA_signal_21789, new_AGEMA_signal_21788, y0_1[24]}), .c ({y0_s3[24], y0_s2[24], y0_s1[24], y0_s0[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_25_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18844, new_AGEMA_signal_18843, new_AGEMA_signal_18842, mcs_out[153]}), .a ({new_AGEMA_signal_19387, new_AGEMA_signal_19386, new_AGEMA_signal_19385, y0_1[25]}), .c ({y0_s3[25], y0_s2[25], y0_s1[25], y0_s0[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_26_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20443, new_AGEMA_signal_20442, new_AGEMA_signal_20441, mcs_out[154]}), .a ({new_AGEMA_signal_20857, new_AGEMA_signal_20856, new_AGEMA_signal_20855, y0_1[26]}), .c ({y0_s3[26], y0_s2[26], y0_s1[26], y0_s0[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_27_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21178, new_AGEMA_signal_21177, new_AGEMA_signal_21176, mcs_out[155]}), .a ({new_AGEMA_signal_21451, new_AGEMA_signal_21450, new_AGEMA_signal_21449, y0_1[27]}), .c ({y0_s3[27], y0_s2[27], y0_s1[27], y0_s0[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_28_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21157, new_AGEMA_signal_21156, new_AGEMA_signal_21155, mcs_out[156]}), .a ({new_AGEMA_signal_21454, new_AGEMA_signal_21453, new_AGEMA_signal_21452, y0_1[28]}), .c ({y0_s3[28], y0_s2[28], y0_s1[28], y0_s0[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_29_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18760, new_AGEMA_signal_18759, new_AGEMA_signal_18758, mcs_out[157]}), .a ({new_AGEMA_signal_19390, new_AGEMA_signal_19389, new_AGEMA_signal_19388, y0_1[29]}), .c ({y0_s3[29], y0_s2[29], y0_s1[29], y0_s0[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_30_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_17407, new_AGEMA_signal_17406, new_AGEMA_signal_17405, mcs_out[158]}), .a ({new_AGEMA_signal_18067, new_AGEMA_signal_18066, new_AGEMA_signal_18065, y0_1[30]}), .c ({y0_s3[30], y0_s2[30], y0_s1[30], y0_s0[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_31_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20398, new_AGEMA_signal_20397, new_AGEMA_signal_20396, mcs_out[159]}), .a ({new_AGEMA_signal_20860, new_AGEMA_signal_20859, new_AGEMA_signal_20858, y0_1[31]}), .c ({y0_s3[31], y0_s2[31], y0_s1[31], y0_s0[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_32_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_17974, new_AGEMA_signal_17973, new_AGEMA_signal_17972, mcs_out[160]}), .a ({new_AGEMA_signal_18070, new_AGEMA_signal_18069, new_AGEMA_signal_18068, y0_1[32]}), .c ({y0_s3[32], y0_s2[32], y0_s1[32], y0_s0[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_33_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18613, new_AGEMA_signal_18612, new_AGEMA_signal_18611, mcs_out[161]}), .a ({new_AGEMA_signal_18688, new_AGEMA_signal_18687, new_AGEMA_signal_18686, y0_1[33]}), .c ({y0_s3[33], y0_s2[33], y0_s1[33], y0_s0[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_34_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18610, new_AGEMA_signal_18609, new_AGEMA_signal_18608, mcs_out[162]}), .a ({new_AGEMA_signal_18691, new_AGEMA_signal_18690, new_AGEMA_signal_18689, y0_1[34]}), .c ({y0_s3[34], y0_s2[34], y0_s1[34], y0_s0[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_35_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18607, new_AGEMA_signal_18606, new_AGEMA_signal_18605, mcs_out[163]}), .a ({new_AGEMA_signal_18694, new_AGEMA_signal_18693, new_AGEMA_signal_18692, y0_1[35]}), .c ({y0_s3[35], y0_s2[35], y0_s1[35], y0_s0[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_36_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19927, new_AGEMA_signal_19926, new_AGEMA_signal_19925, mcs_out[164]}), .a ({new_AGEMA_signal_20098, new_AGEMA_signal_20097, new_AGEMA_signal_20096, y0_1[36]}), .c ({y0_s3[36], y0_s2[36], y0_s1[36], y0_s0[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_37_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_17881, new_AGEMA_signal_17880, new_AGEMA_signal_17879, mcs_out[165]}), .a ({new_AGEMA_signal_18073, new_AGEMA_signal_18072, new_AGEMA_signal_18071, y0_1[37]}), .c ({y0_s3[37], y0_s2[37], y0_s1[37], y0_s0[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_38_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_16396, new_AGEMA_signal_16395, new_AGEMA_signal_16394, mcs_out[166]}), .a ({new_AGEMA_signal_16600, new_AGEMA_signal_16599, new_AGEMA_signal_16598, y0_1[38]}), .c ({y0_s3[38], y0_s2[38], y0_s1[38], y0_s0[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_39_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19207, new_AGEMA_signal_19206, new_AGEMA_signal_19205, mcs_out[167]}), .a ({new_AGEMA_signal_19393, new_AGEMA_signal_19392, new_AGEMA_signal_19391, y0_1[39]}), .c ({y0_s3[39], y0_s2[39], y0_s1[39], y0_s0[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_40_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20641, new_AGEMA_signal_20640, new_AGEMA_signal_20639, mcs_out[168]}), .a ({new_AGEMA_signal_20863, new_AGEMA_signal_20862, new_AGEMA_signal_20861, y0_1[40]}), .c ({y0_s3[40], y0_s2[40], y0_s1[40], y0_s0[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_41_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19855, new_AGEMA_signal_19854, new_AGEMA_signal_19853, mcs_out[169]}), .a ({new_AGEMA_signal_20101, new_AGEMA_signal_20100, new_AGEMA_signal_20099, y0_1[41]}), .c ({y0_s3[41], y0_s2[41], y0_s1[41], y0_s0[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_42_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19852, new_AGEMA_signal_19851, new_AGEMA_signal_19850, mcs_out[170]}), .a ({new_AGEMA_signal_20104, new_AGEMA_signal_20103, new_AGEMA_signal_20102, y0_1[42]}), .c ({y0_s3[42], y0_s2[42], y0_s1[42], y0_s0[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_43_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19849, new_AGEMA_signal_19848, new_AGEMA_signal_19847, mcs_out[171]}), .a ({new_AGEMA_signal_20107, new_AGEMA_signal_20106, new_AGEMA_signal_20105, y0_1[43]}), .c ({y0_s3[43], y0_s2[43], y0_s1[43], y0_s0[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_44_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21265, new_AGEMA_signal_21264, new_AGEMA_signal_21263, mcs_out[172]}), .a ({new_AGEMA_signal_21460, new_AGEMA_signal_21459, new_AGEMA_signal_21458, y0_1[44]}), .c ({y0_s3[44], y0_s2[44], y0_s1[44], y0_s0[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_45_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19054, new_AGEMA_signal_19053, new_AGEMA_signal_19052, mcs_out[173]}), .a ({new_AGEMA_signal_19399, new_AGEMA_signal_19398, new_AGEMA_signal_19397, y0_1[45]}), .c ({y0_s3[45], y0_s2[45], y0_s1[45], y0_s0[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_46_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19051, new_AGEMA_signal_19050, new_AGEMA_signal_19049, mcs_out[174]}), .a ({new_AGEMA_signal_19402, new_AGEMA_signal_19401, new_AGEMA_signal_19400, y0_1[46]}), .c ({y0_s3[46], y0_s2[46], y0_s1[46], y0_s0[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_47_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20596, new_AGEMA_signal_20595, new_AGEMA_signal_20594, mcs_out[175]}), .a ({new_AGEMA_signal_20866, new_AGEMA_signal_20865, new_AGEMA_signal_20864, y0_1[47]}), .c ({y0_s3[47], y0_s2[47], y0_s1[47], y0_s0[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_48_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_17647, new_AGEMA_signal_17646, new_AGEMA_signal_17645, mcs_out[176]}), .a ({new_AGEMA_signal_18076, new_AGEMA_signal_18075, new_AGEMA_signal_18074, y0_1[48]}), .c ({y0_s3[48], y0_s2[48], y0_s1[48], y0_s0[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_49_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18334, new_AGEMA_signal_18333, new_AGEMA_signal_18332, mcs_out[177]}), .a ({new_AGEMA_signal_18697, new_AGEMA_signal_18696, new_AGEMA_signal_18695, y0_1[49]}), .c ({y0_s3[49], y0_s2[49], y0_s1[49], y0_s0[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_50_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18331, new_AGEMA_signal_18330, new_AGEMA_signal_18329, mcs_out[178]}), .a ({new_AGEMA_signal_18700, new_AGEMA_signal_18699, new_AGEMA_signal_18698, y0_1[50]}), .c ({y0_s3[50], y0_s2[50], y0_s1[50], y0_s0[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_51_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18328, new_AGEMA_signal_18327, new_AGEMA_signal_18326, mcs_out[179]}), .a ({new_AGEMA_signal_18703, new_AGEMA_signal_18702, new_AGEMA_signal_18701, y0_1[51]}), .c ({y0_s3[51], y0_s2[51], y0_s1[51], y0_s0[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_52_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19642, new_AGEMA_signal_19641, new_AGEMA_signal_19640, mcs_out[180]}), .a ({new_AGEMA_signal_20110, new_AGEMA_signal_20109, new_AGEMA_signal_20108, y0_1[52]}), .c ({y0_s3[52], y0_s2[52], y0_s1[52], y0_s0[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_53_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_17554, new_AGEMA_signal_17553, new_AGEMA_signal_17552, mcs_out[181]}), .a ({new_AGEMA_signal_18079, new_AGEMA_signal_18078, new_AGEMA_signal_18077, y0_1[53]}), .c ({y0_s3[53], y0_s2[53], y0_s1[53], y0_s0[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_54_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_15955, new_AGEMA_signal_15954, new_AGEMA_signal_15953, mcs_out[182]}), .a ({new_AGEMA_signal_16603, new_AGEMA_signal_16602, new_AGEMA_signal_16601, y0_1[54]}), .c ({y0_s3[54], y0_s2[54], y0_s1[54], y0_s0[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_55_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18910, new_AGEMA_signal_18909, new_AGEMA_signal_18908, mcs_out[183]}), .a ({new_AGEMA_signal_19405, new_AGEMA_signal_19404, new_AGEMA_signal_19403, y0_1[55]}), .c ({y0_s3[55], y0_s2[55], y0_s1[55], y0_s0[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_56_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20434, new_AGEMA_signal_20433, new_AGEMA_signal_20432, mcs_out[184]}), .a ({new_AGEMA_signal_20872, new_AGEMA_signal_20871, new_AGEMA_signal_20870, y0_1[56]}), .c ({y0_s3[56], y0_s2[56], y0_s1[56], y0_s0[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_57_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19570, new_AGEMA_signal_19569, new_AGEMA_signal_19568, mcs_out[185]}), .a ({new_AGEMA_signal_20113, new_AGEMA_signal_20112, new_AGEMA_signal_20111, y0_1[57]}), .c ({y0_s3[57], y0_s2[57], y0_s1[57], y0_s0[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_58_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19567, new_AGEMA_signal_19566, new_AGEMA_signal_19565, mcs_out[186]}), .a ({new_AGEMA_signal_20116, new_AGEMA_signal_20115, new_AGEMA_signal_20114, y0_1[58]}), .c ({y0_s3[58], y0_s2[58], y0_s1[58], y0_s0[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_59_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19564, new_AGEMA_signal_19563, new_AGEMA_signal_19562, mcs_out[187]}), .a ({new_AGEMA_signal_20119, new_AGEMA_signal_20118, new_AGEMA_signal_20117, y0_1[59]}), .c ({y0_s3[59], y0_s2[59], y0_s1[59], y0_s0[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_60_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21154, new_AGEMA_signal_21153, new_AGEMA_signal_21152, mcs_out[188]}), .a ({new_AGEMA_signal_21466, new_AGEMA_signal_21465, new_AGEMA_signal_21464, y0_1[60]}), .c ({y0_s3[60], y0_s2[60], y0_s1[60], y0_s0[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_61_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18757, new_AGEMA_signal_18756, new_AGEMA_signal_18755, mcs_out[189]}), .a ({new_AGEMA_signal_19408, new_AGEMA_signal_19407, new_AGEMA_signal_19406, y0_1[61]}), .c ({y0_s3[61], y0_s2[61], y0_s1[61], y0_s0[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_62_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18754, new_AGEMA_signal_18753, new_AGEMA_signal_18752, mcs_out[190]}), .a ({new_AGEMA_signal_19411, new_AGEMA_signal_19410, new_AGEMA_signal_19409, y0_1[62]}), .c ({y0_s3[62], y0_s2[62], y0_s1[62], y0_s0[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_63_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20389, new_AGEMA_signal_20388, new_AGEMA_signal_20387, mcs_out[191]}), .a ({new_AGEMA_signal_20875, new_AGEMA_signal_20874, new_AGEMA_signal_20873, y0_1[63]}), .c ({y0_s3[63], y0_s2[63], y0_s1[63], y0_s0[63]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_64_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21340, new_AGEMA_signal_21339, new_AGEMA_signal_21338, mcs_out[192]}), .a ({new_AGEMA_signal_21469, new_AGEMA_signal_21468, new_AGEMA_signal_21467, y0_1[64]}), .c ({y0_s3[64], y0_s2[64], y0_s1[64], y0_s0[64]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_65_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20752, new_AGEMA_signal_20751, new_AGEMA_signal_20750, mcs_out[193]}), .a ({new_AGEMA_signal_20878, new_AGEMA_signal_20877, new_AGEMA_signal_20876, y0_1[65]}), .c ({y0_s3[65], y0_s2[65], y0_s1[65], y0_s0[65]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_66_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20749, new_AGEMA_signal_20748, new_AGEMA_signal_20747, mcs_out[194]}), .a ({new_AGEMA_signal_20881, new_AGEMA_signal_20880, new_AGEMA_signal_20879, y0_1[66]}), .c ({y0_s3[66], y0_s2[66], y0_s1[66], y0_s0[66]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_67_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20746, new_AGEMA_signal_20745, new_AGEMA_signal_20744, mcs_out[195]}), .a ({new_AGEMA_signal_20884, new_AGEMA_signal_20883, new_AGEMA_signal_20882, y0_1[67]}), .c ({y0_s3[67], y0_s2[67], y0_s1[67], y0_s0[67]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_68_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20692, new_AGEMA_signal_20691, new_AGEMA_signal_20690, mcs_out[196]}), .a ({new_AGEMA_signal_20887, new_AGEMA_signal_20886, new_AGEMA_signal_20885, y0_1[68]}), .c ({y0_s3[68], y0_s2[68], y0_s1[68], y0_s0[68]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_69_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19921, new_AGEMA_signal_19920, new_AGEMA_signal_19919, mcs_out[197]}), .a ({new_AGEMA_signal_20122, new_AGEMA_signal_20121, new_AGEMA_signal_20120, y0_1[69]}), .c ({y0_s3[69], y0_s2[69], y0_s1[69], y0_s0[69]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_70_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19201, new_AGEMA_signal_19200, new_AGEMA_signal_19199, mcs_out[198]}), .a ({new_AGEMA_signal_19414, new_AGEMA_signal_19413, new_AGEMA_signal_19412, y0_1[70]}), .c ({y0_s3[70], y0_s2[70], y0_s1[70], y0_s0[70]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_71_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20689, new_AGEMA_signal_20688, new_AGEMA_signal_20687, mcs_out[199]}), .a ({new_AGEMA_signal_20890, new_AGEMA_signal_20889, new_AGEMA_signal_20888, y0_1[71]}), .c ({y0_s3[71], y0_s2[71], y0_s1[71], y0_s0[71]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_72_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21838, new_AGEMA_signal_21837, new_AGEMA_signal_21836, mcs_out[200]}), .a ({new_AGEMA_signal_21952, new_AGEMA_signal_21951, new_AGEMA_signal_21950, y0_1[72]}), .c ({y0_s3[72], y0_s2[72], y0_s1[72], y0_s0[72]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_73_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18466, new_AGEMA_signal_18465, new_AGEMA_signal_18464, mcs_out[201]}), .a ({new_AGEMA_signal_18706, new_AGEMA_signal_18705, new_AGEMA_signal_18704, y0_1[73]}), .c ({y0_s3[73], y0_s2[73], y0_s1[73], y0_s0[73]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_74_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19846, new_AGEMA_signal_19845, new_AGEMA_signal_19844, mcs_out[202]}), .a ({new_AGEMA_signal_20125, new_AGEMA_signal_20124, new_AGEMA_signal_20123, y0_1[74]}), .c ({y0_s3[74], y0_s2[74], y0_s1[74], y0_s0[74]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_75_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21286, new_AGEMA_signal_21285, new_AGEMA_signal_21284, mcs_out[203]}), .a ({new_AGEMA_signal_21475, new_AGEMA_signal_21474, new_AGEMA_signal_21473, y0_1[75]}), .c ({y0_s3[75], y0_s2[75], y0_s1[75], y0_s0[75]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_76_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21262, new_AGEMA_signal_21261, new_AGEMA_signal_21260, mcs_out[204]}), .a ({new_AGEMA_signal_21478, new_AGEMA_signal_21477, new_AGEMA_signal_21476, y0_1[76]}), .c ({y0_s3[76], y0_s2[76], y0_s1[76], y0_s0[76]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_77_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21259, new_AGEMA_signal_21258, new_AGEMA_signal_21257, mcs_out[205]}), .a ({new_AGEMA_signal_21481, new_AGEMA_signal_21480, new_AGEMA_signal_21479, y0_1[77]}), .c ({y0_s3[77], y0_s2[77], y0_s1[77], y0_s0[77]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_78_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21256, new_AGEMA_signal_21255, new_AGEMA_signal_21254, mcs_out[206]}), .a ({new_AGEMA_signal_21484, new_AGEMA_signal_21483, new_AGEMA_signal_21482, y0_1[78]}), .c ({y0_s3[78], y0_s2[78], y0_s1[78], y0_s0[78]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_79_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21253, new_AGEMA_signal_21252, new_AGEMA_signal_21251, mcs_out[207]}), .a ({new_AGEMA_signal_21487, new_AGEMA_signal_21486, new_AGEMA_signal_21485, y0_1[79]}), .c ({y0_s3[79], y0_s2[79], y0_s1[79], y0_s0[79]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_80_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21229, new_AGEMA_signal_21228, new_AGEMA_signal_21227, mcs_out[208]}), .a ({new_AGEMA_signal_21490, new_AGEMA_signal_21489, new_AGEMA_signal_21488, y0_1[80]}), .c ({y0_s3[80], y0_s2[80], y0_s1[80], y0_s0[80]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_81_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20545, new_AGEMA_signal_20544, new_AGEMA_signal_20543, mcs_out[209]}), .a ({new_AGEMA_signal_20896, new_AGEMA_signal_20895, new_AGEMA_signal_20894, y0_1[81]}), .c ({y0_s3[81], y0_s2[81], y0_s1[81], y0_s0[81]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_82_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20542, new_AGEMA_signal_20541, new_AGEMA_signal_20540, mcs_out[210]}), .a ({new_AGEMA_signal_20899, new_AGEMA_signal_20898, new_AGEMA_signal_20897, y0_1[82]}), .c ({y0_s3[82], y0_s2[82], y0_s1[82], y0_s0[82]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_83_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20539, new_AGEMA_signal_20538, new_AGEMA_signal_20537, mcs_out[211]}), .a ({new_AGEMA_signal_20902, new_AGEMA_signal_20901, new_AGEMA_signal_20900, y0_1[83]}), .c ({y0_s3[83], y0_s2[83], y0_s1[83], y0_s0[83]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_84_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20485, new_AGEMA_signal_20484, new_AGEMA_signal_20483, mcs_out[212]}), .a ({new_AGEMA_signal_20905, new_AGEMA_signal_20904, new_AGEMA_signal_20903, y0_1[84]}), .c ({y0_s3[84], y0_s2[84], y0_s1[84], y0_s0[84]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_85_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19636, new_AGEMA_signal_19635, new_AGEMA_signal_19634, mcs_out[213]}), .a ({new_AGEMA_signal_20128, new_AGEMA_signal_20127, new_AGEMA_signal_20126, y0_1[85]}), .c ({y0_s3[85], y0_s2[85], y0_s1[85], y0_s0[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_86_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18904, new_AGEMA_signal_18903, new_AGEMA_signal_18902, mcs_out[214]}), .a ({new_AGEMA_signal_19417, new_AGEMA_signal_19416, new_AGEMA_signal_19415, y0_1[86]}), .c ({y0_s3[86], y0_s2[86], y0_s1[86], y0_s0[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_87_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20482, new_AGEMA_signal_20481, new_AGEMA_signal_20480, mcs_out[215]}), .a ({new_AGEMA_signal_20908, new_AGEMA_signal_20907, new_AGEMA_signal_20906, y0_1[87]}), .c ({y0_s3[87], y0_s2[87], y0_s1[87], y0_s0[87]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_88_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21832, new_AGEMA_signal_21831, new_AGEMA_signal_21830, mcs_out[216]}), .a ({new_AGEMA_signal_21955, new_AGEMA_signal_21954, new_AGEMA_signal_21953, y0_1[88]}), .c ({y0_s3[88], y0_s2[88], y0_s1[88], y0_s0[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_89_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18187, new_AGEMA_signal_18186, new_AGEMA_signal_18185, mcs_out[217]}), .a ({new_AGEMA_signal_18709, new_AGEMA_signal_18708, new_AGEMA_signal_18707, y0_1[89]}), .c ({y0_s3[89], y0_s2[89], y0_s1[89], y0_s0[89]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_90_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19561, new_AGEMA_signal_19560, new_AGEMA_signal_19559, mcs_out[218]}), .a ({new_AGEMA_signal_20131, new_AGEMA_signal_20130, new_AGEMA_signal_20129, y0_1[90]}), .c ({y0_s3[90], y0_s2[90], y0_s1[90], y0_s0[90]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_91_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21175, new_AGEMA_signal_21174, new_AGEMA_signal_21173, mcs_out[219]}), .a ({new_AGEMA_signal_21493, new_AGEMA_signal_21492, new_AGEMA_signal_21491, y0_1[91]}), .c ({y0_s3[91], y0_s2[91], y0_s1[91], y0_s0[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_92_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21151, new_AGEMA_signal_21150, new_AGEMA_signal_21149, mcs_out[220]}), .a ({new_AGEMA_signal_21496, new_AGEMA_signal_21495, new_AGEMA_signal_21494, y0_1[92]}), .c ({y0_s3[92], y0_s2[92], y0_s1[92], y0_s0[92]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_93_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21148, new_AGEMA_signal_21147, new_AGEMA_signal_21146, mcs_out[221]}), .a ({new_AGEMA_signal_21499, new_AGEMA_signal_21498, new_AGEMA_signal_21497, y0_1[93]}), .c ({y0_s3[93], y0_s2[93], y0_s1[93], y0_s0[93]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_94_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21145, new_AGEMA_signal_21144, new_AGEMA_signal_21143, mcs_out[222]}), .a ({new_AGEMA_signal_21502, new_AGEMA_signal_21501, new_AGEMA_signal_21500, y0_1[94]}), .c ({y0_s3[94], y0_s2[94], y0_s1[94], y0_s0[94]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_95_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21142, new_AGEMA_signal_21141, new_AGEMA_signal_21140, mcs_out[223]}), .a ({new_AGEMA_signal_21505, new_AGEMA_signal_21504, new_AGEMA_signal_21503, y0_1[95]}), .c ({y0_s3[95], y0_s2[95], y0_s1[95], y0_s0[95]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_96_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20743, new_AGEMA_signal_20742, new_AGEMA_signal_20741, mcs_out[224]}), .a ({new_AGEMA_signal_20911, new_AGEMA_signal_20910, new_AGEMA_signal_20909, y0_1[96]}), .c ({y0_s3[96], y0_s2[96], y0_s1[96], y0_s0[96]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_97_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21337, new_AGEMA_signal_21336, new_AGEMA_signal_21335, mcs_out[225]}), .a ({new_AGEMA_signal_21508, new_AGEMA_signal_21507, new_AGEMA_signal_21506, y0_1[97]}), .c ({y0_s3[97], y0_s2[97], y0_s1[97], y0_s0[97]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_98_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19270, new_AGEMA_signal_19269, new_AGEMA_signal_19268, mcs_out[226]}), .a ({new_AGEMA_signal_19420, new_AGEMA_signal_19419, new_AGEMA_signal_19418, y0_1[98]}), .c ({y0_s3[98], y0_s2[98], y0_s1[98], y0_s0[98]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_99_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21334, new_AGEMA_signal_21333, new_AGEMA_signal_21332, mcs_out[227]}), .a ({new_AGEMA_signal_21511, new_AGEMA_signal_21510, new_AGEMA_signal_21509, y0_1[99]}), .c ({y0_s3[99], y0_s2[99], y0_s1[99], y0_s0[99]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_100_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19915, new_AGEMA_signal_19914, new_AGEMA_signal_19913, mcs_out[228]}), .a ({new_AGEMA_signal_20080, new_AGEMA_signal_20079, new_AGEMA_signal_20078, y0_1[100]}), .c ({y0_s3[100], y0_s2[100], y0_s1[100], y0_s0[100]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_101_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20686, new_AGEMA_signal_20685, new_AGEMA_signal_20684, mcs_out[229]}), .a ({new_AGEMA_signal_20830, new_AGEMA_signal_20829, new_AGEMA_signal_20828, y0_1[101]}), .c ({y0_s3[101], y0_s2[101], y0_s1[101], y0_s0[101]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_102_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21310, new_AGEMA_signal_21309, new_AGEMA_signal_21308, mcs_out[230]}), .a ({new_AGEMA_signal_21409, new_AGEMA_signal_21408, new_AGEMA_signal_21407, y0_1[102]}), .c ({y0_s3[102], y0_s2[102], y0_s1[102], y0_s0[102]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_103_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21307, new_AGEMA_signal_21306, new_AGEMA_signal_21305, mcs_out[231]}), .a ({new_AGEMA_signal_21412, new_AGEMA_signal_21411, new_AGEMA_signal_21410, y0_1[103]}), .c ({y0_s3[103], y0_s2[103], y0_s1[103], y0_s0[103]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_104_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21283, new_AGEMA_signal_21282, new_AGEMA_signal_21281, mcs_out[232]}), .a ({new_AGEMA_signal_21415, new_AGEMA_signal_21414, new_AGEMA_signal_21413, y0_1[104]}), .c ({y0_s3[104], y0_s2[104], y0_s1[104], y0_s0[104]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_105_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19126, new_AGEMA_signal_19125, new_AGEMA_signal_19124, mcs_out[233]}), .a ({new_AGEMA_signal_19372, new_AGEMA_signal_19371, new_AGEMA_signal_19370, y0_1[105]}), .c ({y0_s3[105], y0_s2[105], y0_s1[105], y0_s0[105]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_106_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19840, new_AGEMA_signal_19839, new_AGEMA_signal_19838, mcs_out[234]}), .a ({new_AGEMA_signal_20083, new_AGEMA_signal_20082, new_AGEMA_signal_20081, y0_1[106]}), .c ({y0_s3[106], y0_s2[106], y0_s1[106], y0_s0[106]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_107_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20632, new_AGEMA_signal_20631, new_AGEMA_signal_20630, mcs_out[235]}), .a ({new_AGEMA_signal_20833, new_AGEMA_signal_20832, new_AGEMA_signal_20831, y0_1[107]}), .c ({y0_s3[107], y0_s2[107], y0_s1[107], y0_s0[107]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_108_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_17731, new_AGEMA_signal_17730, new_AGEMA_signal_17729, mcs_out[236]}), .a ({new_AGEMA_signal_18052, new_AGEMA_signal_18051, new_AGEMA_signal_18050, y0_1[108]}), .c ({y0_s3[108], y0_s2[108], y0_s1[108], y0_s0[108]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_109_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18403, new_AGEMA_signal_18402, new_AGEMA_signal_18401, mcs_out[237]}), .a ({new_AGEMA_signal_18676, new_AGEMA_signal_18675, new_AGEMA_signal_18674, y0_1[109]}), .c ({y0_s3[109], y0_s2[109], y0_s1[109], y0_s0[109]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_110_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18400, new_AGEMA_signal_18399, new_AGEMA_signal_18398, mcs_out[238]}), .a ({new_AGEMA_signal_18679, new_AGEMA_signal_18678, new_AGEMA_signal_18677, y0_1[110]}), .c ({y0_s3[110], y0_s2[110], y0_s1[110], y0_s0[110]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_111_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_17722, new_AGEMA_signal_17721, new_AGEMA_signal_17720, mcs_out[239]}), .a ({new_AGEMA_signal_18055, new_AGEMA_signal_18054, new_AGEMA_signal_18053, y0_1[111]}), .c ({y0_s3[111], y0_s2[111], y0_s1[111], y0_s0[111]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_112_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20536, new_AGEMA_signal_20535, new_AGEMA_signal_20534, mcs_out[240]}), .a ({new_AGEMA_signal_20839, new_AGEMA_signal_20838, new_AGEMA_signal_20837, y0_1[112]}), .c ({y0_s3[112], y0_s2[112], y0_s1[112], y0_s0[112]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_113_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21226, new_AGEMA_signal_21225, new_AGEMA_signal_21224, mcs_out[241]}), .a ({new_AGEMA_signal_21418, new_AGEMA_signal_21417, new_AGEMA_signal_21416, y0_1[113]}), .c ({y0_s3[113], y0_s2[113], y0_s1[113], y0_s0[113]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_114_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18973, new_AGEMA_signal_18972, new_AGEMA_signal_18971, mcs_out[242]}), .a ({new_AGEMA_signal_19375, new_AGEMA_signal_19374, new_AGEMA_signal_19373, y0_1[114]}), .c ({y0_s3[114], y0_s2[114], y0_s1[114], y0_s0[114]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_115_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21223, new_AGEMA_signal_21222, new_AGEMA_signal_21221, mcs_out[243]}), .a ({new_AGEMA_signal_21421, new_AGEMA_signal_21420, new_AGEMA_signal_21419, y0_1[115]}), .c ({y0_s3[115], y0_s2[115], y0_s1[115], y0_s0[115]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_116_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19630, new_AGEMA_signal_19629, new_AGEMA_signal_19628, mcs_out[244]}), .a ({new_AGEMA_signal_20086, new_AGEMA_signal_20085, new_AGEMA_signal_20084, y0_1[116]}), .c ({y0_s3[116], y0_s2[116], y0_s1[116], y0_s0[116]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_117_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20479, new_AGEMA_signal_20478, new_AGEMA_signal_20477, mcs_out[245]}), .a ({new_AGEMA_signal_20842, new_AGEMA_signal_20841, new_AGEMA_signal_20840, y0_1[117]}), .c ({y0_s3[117], y0_s2[117], y0_s1[117], y0_s0[117]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_118_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21199, new_AGEMA_signal_21198, new_AGEMA_signal_21197, mcs_out[246]}), .a ({new_AGEMA_signal_21424, new_AGEMA_signal_21423, new_AGEMA_signal_21422, y0_1[118]}), .c ({y0_s3[118], y0_s2[118], y0_s1[118], y0_s0[118]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_119_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21196, new_AGEMA_signal_21195, new_AGEMA_signal_21194, mcs_out[247]}), .a ({new_AGEMA_signal_21427, new_AGEMA_signal_21426, new_AGEMA_signal_21425, y0_1[119]}), .c ({y0_s3[119], y0_s2[119], y0_s1[119], y0_s0[119]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_120_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_21172, new_AGEMA_signal_21171, new_AGEMA_signal_21170, mcs_out[248]}), .a ({new_AGEMA_signal_21433, new_AGEMA_signal_21432, new_AGEMA_signal_21431, y0_1[120]}), .c ({y0_s3[120], y0_s2[120], y0_s1[120], y0_s0[120]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_121_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18829, new_AGEMA_signal_18828, new_AGEMA_signal_18827, mcs_out[249]}), .a ({new_AGEMA_signal_19378, new_AGEMA_signal_19377, new_AGEMA_signal_19376, y0_1[121]}), .c ({y0_s3[121], y0_s2[121], y0_s1[121], y0_s0[121]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_122_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_19555, new_AGEMA_signal_19554, new_AGEMA_signal_19553, mcs_out[250]}), .a ({new_AGEMA_signal_20089, new_AGEMA_signal_20088, new_AGEMA_signal_20087, y0_1[122]}), .c ({y0_s3[122], y0_s2[122], y0_s1[122], y0_s0[122]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_123_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_20425, new_AGEMA_signal_20424, new_AGEMA_signal_20423, mcs_out[251]}), .a ({new_AGEMA_signal_20845, new_AGEMA_signal_20844, new_AGEMA_signal_20843, y0_1[123]}), .c ({y0_s3[123], y0_s2[123], y0_s1[123], y0_s0[123]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_124_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_17404, new_AGEMA_signal_17403, new_AGEMA_signal_17402, mcs_out[252]}), .a ({new_AGEMA_signal_18058, new_AGEMA_signal_18057, new_AGEMA_signal_18056, y0_1[124]}), .c ({y0_s3[124], y0_s2[124], y0_s1[124], y0_s0[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_125_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18124, new_AGEMA_signal_18123, new_AGEMA_signal_18122, mcs_out[253]}), .a ({new_AGEMA_signal_18682, new_AGEMA_signal_18681, new_AGEMA_signal_18680, y0_1[125]}), .c ({y0_s3[125], y0_s2[125], y0_s1[125], y0_s0[125]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_126_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_18121, new_AGEMA_signal_18120, new_AGEMA_signal_18119, mcs_out[254]}), .a ({new_AGEMA_signal_18685, new_AGEMA_signal_18684, new_AGEMA_signal_18683, y0_1[126]}), .c ({y0_s3[126], y0_s2[126], y0_s1[126], y0_s0[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) MUX_inst2_MUXInst_127_U1 ( .s (p256_sel), .b ({new_AGEMA_signal_17395, new_AGEMA_signal_17394, new_AGEMA_signal_17393, mcs_out[255]}), .a ({new_AGEMA_signal_18061, new_AGEMA_signal_18060, new_AGEMA_signal_18059, y0_1[127]}), .c ({y0_s3[127], y0_s2[127], y0_s1[127], y0_s0[127]}) ) ;

endmodule
